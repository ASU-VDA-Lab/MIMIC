module real_aes_6224_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_1106;
wire n_1170;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_1175;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_635;
wire n_503;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_1192;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_979;
wire n_759;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1197;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_1113;
wire n_852;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1137;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_1040;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_892;
wire n_495;
wire n_994;
wire n_1072;
wire n_1078;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_1182;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_1189;
wire n_1180;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_656;
wire n_532;
wire n_1025;
wire n_755;
wire n_1168;
wire n_1148;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_455;
wire n_504;
wire n_973;
wire n_725;
wire n_671;
wire n_1084;
wire n_960;
wire n_1081;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1196;
wire n_737;
wire n_1013;
wire n_1017;
wire n_936;
wire n_581;
wire n_610;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_1100;
wire n_1167;
wire n_1174;
wire n_1193;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_754;
wire n_607;
wire n_449;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_1031;
wire n_432;
wire n_880;
wire n_1037;
wire n_1131;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_999;
wire n_913;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_1179;
wire n_1171;
wire n_569;
wire n_563;
wire n_785;
wire n_997;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1157;
wire n_1158;
wire n_1132;
wire n_853;
wire n_1079;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1003;
wire n_1028;
wire n_1000;
wire n_1014;
wire n_1187;
wire n_1083;
wire n_727;
wire n_649;
wire n_663;
wire n_1056;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_1043;
wire n_850;
wire n_1136;
wire n_720;
wire n_1127;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_717;
wire n_456;
wire n_1090;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_705;
wire n_1191;
wire n_1195;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1186;
wire n_1010;
wire n_811;
wire n_823;
wire n_459;
wire n_558;
wire n_1015;
wire n_1172;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1184;
wire n_1166;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_1143;
wire n_929;
wire n_1190;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_1156;
wire n_1159;
wire n_829;
wire n_1030;
wire n_988;
wire n_1088;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1176;
wire n_1151;
wire n_1036;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_968;
wire n_652;
wire n_703;
wire n_1097;
wire n_601;
wire n_1101;
wire n_1102;
wire n_661;
wire n_500;
wire n_463;
wire n_804;
wire n_1076;
wire n_447;
wire n_1185;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_1039;
wire n_424;
wire n_802;
wire n_868;
wire n_877;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_1061;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx20_ASAP7_75t_R g1153 ( .A(n_0), .Y(n_1153) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_1), .A2(n_165), .B1(n_546), .B2(n_549), .Y(n_899) );
INVx1_ASAP7_75t_L g894 ( .A(n_2), .Y(n_894) );
AOI22xp33_ASAP7_75t_SL g954 ( .A1(n_3), .A2(n_134), .B1(n_549), .B2(n_754), .Y(n_954) );
CKINVDCx20_ASAP7_75t_R g880 ( .A(n_4), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_5), .A2(n_103), .B1(n_656), .B2(n_777), .Y(n_1040) );
AO22x2_ASAP7_75t_L g428 ( .A1(n_6), .A2(n_233), .B1(n_420), .B2(n_425), .Y(n_428) );
INVx1_ASAP7_75t_L g1139 ( .A(n_6), .Y(n_1139) );
CKINVDCx20_ASAP7_75t_R g984 ( .A(n_7), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_8), .A2(n_152), .B1(n_440), .B2(n_471), .Y(n_748) );
AOI222xp33_ASAP7_75t_L g958 ( .A1(n_9), .A2(n_335), .B1(n_347), .B2(n_486), .C1(n_578), .C2(n_847), .Y(n_958) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_10), .Y(n_910) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_11), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g982 ( .A(n_12), .Y(n_982) );
INVx1_ASAP7_75t_L g740 ( .A(n_13), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_14), .A2(n_56), .B1(n_908), .B2(n_909), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_15), .A2(n_129), .B1(n_555), .B2(n_560), .Y(n_1157) );
AOI22xp33_ASAP7_75t_SL g598 ( .A1(n_16), .A2(n_116), .B1(n_599), .B2(n_601), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g1011 ( .A1(n_17), .A2(n_205), .B1(n_650), .B2(n_805), .C(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g721 ( .A(n_18), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g577 ( .A1(n_19), .A2(n_293), .B1(n_486), .B2(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g728 ( .A(n_20), .Y(n_728) );
INVx1_ASAP7_75t_L g1073 ( .A(n_21), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_22), .A2(n_328), .B1(n_466), .B2(n_469), .Y(n_465) );
AOI22xp5_ASAP7_75t_SL g765 ( .A1(n_23), .A2(n_199), .B1(n_628), .B2(n_766), .Y(n_765) );
AOI22xp33_ASAP7_75t_SL g595 ( .A1(n_24), .A2(n_268), .B1(n_444), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_25), .A2(n_95), .B1(n_486), .B2(n_578), .Y(n_876) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_26), .A2(n_217), .B1(n_439), .B2(n_444), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1184 ( .A1(n_27), .A2(n_381), .B1(n_619), .B2(n_654), .Y(n_1184) );
AOI22xp33_ASAP7_75t_SL g895 ( .A1(n_28), .A2(n_200), .B1(n_580), .B2(n_614), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_29), .A2(n_158), .B1(n_622), .B2(n_941), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_30), .A2(n_110), .B1(n_526), .B2(n_633), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_31), .A2(n_331), .B1(n_909), .B2(n_1113), .Y(n_1112) );
CKINVDCx20_ASAP7_75t_R g1005 ( .A(n_32), .Y(n_1005) );
AOI22xp33_ASAP7_75t_SL g1042 ( .A1(n_33), .A2(n_138), .B1(n_529), .B2(n_1043), .Y(n_1042) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_34), .A2(n_84), .B1(n_544), .B2(n_548), .Y(n_617) );
AO22x2_ASAP7_75t_L g430 ( .A1(n_35), .A2(n_115), .B1(n_420), .B2(n_421), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_36), .A2(n_258), .B1(n_544), .B2(n_549), .Y(n_841) );
AOI222xp33_ASAP7_75t_L g759 ( .A1(n_37), .A2(n_198), .B1(n_307), .B2(n_548), .C1(n_580), .C2(n_611), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g1008 ( .A(n_38), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_39), .A2(n_224), .B1(n_531), .B2(n_1190), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_40), .A2(n_322), .B1(n_433), .B2(n_861), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_41), .B(n_1039), .Y(n_1038) );
CKINVDCx20_ASAP7_75t_R g1154 ( .A(n_42), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_43), .A2(n_67), .B1(n_472), .B2(n_632), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_44), .A2(n_267), .B1(n_726), .B2(n_941), .Y(n_940) );
CKINVDCx20_ASAP7_75t_R g1056 ( .A(n_45), .Y(n_1056) );
CKINVDCx20_ASAP7_75t_R g1016 ( .A(n_46), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g1095 ( .A(n_47), .Y(n_1095) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_48), .A2(n_117), .B1(n_592), .B2(n_593), .Y(n_591) );
AOI22xp33_ASAP7_75t_SL g621 ( .A1(n_49), .A2(n_378), .B1(n_622), .B2(n_623), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g1161 ( .A1(n_50), .A2(n_180), .B1(n_469), .B2(n_1048), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_51), .A2(n_80), .B1(n_689), .B2(n_975), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_52), .B(n_567), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_53), .A2(n_100), .B1(n_692), .B2(n_829), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_54), .Y(n_464) );
INVx1_ASAP7_75t_L g714 ( .A(n_55), .Y(n_714) );
INVx1_ASAP7_75t_L g556 ( .A(n_57), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_58), .A2(n_144), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22x1_ASAP7_75t_L g1078 ( .A1(n_59), .A2(n_1079), .B1(n_1101), .B2(n_1102), .Y(n_1078) );
CKINVDCx20_ASAP7_75t_R g1101 ( .A(n_59), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_60), .A2(n_88), .B1(n_439), .B2(n_628), .Y(n_1158) );
AOI22xp33_ASAP7_75t_SL g630 ( .A1(n_61), .A2(n_120), .B1(n_631), .B2(n_632), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g972 ( .A(n_62), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_63), .A2(n_238), .B1(n_564), .B2(n_692), .Y(n_906) );
AO22x1_ASAP7_75t_L g994 ( .A1(n_64), .A2(n_995), .B1(n_1026), .B2(n_1027), .Y(n_994) );
INVx1_ASAP7_75t_L g1026 ( .A(n_64), .Y(n_1026) );
AOI222xp33_ASAP7_75t_L g812 ( .A1(n_65), .A2(n_181), .B1(n_357), .B2(n_495), .C1(n_615), .C2(n_783), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_66), .A2(n_97), .B1(n_855), .B2(n_885), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_68), .A2(n_321), .B1(n_450), .B2(n_564), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g980 ( .A(n_69), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_70), .A2(n_193), .B1(n_544), .B2(n_656), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_71), .A2(n_86), .B1(n_587), .B2(n_1118), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_72), .A2(n_382), .B1(n_689), .B2(n_855), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_73), .B(n_587), .Y(n_953) );
AOI22xp33_ASAP7_75t_SL g1047 ( .A1(n_74), .A2(n_395), .B1(n_769), .B2(n_1048), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_75), .A2(n_348), .B1(n_802), .B2(n_805), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_76), .A2(n_342), .B1(n_858), .B2(n_859), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_77), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_78), .A2(n_390), .B1(n_544), .B2(n_548), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g1063 ( .A(n_79), .Y(n_1063) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_81), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_82), .A2(n_209), .B1(n_858), .B2(n_909), .Y(n_1160) );
CKINVDCx20_ASAP7_75t_R g968 ( .A(n_83), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_85), .A2(n_287), .B1(n_549), .B2(n_1120), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_87), .A2(n_260), .B1(n_622), .B2(n_692), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_89), .Y(n_794) );
AO22x2_ASAP7_75t_L g424 ( .A1(n_90), .A2(n_266), .B1(n_420), .B2(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g1136 ( .A(n_90), .Y(n_1136) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_91), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g1082 ( .A(n_92), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_93), .A2(n_147), .B1(n_777), .B2(n_844), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_94), .A2(n_107), .B1(n_469), .B2(n_555), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_96), .A2(n_229), .B1(n_777), .B2(n_778), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_98), .A2(n_289), .B1(n_452), .B2(n_564), .Y(n_888) );
CKINVDCx20_ASAP7_75t_R g1093 ( .A(n_99), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_101), .A2(n_194), .B1(n_583), .B2(n_654), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_102), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_104), .A2(n_790), .B1(n_813), .B2(n_814), .Y(n_789) );
CKINVDCx16_ASAP7_75t_R g813 ( .A(n_104), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_105), .A2(n_387), .B1(n_487), .B2(n_754), .Y(n_753) );
AOI222xp33_ASAP7_75t_L g831 ( .A1(n_106), .A2(n_112), .B1(n_184), .B2(n_494), .C1(n_578), .C2(n_589), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_108), .A2(n_836), .B1(n_862), .B2(n_863), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_108), .Y(n_862) );
XOR2x2_ASAP7_75t_L g923 ( .A(n_109), .B(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g781 ( .A(n_111), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_113), .A2(n_285), .B1(n_592), .B2(n_624), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_114), .A2(n_275), .B1(n_472), .B2(n_757), .Y(n_764) );
INVx1_ASAP7_75t_L g1140 ( .A(n_115), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_118), .A2(n_270), .B1(n_770), .B2(n_1085), .Y(n_1084) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_119), .A2(n_309), .B1(n_769), .B2(n_770), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g1146 ( .A(n_121), .Y(n_1146) );
CKINVDCx20_ASAP7_75t_R g1096 ( .A(n_122), .Y(n_1096) );
CKINVDCx20_ASAP7_75t_R g1181 ( .A(n_123), .Y(n_1181) );
XOR2x2_ASAP7_75t_L g571 ( .A(n_124), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_125), .B(n_936), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_126), .A2(n_282), .B1(n_726), .B2(n_772), .Y(n_887) );
CKINVDCx20_ASAP7_75t_R g998 ( .A(n_127), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_128), .Y(n_809) );
AO22x1_ASAP7_75t_L g1105 ( .A1(n_130), .A2(n_1106), .B1(n_1107), .B2(n_1122), .Y(n_1105) );
CKINVDCx20_ASAP7_75t_R g1122 ( .A(n_130), .Y(n_1122) );
CKINVDCx20_ASAP7_75t_R g1092 ( .A(n_131), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_132), .A2(n_149), .B1(n_445), .B2(n_627), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_133), .B(n_934), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_135), .A2(n_361), .B1(n_452), .B2(n_467), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_136), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g839 ( .A(n_137), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_139), .A2(n_143), .B1(n_592), .B2(n_624), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g1100 ( .A(n_140), .Y(n_1100) );
AOI22xp33_ASAP7_75t_SL g1183 ( .A1(n_141), .A2(n_218), .B1(n_656), .B2(n_1120), .Y(n_1183) );
CKINVDCx20_ASAP7_75t_R g1009 ( .A(n_142), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_145), .A2(n_359), .B1(n_533), .B2(n_596), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_146), .A2(n_162), .B1(n_628), .B2(n_855), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_148), .A2(n_370), .B1(n_635), .B2(n_805), .Y(n_942) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_150), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g1150 ( .A(n_151), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_153), .A2(n_206), .B1(n_614), .B2(n_615), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_154), .A2(n_215), .B1(n_548), .B2(n_754), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_155), .A2(n_312), .B1(n_555), .B2(n_633), .Y(n_949) );
AOI22xp33_ASAP7_75t_SL g634 ( .A1(n_156), .A2(n_353), .B1(n_635), .B2(n_637), .Y(n_634) );
AOI22xp33_ASAP7_75t_SL g884 ( .A1(n_157), .A2(n_257), .B1(n_596), .B2(n_885), .Y(n_884) );
AND2x6_ASAP7_75t_L g403 ( .A(n_159), .B(n_404), .Y(n_403) );
HB1xp67_ASAP7_75t_L g1133 ( .A(n_159), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_160), .A2(n_292), .B1(n_531), .B2(n_533), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_161), .A2(n_343), .B1(n_487), .B2(n_580), .Y(n_1061) );
AOI22xp33_ASAP7_75t_SL g1035 ( .A1(n_163), .A2(n_271), .B1(n_567), .B2(n_735), .Y(n_1035) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_164), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_166), .A2(n_346), .B1(n_628), .B2(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_167), .A2(n_333), .B1(n_531), .B2(n_689), .Y(n_688) );
AOI222xp33_ASAP7_75t_L g566 ( .A1(n_168), .A2(n_246), .B1(n_265), .B2(n_487), .C1(n_495), .C2(n_567), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_169), .Y(n_959) );
INVx1_ASAP7_75t_L g568 ( .A(n_170), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_171), .A2(n_320), .B1(n_526), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_SL g1050 ( .A1(n_172), .A2(n_350), .B1(n_723), .B2(n_772), .Y(n_1050) );
CKINVDCx20_ASAP7_75t_R g1087 ( .A(n_173), .Y(n_1087) );
AOI22xp33_ASAP7_75t_SL g904 ( .A1(n_174), .A2(n_372), .B1(n_627), .B2(n_750), .Y(n_904) );
INVx1_ASAP7_75t_L g1025 ( .A(n_175), .Y(n_1025) );
INVx1_ASAP7_75t_L g738 ( .A(n_176), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_177), .A2(n_326), .B1(n_650), .B2(n_772), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g1003 ( .A(n_178), .Y(n_1003) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_179), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_182), .A2(n_262), .B1(n_439), .B2(n_444), .Y(n_1089) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_183), .A2(n_253), .B1(n_531), .B2(n_662), .Y(n_944) );
CKINVDCx20_ASAP7_75t_R g973 ( .A(n_185), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_186), .A2(n_360), .B1(n_624), .B2(n_903), .Y(n_1072) );
AO22x2_ASAP7_75t_L g419 ( .A1(n_187), .A2(n_254), .B1(n_420), .B2(n_421), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g1137 ( .A(n_187), .B(n_1138), .Y(n_1137) );
CKINVDCx20_ASAP7_75t_R g987 ( .A(n_188), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_189), .A2(n_226), .B1(n_461), .B2(n_533), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_190), .Y(n_952) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_191), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_192), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_195), .A2(n_385), .B1(n_661), .B2(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g1034 ( .A(n_196), .Y(n_1034) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_197), .Y(n_576) );
AOI222xp33_ASAP7_75t_L g1121 ( .A1(n_201), .A2(n_341), .B1(n_349), .B2(n_494), .C1(n_614), .C2(n_664), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_202), .A2(n_259), .B1(n_555), .B2(n_659), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g1147 ( .A(n_203), .Y(n_1147) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_204), .A2(n_355), .B1(n_626), .B2(n_628), .Y(n_625) );
XOR2x2_ASAP7_75t_L g816 ( .A(n_207), .B(n_817), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_208), .A2(n_283), .B1(n_540), .B2(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_210), .A2(n_315), .B1(n_583), .B2(n_775), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_211), .Y(n_760) );
OA22x2_ASAP7_75t_L g709 ( .A1(n_212), .A2(n_710), .B1(n_711), .B2(n_743), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_212), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_213), .Y(n_810) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_214), .A2(n_399), .B(n_408), .C(n_1141), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g1019 ( .A1(n_216), .A2(n_304), .B1(n_526), .B2(n_1020), .C(n_1022), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_219), .A2(n_397), .B1(n_462), .B2(n_804), .Y(n_1192) );
CKINVDCx20_ASAP7_75t_R g1178 ( .A(n_220), .Y(n_1178) );
INVx1_ASAP7_75t_L g558 ( .A(n_221), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_222), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_223), .A2(n_310), .B1(n_775), .B2(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_225), .B(n_615), .Y(n_985) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_227), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g1097 ( .A(n_228), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_230), .A2(n_274), .B1(n_467), .B2(n_627), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_231), .B(n_583), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_232), .A2(n_302), .B1(n_593), .B2(n_825), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_234), .A2(n_325), .B1(n_549), .B2(n_732), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_235), .A2(n_291), .B1(n_529), .B2(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_236), .A2(n_305), .B1(n_544), .B2(n_589), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_237), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_239), .A2(n_384), .B1(n_445), .B2(n_757), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g1083 ( .A(n_240), .Y(n_1083) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_241), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g988 ( .A(n_242), .Y(n_988) );
INVx1_ASAP7_75t_L g552 ( .A(n_243), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_244), .A2(n_345), .B1(n_487), .B2(n_754), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_245), .A2(n_269), .B1(n_445), .B2(n_627), .Y(n_806) );
AOI222xp33_ASAP7_75t_L g663 ( .A1(n_247), .A2(n_362), .B1(n_373), .B2(n_495), .C1(n_614), .C2(n_664), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_248), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_249), .A2(n_383), .B1(n_903), .B2(n_1188), .Y(n_1187) );
INVx2_ASAP7_75t_L g407 ( .A(n_250), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_251), .A2(n_288), .B1(n_500), .B2(n_930), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g1142 ( .A1(n_252), .A2(n_1143), .B1(n_1162), .B2(n_1163), .Y(n_1142) );
CKINVDCx20_ASAP7_75t_R g1162 ( .A(n_252), .Y(n_1162) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_255), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_256), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_261), .A2(n_867), .B1(n_868), .B2(n_889), .Y(n_866) );
CKINVDCx14_ASAP7_75t_R g889 ( .A(n_261), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_263), .A2(n_308), .B1(n_580), .B2(n_783), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_264), .A2(n_377), .B1(n_466), .B2(n_1020), .Y(n_1109) );
INVx1_ASAP7_75t_L g1065 ( .A(n_272), .Y(n_1065) );
CKINVDCx20_ASAP7_75t_R g1149 ( .A(n_273), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_276), .A2(n_299), .B1(n_631), .B2(n_772), .Y(n_969) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_277), .Y(n_848) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_278), .Y(n_873) );
INVx1_ASAP7_75t_L g715 ( .A(n_279), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g602 ( .A1(n_280), .A2(n_393), .B1(n_471), .B2(n_603), .Y(n_602) );
XOR2x2_ASAP7_75t_L g1030 ( .A(n_281), .B(n_1031), .Y(n_1030) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_284), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g1171 ( .A(n_286), .Y(n_1171) );
OA22x2_ASAP7_75t_L g1172 ( .A1(n_286), .A2(n_1171), .B1(n_1173), .B2(n_1194), .Y(n_1172) );
INVx1_ASAP7_75t_L g420 ( .A(n_290), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_290), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_294), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_295), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_296), .A2(n_380), .B1(n_439), .B2(n_444), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_297), .A2(n_351), .B1(n_601), .B2(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_298), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g742 ( .A(n_300), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_301), .B(n_820), .Y(n_897) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_303), .A2(n_412), .B1(n_517), .B2(n_518), .Y(n_411) );
INVx1_ASAP7_75t_L g517 ( .A(n_303), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_306), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g1177 ( .A(n_311), .Y(n_1177) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_313), .Y(n_475) );
INVx1_ASAP7_75t_L g730 ( .A(n_314), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_316), .Y(n_798) );
INVx1_ASAP7_75t_L g1023 ( .A(n_317), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_318), .B(n_540), .Y(n_898) );
OA22x2_ASAP7_75t_L g605 ( .A1(n_319), .A2(n_606), .B1(n_607), .B2(n_639), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_319), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_323), .A2(n_391), .B1(n_585), .B2(n_587), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_324), .A2(n_363), .B1(n_638), .B2(n_694), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_327), .Y(n_687) );
INVx1_ASAP7_75t_L g406 ( .A(n_329), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_330), .Y(n_458) );
INVx1_ASAP7_75t_L g404 ( .A(n_332), .Y(n_404) );
INVx1_ASAP7_75t_L g784 ( .A(n_334), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g1099 ( .A(n_336), .Y(n_1099) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_337), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_338), .A2(n_344), .B1(n_433), .B2(n_757), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g1060 ( .A(n_339), .Y(n_1060) );
INVx1_ASAP7_75t_L g562 ( .A(n_340), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g1000 ( .A(n_352), .Y(n_1000) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_354), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g1088 ( .A(n_356), .Y(n_1088) );
CKINVDCx20_ASAP7_75t_R g979 ( .A(n_358), .Y(n_979) );
INVx1_ASAP7_75t_L g535 ( .A(n_364), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_365), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_366), .B(n_664), .Y(n_1006) );
AOI22xp33_ASAP7_75t_SL g902 ( .A1(n_367), .A2(n_389), .B1(n_659), .B2(n_903), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_368), .B(n_583), .Y(n_582) );
XOR2x2_ASAP7_75t_L g646 ( .A(n_369), .B(n_647), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_371), .A2(n_666), .B1(n_696), .B2(n_697), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_371), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_374), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_375), .B(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_376), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_379), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_386), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_388), .Y(n_1013) );
INVx1_ASAP7_75t_L g724 ( .A(n_392), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_394), .A2(n_963), .B1(n_989), .B2(n_990), .Y(n_962) );
CKINVDCx20_ASAP7_75t_R g989 ( .A(n_394), .Y(n_989) );
CKINVDCx20_ASAP7_75t_R g1058 ( .A(n_396), .Y(n_1058) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_400), .Y(n_399) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
HB1xp67_ASAP7_75t_L g1132 ( .A(n_404), .Y(n_1132) );
OAI21xp5_ASAP7_75t_L g1169 ( .A1(n_405), .A2(n_1131), .B(n_1170), .Y(n_1169) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_703), .B1(n_1126), .B2(n_1127), .C(n_1128), .Y(n_408) );
INVx1_ASAP7_75t_L g1127 ( .A(n_409), .Y(n_1127) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_519), .B1(n_701), .B2(n_702), .Y(n_409) );
INVx1_ASAP7_75t_L g701 ( .A(n_410), .Y(n_701) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g518 ( .A(n_412), .Y(n_518) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_473), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_448), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_431), .B1(n_432), .B2(n_437), .C(n_438), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g553 ( .A(n_416), .Y(n_553) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_426), .Y(n_417) );
AND2x2_ASAP7_75t_L g442 ( .A(n_418), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g600 ( .A(n_418), .B(n_426), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g1015 ( .A(n_418), .B(n_443), .Y(n_1015) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_423), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_419), .B(n_424), .Y(n_436) );
INVx2_ASAP7_75t_L g456 ( .A(n_419), .Y(n_456) );
AND2x2_ASAP7_75t_L g491 ( .A(n_419), .B(n_428), .Y(n_491) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_422), .Y(n_425) );
INVx1_ASAP7_75t_L g516 ( .A(n_423), .Y(n_516) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g457 ( .A(n_424), .Y(n_457) );
AND2x2_ASAP7_75t_L g463 ( .A(n_424), .B(n_456), .Y(n_463) );
INVx1_ASAP7_75t_L g490 ( .A(n_424), .Y(n_490) );
AND2x4_ASAP7_75t_L g434 ( .A(n_426), .B(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g462 ( .A(n_426), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g468 ( .A(n_426), .B(n_455), .Y(n_468) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
AND2x2_ASAP7_75t_L g443 ( .A(n_427), .B(n_430), .Y(n_443) );
OR2x2_ASAP7_75t_L g454 ( .A(n_427), .B(n_430), .Y(n_454) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g496 ( .A(n_428), .B(n_430), .Y(n_496) );
AND2x2_ASAP7_75t_L g489 ( .A(n_429), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g509 ( .A(n_429), .Y(n_509) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g447 ( .A(n_430), .Y(n_447) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
HB1xp67_ASAP7_75t_L g1085 ( .A(n_433), .Y(n_1085) );
BUFx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g555 ( .A(n_434), .Y(n_555) );
BUFx2_ASAP7_75t_SL g601 ( .A(n_434), .Y(n_601) );
BUFx3_ASAP7_75t_L g638 ( .A(n_434), .Y(n_638) );
BUFx2_ASAP7_75t_SL g772 ( .A(n_434), .Y(n_772) );
BUFx3_ASAP7_75t_L g805 ( .A(n_434), .Y(n_805) );
INVx1_ASAP7_75t_L g826 ( .A(n_434), .Y(n_826) );
BUFx2_ASAP7_75t_L g903 ( .A(n_434), .Y(n_903) );
AND2x2_ASAP7_75t_L g750 ( .A(n_435), .B(n_509), .Y(n_750) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OR2x6_ASAP7_75t_L g446 ( .A(n_436), .B(n_447), .Y(n_446) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_440), .Y(n_596) );
INVx5_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx3_ASAP7_75t_L g532 ( .A(n_441), .Y(n_532) );
INVx2_ASAP7_75t_L g627 ( .A(n_441), .Y(n_627) );
INVx4_ASAP7_75t_L g719 ( .A(n_441), .Y(n_719) );
INVx3_ASAP7_75t_L g855 ( .A(n_441), .Y(n_855) );
INVx1_ASAP7_75t_L g976 ( .A(n_441), .Y(n_976) );
INVx8_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g472 ( .A(n_443), .B(n_455), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g483 ( .A(n_443), .B(n_463), .Y(n_483) );
AND2x6_ASAP7_75t_L g585 ( .A(n_443), .B(n_463), .Y(n_585) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g533 ( .A(n_445), .Y(n_533) );
BUFx2_ASAP7_75t_L g628 ( .A(n_445), .Y(n_628) );
BUFx2_ASAP7_75t_L g885 ( .A(n_445), .Y(n_885) );
BUFx4f_ASAP7_75t_SL g1018 ( .A(n_445), .Y(n_1018) );
INVx6_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g689 ( .A(n_446), .Y(n_689) );
INVx1_ASAP7_75t_SL g1190 ( .A(n_446), .Y(n_1190) );
INVx1_ASAP7_75t_L g547 ( .A(n_447), .Y(n_547) );
OAI221xp5_ASAP7_75t_SL g448 ( .A1(n_449), .A2(n_458), .B1(n_459), .B2(n_464), .C(n_465), .Y(n_448) );
OAI221xp5_ASAP7_75t_SL g851 ( .A1(n_449), .A2(n_528), .B1(n_852), .B2(n_853), .C(n_854), .Y(n_851) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx4_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g661 ( .A(n_451), .Y(n_661) );
INVx2_ASAP7_75t_L g770 ( .A(n_451), .Y(n_770) );
INVx5_ASAP7_75t_SL g804 ( .A(n_451), .Y(n_804) );
INVx2_ASAP7_75t_SL g941 ( .A(n_451), .Y(n_941) );
HB1xp67_ASAP7_75t_L g1114 ( .A(n_451), .Y(n_1114) );
INVx11_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx11_ASAP7_75t_L g561 ( .A(n_452), .Y(n_561) );
AND2x6_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
AND2x4_ASAP7_75t_L g542 ( .A(n_453), .B(n_463), .Y(n_542) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g478 ( .A(n_454), .B(n_479), .Y(n_478) );
AND2x6_ASAP7_75t_L g495 ( .A(n_455), .B(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
OAI221xp5_ASAP7_75t_SL g1081 ( .A1(n_459), .A2(n_713), .B1(n_1082), .B2(n_1083), .C(n_1084), .Y(n_1081) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_462), .Y(n_529) );
INVx2_ASAP7_75t_L g594 ( .A(n_462), .Y(n_594) );
BUFx3_ASAP7_75t_L g624 ( .A(n_462), .Y(n_624) );
BUFx3_ASAP7_75t_L g909 ( .A(n_462), .Y(n_909) );
INVx1_ASAP7_75t_L g479 ( .A(n_463), .Y(n_479) );
BUFx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g713 ( .A(n_467), .Y(n_713) );
BUFx6f_ASAP7_75t_L g769 ( .A(n_467), .Y(n_769) );
BUFx3_ASAP7_75t_L g858 ( .A(n_467), .Y(n_858) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_SL g526 ( .A(n_468), .Y(n_526) );
BUFx2_ASAP7_75t_SL g592 ( .A(n_468), .Y(n_592) );
INVx2_ASAP7_75t_L g636 ( .A(n_468), .Y(n_636) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx6_ASAP7_75t_L g565 ( .A(n_472), .Y(n_565) );
BUFx3_ASAP7_75t_L g622 ( .A(n_472), .Y(n_622) );
BUFx3_ASAP7_75t_L g829 ( .A(n_472), .Y(n_829) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .C(n_504), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B1(n_480), .B2(n_481), .Y(n_474) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_476), .A2(n_728), .B1(n_729), .B2(n_730), .C(n_731), .Y(n_727) );
OAI221xp5_ASAP7_75t_SL g838 ( .A1(n_476), .A2(n_729), .B1(n_839), .B2(n_840), .C(n_841), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_476), .A2(n_481), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g872 ( .A(n_477), .Y(n_872) );
INVx1_ASAP7_75t_SL g999 ( .A(n_477), .Y(n_999) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_478), .Y(n_670) );
BUFx3_ASAP7_75t_L g1057 ( .A(n_478), .Y(n_1057) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g729 ( .A(n_482), .Y(n_729) );
INVx1_ASAP7_75t_SL g1001 ( .A(n_482), .Y(n_1001) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx3_ASAP7_75t_L g537 ( .A(n_483), .Y(n_537) );
OAI222xp33_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_492), .B1(n_493), .B2(n_497), .C1(n_498), .C2(n_503), .Y(n_484) );
OAI221xp5_ASAP7_75t_SL g1148 ( .A1(n_485), .A2(n_846), .B1(n_1149), .B2(n_1150), .C(n_1151), .Y(n_1148) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_SL g1004 ( .A(n_486), .Y(n_1004) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx4f_ASAP7_75t_SL g614 ( .A(n_488), .Y(n_614) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_488), .Y(n_737) );
BUFx2_ASAP7_75t_L g783 ( .A(n_488), .Y(n_783) );
BUFx6f_ASAP7_75t_L g844 ( .A(n_488), .Y(n_844) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
INVx1_ASAP7_75t_L g502 ( .A(n_490), .Y(n_502) );
AND2x4_ASAP7_75t_L g501 ( .A(n_491), .B(n_502), .Y(n_501) );
NAND2x1p5_ASAP7_75t_L g508 ( .A(n_491), .B(n_509), .Y(n_508) );
AND2x4_ASAP7_75t_L g546 ( .A(n_491), .B(n_547), .Y(n_546) );
OAI222xp33_ASAP7_75t_L g674 ( .A1(n_493), .A2(n_675), .B1(n_676), .B2(n_677), .C1(n_678), .C2(n_679), .Y(n_674) );
OAI222xp33_ASAP7_75t_L g1094 ( .A1(n_493), .A2(n_741), .B1(n_983), .B2(n_1095), .C1(n_1096), .C2(n_1097), .Y(n_1094) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_SL g575 ( .A(n_494), .Y(n_575) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx3_ASAP7_75t_L g611 ( .A(n_495), .Y(n_611) );
INVx4_ASAP7_75t_L g739 ( .A(n_495), .Y(n_739) );
INVx2_ASAP7_75t_SL g927 ( .A(n_495), .Y(n_927) );
INVx1_ASAP7_75t_L g514 ( .A(n_496), .Y(n_514) );
AND2x4_ASAP7_75t_L g549 ( .A(n_496), .B(n_516), .Y(n_549) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g615 ( .A(n_500), .Y(n_615) );
INVx2_ASAP7_75t_L g678 ( .A(n_500), .Y(n_678) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_501), .Y(n_567) );
BUFx12f_ASAP7_75t_L g580 ( .A(n_501), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B1(n_510), .B2(n_511), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_506), .A2(n_511), .B1(n_681), .B2(n_682), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_506), .A2(n_511), .B1(n_987), .B2(n_988), .Y(n_986) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_506), .A2(n_1008), .B1(n_1009), .B2(n_1010), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_506), .A2(n_511), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx4_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_508), .Y(n_879) );
BUFx3_ASAP7_75t_L g1064 ( .A(n_508), .Y(n_1064) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g1010 ( .A(n_512), .Y(n_1010) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_513), .A2(n_878), .B1(n_879), .B2(n_880), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_513), .A2(n_1063), .B1(n_1064), .B2(n_1065), .Y(n_1062) );
OR2x6_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g702 ( .A(n_519), .Y(n_702) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_642), .B1(n_699), .B2(n_700), .Y(n_520) );
INVx1_ASAP7_75t_L g699 ( .A(n_521), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_569), .B1(n_570), .B2(n_641), .Y(n_521) );
INVx2_ASAP7_75t_L g641 ( .A(n_522), .Y(n_641) );
XOR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_568), .Y(n_522) );
NAND4xp75_ASAP7_75t_L g523 ( .A(n_524), .B(n_534), .C(n_550), .D(n_566), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_530), .Y(n_524) );
INVx1_ASAP7_75t_L g685 ( .A(n_526), .Y(n_685) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx4_ASAP7_75t_L g650 ( .A(n_528), .Y(n_650) );
OAI221xp5_ASAP7_75t_SL g684 ( .A1(n_528), .A2(n_685), .B1(n_686), .B2(n_687), .C(n_688), .Y(n_684) );
OAI221xp5_ASAP7_75t_SL g712 ( .A1(n_528), .A2(n_713), .B1(n_714), .B2(n_715), .C(n_716), .Y(n_712) );
INVx4_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OA211x2_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B(n_538), .C(n_543), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_536), .A2(n_871), .B1(n_872), .B2(n_873), .Y(n_870) );
OA211x2_ASAP7_75t_L g951 ( .A1(n_536), .A2(n_952), .B(n_953), .C(n_954), .Y(n_951) );
BUFx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g673 ( .A(n_537), .Y(n_673) );
BUFx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx5_ASAP7_75t_L g587 ( .A(n_541), .Y(n_587) );
INVx2_ASAP7_75t_L g775 ( .A(n_541), .Y(n_775) );
INVx2_ASAP7_75t_L g1039 ( .A(n_541), .Y(n_1039) );
INVx4_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g732 ( .A(n_545), .Y(n_732) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
BUFx3_ASAP7_75t_L g754 ( .A(n_546), .Y(n_754) );
BUFx2_ASAP7_75t_L g777 ( .A(n_546), .Y(n_777) );
BUFx2_ASAP7_75t_L g1120 ( .A(n_546), .Y(n_1120) );
BUFx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx2_ASAP7_75t_SL g589 ( .A(n_549), .Y(n_589) );
BUFx2_ASAP7_75t_SL g656 ( .A(n_549), .Y(n_656) );
BUFx6f_ASAP7_75t_L g778 ( .A(n_549), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_557), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B1(n_554), .B2(n_556), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_553), .A2(n_722), .B1(n_793), .B2(n_794), .Y(n_792) );
OAI221xp5_ASAP7_75t_SL g970 ( .A1(n_553), .A2(n_971), .B1(n_972), .B2(n_973), .C(n_974), .Y(n_970) );
OAI221xp5_ASAP7_75t_SL g1086 ( .A1(n_553), .A2(n_722), .B1(n_1087), .B2(n_1088), .C(n_1089), .Y(n_1086) );
INVxp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_562), .B2(n_563), .Y(n_557) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g603 ( .A(n_561), .Y(n_603) );
INVx4_ASAP7_75t_L g631 ( .A(n_561), .Y(n_631) );
INVx4_ASAP7_75t_L g692 ( .A(n_561), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g720 ( .A1(n_561), .A2(n_721), .B1(n_722), .B2(n_724), .C(n_725), .Y(n_720) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g662 ( .A(n_565), .Y(n_662) );
INVx2_ASAP7_75t_L g723 ( .A(n_565), .Y(n_723) );
INVx2_ASAP7_75t_L g859 ( .A(n_565), .Y(n_859) );
BUFx4f_ASAP7_75t_L g1180 ( .A(n_567), .Y(n_1180) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI22xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_604), .B1(n_605), .B2(n_640), .Y(n_570) );
INVx1_ASAP7_75t_L g640 ( .A(n_571), .Y(n_640) );
XNOR2xp5_ASAP7_75t_L g645 ( .A(n_571), .B(n_646), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_590), .C(n_597), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_581), .Y(n_573) );
OAI21xp5_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_576), .B(n_577), .Y(n_574) );
OAI222xp33_ASAP7_75t_L g1175 ( .A1(n_575), .A2(n_1176), .B1(n_1177), .B2(n_1178), .C1(n_1179), .C2(n_1181), .Y(n_1175) );
INVx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx4f_ASAP7_75t_SL g664 ( .A(n_580), .Y(n_664) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_586), .C(n_588), .Y(n_581) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g619 ( .A(n_584), .Y(n_619) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
BUFx4f_ASAP7_75t_L g820 ( .A(n_585), .Y(n_820) );
BUFx2_ASAP7_75t_L g936 ( .A(n_585), .Y(n_936) );
BUFx2_ASAP7_75t_L g1118 ( .A(n_585), .Y(n_1118) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_587), .Y(n_654) );
HB1xp67_ASAP7_75t_L g934 ( .A(n_587), .Y(n_934) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_595), .Y(n_590) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_602), .Y(n_597) );
INVx1_ASAP7_75t_L g695 ( .A(n_599), .Y(n_695) );
BUFx4f_ASAP7_75t_SL g726 ( .A(n_599), .Y(n_726) );
BUFx3_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx3_ASAP7_75t_L g633 ( .A(n_600), .Y(n_633) );
BUFx3_ASAP7_75t_L g659 ( .A(n_600), .Y(n_659) );
BUFx3_ASAP7_75t_L g757 ( .A(n_600), .Y(n_757) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g639 ( .A(n_607), .Y(n_639) );
NAND3x1_ASAP7_75t_L g607 ( .A(n_608), .B(n_620), .C(n_629), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_616), .Y(n_608) );
OAI21xp5_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_612), .B(n_613), .Y(n_609) );
OAI21xp5_ASAP7_75t_SL g893 ( .A1(n_610), .A2(n_894), .B(n_895), .Y(n_893) );
OAI221xp5_ASAP7_75t_L g1002 ( .A1(n_610), .A2(n_1003), .B1(n_1004), .B2(n_1005), .C(n_1006), .Y(n_1002) );
OAI21xp33_ASAP7_75t_L g1059 ( .A1(n_610), .A2(n_1060), .B(n_1061), .Y(n_1059) );
INVx3_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g675 ( .A(n_614), .Y(n_675) );
INVx1_ASAP7_75t_L g983 ( .A(n_614), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_625), .Y(n_620) );
INVx1_ASAP7_75t_L g971 ( .A(n_622), .Y(n_971) );
INVx1_ASAP7_75t_L g967 ( .A(n_623), .Y(n_967) );
BUFx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVxp67_ASAP7_75t_L g799 ( .A(n_624), .Y(n_799) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_634), .Y(n_629) );
INVx1_ASAP7_75t_L g1024 ( .A(n_631), .Y(n_1024) );
BUFx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx3_ASAP7_75t_L g908 ( .A(n_636), .Y(n_908) );
BUFx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g700 ( .A(n_642), .Y(n_700) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B1(n_665), .B2(n_698), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND4xp75_ASAP7_75t_L g647 ( .A(n_648), .B(n_652), .C(n_657), .D(n_663), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
AND2x2_ASAP7_75t_SL g652 ( .A(n_653), .B(n_655), .Y(n_652) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
BUFx2_ASAP7_75t_L g861 ( .A(n_659), .Y(n_861) );
INVx1_ASAP7_75t_L g1021 ( .A(n_659), .Y(n_1021) );
INVx1_ASAP7_75t_L g741 ( .A(n_664), .Y(n_741) );
INVx1_ASAP7_75t_L g698 ( .A(n_665), .Y(n_698) );
INVx1_ASAP7_75t_L g697 ( .A(n_666), .Y(n_697) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_683), .Y(n_666) );
NOR3xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_674), .C(n_680), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B1(n_671), .B2(n_672), .Y(n_668) );
OAI221xp5_ASAP7_75t_SL g808 ( .A1(n_670), .A2(n_672), .B1(n_809), .B2(n_810), .C(n_811), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g1145 ( .A1(n_672), .A2(n_999), .B1(n_1146), .B2(n_1147), .Y(n_1145) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_690), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_691), .B(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g1126 ( .A(n_703), .Y(n_1126) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_917), .B2(n_1125), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B1(n_787), .B2(n_916), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_744), .B1(n_785), .B2(n_786), .Y(n_708) );
INVx1_ASAP7_75t_L g785 ( .A(n_709), .Y(n_785) );
INVx1_ASAP7_75t_L g743 ( .A(n_711), .Y(n_743) );
OR4x1_ASAP7_75t_L g711 ( .A(n_712), .B(n_720), .C(n_727), .D(n_733), .Y(n_711) );
OAI221xp5_ASAP7_75t_SL g965 ( .A1(n_713), .A2(n_966), .B1(n_967), .B2(n_968), .C(n_969), .Y(n_965) );
INVx2_ASAP7_75t_L g1188 ( .A(n_713), .Y(n_1188) );
INVx3_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_719), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_722), .A2(n_1023), .B1(n_1024), .B2(n_1025), .Y(n_1022) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_729), .A2(n_872), .B1(n_979), .B2(n_980), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_729), .A2(n_1056), .B1(n_1057), .B2(n_1058), .Y(n_1055) );
OAI222xp33_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_738), .B1(n_739), .B2(n_740), .C1(n_741), .C2(n_742), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx3_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx4_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g1176 ( .A(n_737), .Y(n_1176) );
BUFx2_ASAP7_75t_L g780 ( .A(n_739), .Y(n_780) );
INVx4_ASAP7_75t_L g847 ( .A(n_739), .Y(n_847) );
OAI222xp33_ASAP7_75t_L g842 ( .A1(n_741), .A2(n_843), .B1(n_845), .B2(n_846), .C1(n_848), .C2(n_849), .Y(n_842) );
INVx1_ASAP7_75t_L g786 ( .A(n_744), .Y(n_786) );
XNOR2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_761), .Y(n_744) );
XOR2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_760), .Y(n_745) );
NAND4xp75_ASAP7_75t_L g746 ( .A(n_747), .B(n_751), .C(n_755), .D(n_759), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
AND2x2_ASAP7_75t_SL g751 ( .A(n_752), .B(n_753), .Y(n_751) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_758), .Y(n_755) );
INVx1_ASAP7_75t_L g1049 ( .A(n_757), .Y(n_1049) );
XOR2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_784), .Y(n_761) );
NOR4xp75_ASAP7_75t_L g762 ( .A(n_763), .B(n_767), .C(n_773), .D(n_779), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g763 ( .A(n_764), .B(n_765), .Y(n_763) );
NAND2x1_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .Y(n_767) );
INVx1_ASAP7_75t_SL g797 ( .A(n_769), .Y(n_797) );
NAND2xp5_ASAP7_75t_SL g773 ( .A(n_774), .B(n_776), .Y(n_773) );
INVx1_ASAP7_75t_SL g931 ( .A(n_778), .Y(n_931) );
OAI21xp5_ASAP7_75t_SL g779 ( .A1(n_780), .A2(n_781), .B(n_782), .Y(n_779) );
OAI21xp5_ASAP7_75t_SL g874 ( .A1(n_780), .A2(n_875), .B(n_876), .Y(n_874) );
INVx1_ASAP7_75t_SL g916 ( .A(n_787), .Y(n_916) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_834), .B1(n_914), .B2(n_915), .Y(n_787) );
INVx1_ASAP7_75t_L g915 ( .A(n_788), .Y(n_915) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_815), .B1(n_832), .B2(n_833), .Y(n_788) );
INVx1_ASAP7_75t_L g832 ( .A(n_789), .Y(n_832) );
INVx2_ASAP7_75t_SL g814 ( .A(n_790), .Y(n_814) );
AND4x1_ASAP7_75t_L g790 ( .A(n_791), .B(n_800), .C(n_807), .D(n_812), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_792), .B(n_795), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_797), .B1(n_798), .B2(n_799), .Y(n_795) );
AND2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_806), .Y(n_800) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVxp67_ASAP7_75t_L g833 ( .A(n_815), .Y(n_833) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
XOR2x2_ASAP7_75t_L g1123 ( .A(n_816), .B(n_923), .Y(n_1123) );
NAND4xp75_ASAP7_75t_L g817 ( .A(n_818), .B(n_822), .C(n_827), .D(n_831), .Y(n_817) );
AND2x2_ASAP7_75t_SL g818 ( .A(n_819), .B(n_821), .Y(n_818) );
AND2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AND2x2_ASAP7_75t_L g827 ( .A(n_828), .B(n_830), .Y(n_827) );
INVx1_ASAP7_75t_L g914 ( .A(n_834), .Y(n_914) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_864), .B1(n_865), .B2(n_913), .Y(n_834) );
INVx1_ASAP7_75t_SL g913 ( .A(n_835), .Y(n_913) );
INVx1_ASAP7_75t_L g863 ( .A(n_836), .Y(n_863) );
AND2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_850), .Y(n_836) );
NOR2xp33_ASAP7_75t_SL g837 ( .A(n_838), .B(n_842), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_844), .Y(n_843) );
OAI21xp5_ASAP7_75t_SL g1033 ( .A1(n_846), .A2(n_1034), .B(n_1035), .Y(n_1033) );
INVx2_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_856), .Y(n_850) );
NAND2xp33_ASAP7_75t_SL g856 ( .A(n_857), .B(n_860), .Y(n_856) );
INVx2_ASAP7_75t_SL g864 ( .A(n_865), .Y(n_864) );
AO22x1_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_890), .B1(n_911), .B2(n_912), .Y(n_865) );
INVx1_ASAP7_75t_L g912 ( .A(n_866), .Y(n_912) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_881), .Y(n_868) );
NOR3xp33_ASAP7_75t_L g869 ( .A(n_870), .B(n_874), .C(n_877), .Y(n_869) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_886), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_883), .B(n_884), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .Y(n_886) );
INVx3_ASAP7_75t_SL g911 ( .A(n_890), .Y(n_911) );
XOR2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_910), .Y(n_890) );
NAND2xp5_ASAP7_75t_SL g891 ( .A(n_892), .B(n_900), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_893), .B(n_896), .Y(n_892) );
NAND3xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .C(n_899), .Y(n_896) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_905), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_904), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_906), .B(n_907), .Y(n_905) );
INVx1_ASAP7_75t_L g1125 ( .A(n_917), .Y(n_1125) );
AOI22xp5_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_919), .B1(n_1075), .B2(n_1076), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_920), .A2(n_921), .B1(n_991), .B2(n_992), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
XNOR2xp5_ASAP7_75t_L g921 ( .A(n_922), .B(n_962), .Y(n_921) );
AO22x2_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_946), .B1(n_960), .B2(n_961), .Y(n_922) );
INVx2_ASAP7_75t_L g960 ( .A(n_923), .Y(n_960) );
NAND2xp5_ASAP7_75t_SL g924 ( .A(n_925), .B(n_938), .Y(n_924) );
NOR2xp33_ASAP7_75t_SL g925 ( .A(n_926), .B(n_932), .Y(n_925) );
OAI21xp5_ASAP7_75t_SL g926 ( .A1(n_927), .A2(n_928), .B(n_929), .Y(n_926) );
OAI221xp5_ASAP7_75t_L g981 ( .A1(n_927), .A2(n_982), .B1(n_983), .B2(n_984), .C(n_985), .Y(n_981) );
INVx2_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
NAND3xp33_ASAP7_75t_L g932 ( .A(n_933), .B(n_935), .C(n_937), .Y(n_932) );
NOR2x1_ASAP7_75t_L g938 ( .A(n_939), .B(n_943), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_940), .B(n_942), .Y(n_939) );
INVx1_ASAP7_75t_L g1044 ( .A(n_941), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_944), .B(n_945), .Y(n_943) );
INVx3_ASAP7_75t_SL g961 ( .A(n_946), .Y(n_961) );
XOR2x2_ASAP7_75t_L g946 ( .A(n_947), .B(n_959), .Y(n_946) );
NAND4xp75_ASAP7_75t_L g947 ( .A(n_948), .B(n_951), .C(n_955), .D(n_958), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_949), .B(n_950), .Y(n_948) );
AND2x2_ASAP7_75t_L g955 ( .A(n_956), .B(n_957), .Y(n_955) );
INVx2_ASAP7_75t_L g990 ( .A(n_963), .Y(n_990) );
AND2x2_ASAP7_75t_SL g963 ( .A(n_964), .B(n_977), .Y(n_963) );
NOR2xp33_ASAP7_75t_L g964 ( .A(n_965), .B(n_970), .Y(n_964) );
HB1xp67_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
NOR3xp33_ASAP7_75t_L g977 ( .A(n_978), .B(n_981), .C(n_986), .Y(n_977) );
INVx1_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
AOI22xp5_ASAP7_75t_L g992 ( .A1(n_993), .A2(n_994), .B1(n_1028), .B2(n_1029), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g1027 ( .A(n_995), .Y(n_1027) );
AND3x1_ASAP7_75t_L g995 ( .A(n_996), .B(n_1011), .C(n_1019), .Y(n_995) );
NOR3xp33_ASAP7_75t_L g996 ( .A(n_997), .B(n_1002), .C(n_1007), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_999), .B1(n_1000), .B2(n_1001), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g1152 ( .A1(n_1010), .A2(n_1064), .B1(n_1153), .B2(n_1154), .Y(n_1152) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1014), .B1(n_1016), .B2(n_1017), .Y(n_1012) );
BUFx2_ASAP7_75t_R g1014 ( .A(n_1015), .Y(n_1014) );
CKINVDCx20_ASAP7_75t_R g1017 ( .A(n_1018), .Y(n_1017) );
INVx2_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx2_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_1030), .A2(n_1051), .B1(n_1052), .B2(n_1074), .Y(n_1029) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1030), .Y(n_1074) );
NAND3x2_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1041), .C(n_1046), .Y(n_1031) );
NOR2x1_ASAP7_75t_SL g1032 ( .A(n_1033), .B(n_1036), .Y(n_1032) );
NAND3xp33_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1038), .C(n_1040), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1045), .Y(n_1041) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1050), .Y(n_1046) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
INVx2_ASAP7_75t_SL g1051 ( .A(n_1052), .Y(n_1051) );
XOR2x2_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1073), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1066), .Y(n_1053) );
NOR3xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1059), .C(n_1062), .Y(n_1054) );
NOR2xp33_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1070), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1069), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1072), .Y(n_1070) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
AOI22xp5_ASAP7_75t_L g1076 ( .A1(n_1077), .A2(n_1078), .B1(n_1103), .B2(n_1124), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1079), .Y(n_1102) );
AND2x2_ASAP7_75t_SL g1079 ( .A(n_1080), .B(n_1090), .Y(n_1079) );
NOR2xp33_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1086), .Y(n_1080) );
NOR3xp33_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1094), .C(n_1098), .Y(n_1090) );
INVx2_ASAP7_75t_L g1124 ( .A(n_1103), .Y(n_1124) );
XNOR2x1_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1123), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_SL g1106 ( .A(n_1107), .Y(n_1106) );
NAND4xp75_ASAP7_75t_SL g1107 ( .A(n_1108), .B(n_1111), .C(n_1116), .D(n_1121), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1110), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1115), .Y(n_1111) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
AND2x2_ASAP7_75t_SL g1116 ( .A(n_1117), .B(n_1119), .Y(n_1116) );
INVx1_ASAP7_75t_SL g1128 ( .A(n_1129), .Y(n_1128) );
NOR2x1_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1134), .Y(n_1129) );
OR2x2_ASAP7_75t_SL g1197 ( .A(n_1130), .B(n_1135), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1133), .Y(n_1130) );
CKINVDCx20_ASAP7_75t_R g1165 ( .A(n_1131), .Y(n_1165) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1132), .B(n_1167), .Y(n_1170) );
CKINVDCx16_ASAP7_75t_R g1167 ( .A(n_1133), .Y(n_1167) );
CKINVDCx20_ASAP7_75t_R g1134 ( .A(n_1135), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1137), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1140), .Y(n_1138) );
OAI322xp33_ASAP7_75t_L g1141 ( .A1(n_1142), .A2(n_1164), .A3(n_1166), .B1(n_1168), .B2(n_1171), .C1(n_1172), .C2(n_1195), .Y(n_1141) );
INVx1_ASAP7_75t_SL g1163 ( .A(n_1143), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1155), .Y(n_1143) );
NOR3xp33_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1148), .C(n_1152), .Y(n_1144) );
NOR2xp33_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1159), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1158), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1161), .Y(n_1159) );
BUFx2_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
CKINVDCx20_ASAP7_75t_R g1168 ( .A(n_1169), .Y(n_1168) );
INVx1_ASAP7_75t_SL g1194 ( .A(n_1173), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1185), .Y(n_1173) );
NOR2x1_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1182), .Y(n_1174) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1184), .Y(n_1182) );
NOR2xp33_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1191), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1189), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1193), .Y(n_1191) );
CKINVDCx20_ASAP7_75t_R g1195 ( .A(n_1196), .Y(n_1195) );
CKINVDCx20_ASAP7_75t_R g1196 ( .A(n_1197), .Y(n_1196) );
endmodule