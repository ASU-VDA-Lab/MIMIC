module fake_jpeg_6233_n_290 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_43),
.B(n_60),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_0),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_48),
.Y(n_72)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_25),
.B(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_53),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_58),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_57),
.B(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_61),
.Y(n_100)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_34),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_1),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_70),
.A2(n_82),
.B1(n_21),
.B2(n_3),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_39),
.B1(n_36),
.B2(n_35),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_71),
.A2(n_33),
.B1(n_37),
.B2(n_35),
.Y(n_124)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_77),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_76),
.B(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_54),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_81),
.A2(n_1),
.B(n_4),
.Y(n_136)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_90),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_97),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_61),
.B1(n_56),
.B2(n_49),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_88),
.B1(n_74),
.B2(n_93),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_38),
.B1(n_26),
.B2(n_22),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_94),
.Y(n_139)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_96),
.Y(n_140)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_42),
.B(n_28),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_98),
.B(n_102),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

BUFx16f_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_24),
.Y(n_105)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_37),
.Y(n_106)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_41),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_121),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_126),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_98),
.B(n_41),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_117),
.B(n_132),
.C(n_138),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_129),
.B1(n_74),
.B2(n_93),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_32),
.C(n_29),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_116),
.A2(n_80),
.B(n_79),
.Y(n_171)
);

OR2x2_ASAP7_75t_SL g117 ( 
.A(n_88),
.B(n_16),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_88),
.A2(n_39),
.B1(n_33),
.B2(n_29),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_101),
.B1(n_92),
.B2(n_96),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_41),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_124),
.A2(n_130),
.B1(n_83),
.B2(n_107),
.Y(n_155)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_38),
.B1(n_26),
.B2(n_22),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_142),
.B1(n_75),
.B2(n_87),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_69),
.A2(n_38),
.B1(n_26),
.B2(n_22),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_17),
.C(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_94),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_121),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_99),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_78),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_136),
.A2(n_66),
.B(n_7),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_70),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_86),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_104),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_144),
.B(n_123),
.C(n_118),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_150),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_149),
.B1(n_154),
.B2(n_155),
.Y(n_178)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_142),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_152),
.B(n_160),
.Y(n_177)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_163),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_100),
.B1(n_89),
.B2(n_72),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_159),
.A2(n_167),
.B1(n_168),
.B2(n_143),
.Y(n_200)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_161),
.B(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_82),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_109),
.B(n_131),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_174),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_128),
.A2(n_95),
.B1(n_104),
.B2(n_102),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_128),
.A2(n_90),
.B1(n_68),
.B2(n_103),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_134),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_170),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_176),
.B1(n_142),
.B2(n_110),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_116),
.B(n_110),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_131),
.B(n_6),
.Y(n_173)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_80),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_150),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_66),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_142),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_190),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_200),
.B1(n_154),
.B2(n_168),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_185),
.A2(n_186),
.B(n_203),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_144),
.A2(n_113),
.B(n_79),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_188),
.Y(n_224)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_144),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_195),
.Y(n_209)
);

AO22x2_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_117),
.B1(n_138),
.B2(n_123),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_193),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_211)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_135),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_9),
.Y(n_220)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_201),
.B(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_13),
.Y(n_226)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_149),
.B1(n_175),
.B2(n_176),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_211),
.B1(n_225),
.B2(n_181),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_172),
.B(n_157),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_174),
.B(n_171),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_213),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_217),
.B1(n_218),
.B2(n_221),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_167),
.B(n_163),
.Y(n_213)
);

OA21x2_ASAP7_75t_SL g214 ( 
.A1(n_193),
.A2(n_153),
.B(n_118),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_197),
.B(n_196),
.Y(n_233)
);

OAI211xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_215),
.B(n_216),
.Y(n_238)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_165),
.B1(n_119),
.B2(n_111),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_119),
.B1(n_111),
.B2(n_125),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_219),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_223),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_221)
);

NAND2x1p5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_180),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_193),
.A2(n_10),
.B1(n_13),
.B2(n_15),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_199),
.C(n_190),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_231),
.C(n_241),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_195),
.C(n_201),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_237),
.Y(n_249)
);

BUFx12f_ASAP7_75t_SL g250 ( 
.A(n_233),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_204),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_209),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_240),
.A2(n_223),
.B1(n_210),
.B2(n_214),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_203),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_177),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_245),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_179),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_247),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_244),
.B(n_194),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_223),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_245),
.B(n_181),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_234),
.Y(n_258)
);

OAI22x1_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_221),
.B1(n_225),
.B2(n_213),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_253),
.A2(n_242),
.B1(n_239),
.B2(n_228),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_211),
.B1(n_227),
.B2(n_207),
.Y(n_254)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

NOR3xp33_ASAP7_75t_SL g257 ( 
.A(n_250),
.B(n_253),
.C(n_240),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_257),
.A2(n_258),
.B(n_261),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_262),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_232),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_236),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_230),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_267),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_264),
.A2(n_265),
.B1(n_254),
.B2(n_256),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_241),
.C(n_231),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_220),
.C(n_252),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_242),
.B(n_237),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_236),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_270),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_260),
.B(n_266),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_249),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_217),
.B1(n_218),
.B2(n_252),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_272),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_185),
.C(n_238),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_278),
.B(n_279),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_229),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_184),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_275),
.C(n_273),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_224),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_283),
.B(n_285),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_SL g284 ( 
.A(n_276),
.B(n_274),
.Y(n_284)
);

AOI21x1_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_282),
.B(n_277),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_277),
.C(n_281),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_288),
.B(n_273),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_287),
.Y(n_290)
);


endmodule