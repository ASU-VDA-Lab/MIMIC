module fake_jpeg_1944_n_710 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_710);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_710;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g142 ( 
.A(n_60),
.B(n_105),
.Y(n_142)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_61),
.Y(n_201)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_63),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_64),
.B(n_108),
.Y(n_182)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_65),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_69),
.A2(n_89),
.B1(n_45),
.B2(n_30),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_71),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_74),
.Y(n_217)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_76),
.Y(n_173)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_77),
.Y(n_180)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_79),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_80),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_10),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_81),
.B(n_82),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_27),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_83),
.Y(n_212)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_85),
.Y(n_196)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_86),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_87),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_88),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_32),
.A2(n_28),
.B1(n_47),
.B2(n_37),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_90),
.Y(n_231)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_91),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_92),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_34),
.Y(n_93)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_96),
.Y(n_220)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_97),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx6_ASAP7_75t_SL g101 ( 
.A(n_21),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g181 ( 
.A(n_101),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

BUFx12f_ASAP7_75t_SL g105 ( 
.A(n_21),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_107),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_33),
.B(n_10),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_33),
.B(n_12),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_110),
.B(n_123),
.Y(n_225)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_40),
.Y(n_112)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_112),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_113),
.Y(n_219)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_122),
.Y(n_150)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_22),
.Y(n_118)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_118),
.Y(n_171)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_22),
.Y(n_120)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_39),
.Y(n_121)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_25),
.B(n_12),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_26),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_58),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_22),
.Y(n_125)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_59),
.Y(n_127)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_49),
.Y(n_129)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_40),
.Y(n_131)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_40),
.Y(n_132)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_SL g133 ( 
.A(n_60),
.Y(n_133)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_133),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_81),
.B(n_25),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_139),
.B(n_174),
.Y(n_262)
);

BUFx8_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

CKINVDCx6p67_ASAP7_75t_R g283 ( 
.A(n_148),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_131),
.A2(n_45),
.B1(n_39),
.B2(n_38),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_151),
.A2(n_125),
.B1(n_72),
.B2(n_76),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_152),
.B(n_163),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_31),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_165),
.A2(n_70),
.B1(n_5),
.B2(n_6),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_93),
.B(n_38),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_117),
.B(n_50),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_175),
.B(n_183),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_127),
.A2(n_49),
.B1(n_36),
.B2(n_54),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_177),
.A2(n_188),
.B1(n_192),
.B2(n_199),
.Y(n_236)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_75),
.Y(n_178)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_179),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_31),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_69),
.B(n_58),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_184),
.B(n_187),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_61),
.B(n_57),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_102),
.A2(n_20),
.B1(n_54),
.B2(n_53),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_102),
.A2(n_42),
.B1(n_53),
.B2(n_51),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_193),
.Y(n_258)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_80),
.A2(n_42),
.B1(n_51),
.B2(n_36),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_65),
.A2(n_20),
.B1(n_43),
.B2(n_35),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_200),
.A2(n_216),
.B1(n_84),
.B2(n_73),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_120),
.B(n_50),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_206),
.B(n_215),
.Y(n_292)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_85),
.Y(n_207)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_207),
.Y(n_277)
);

INVx6_ASAP7_75t_SL g210 ( 
.A(n_86),
.Y(n_210)
);

BUFx4f_ASAP7_75t_SL g295 ( 
.A(n_210),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_91),
.B(n_57),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_74),
.A2(n_43),
.B1(n_35),
.B2(n_26),
.Y(n_216)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_87),
.Y(n_221)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_221),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_129),
.B(n_12),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_222),
.B(n_224),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_106),
.B(n_9),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_107),
.Y(n_226)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_111),
.B(n_19),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_227),
.B(n_228),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_126),
.B(n_9),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_88),
.B(n_18),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_0),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_232),
.B(n_241),
.Y(n_341)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_234),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_128),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_235),
.B(n_290),
.C(n_218),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_134),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_237),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_141),
.B(n_116),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_238),
.B(n_242),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_148),
.Y(n_240)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_240),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_150),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_0),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_154),
.Y(n_244)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_244),
.Y(n_342)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_134),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_245),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_140),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_246),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_247),
.A2(n_300),
.B1(n_159),
.B2(n_173),
.Y(n_360)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_181),
.Y(n_249)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_249),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_250),
.A2(n_259),
.B1(n_272),
.B2(n_312),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_3),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_251),
.B(n_254),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_153),
.Y(n_252)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_252),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_137),
.B(n_4),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_170),
.Y(n_255)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_255),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_140),
.Y(n_256)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_256),
.Y(n_349)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_154),
.Y(n_257)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_257),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_142),
.A2(n_68),
.B1(n_67),
.B2(n_66),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_133),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_260),
.B(n_268),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_138),
.B(n_4),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_261),
.B(n_267),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_264),
.A2(n_265),
.B1(n_302),
.B2(n_303),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_184),
.A2(n_13),
.B1(n_17),
.B2(n_16),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_143),
.Y(n_266)
);

INVx8_ASAP7_75t_L g378 ( 
.A(n_266),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_145),
.B(n_4),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_187),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_167),
.Y(n_269)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_269),
.Y(n_337)
);

INVx3_ASAP7_75t_SL g270 ( 
.A(n_160),
.Y(n_270)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_270),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_166),
.B(n_4),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_271),
.B(n_288),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_191),
.A2(n_13),
.B1(n_17),
.B2(n_16),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_199),
.A2(n_162),
.B1(n_157),
.B2(n_214),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_273),
.A2(n_176),
.B1(n_223),
.B2(n_196),
.Y(n_317)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_201),
.Y(n_274)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_274),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_202),
.A2(n_13),
.B1(n_16),
.B2(n_15),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_275),
.A2(n_197),
.B(n_185),
.Y(n_351)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_160),
.B(n_4),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_276),
.Y(n_352)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_170),
.Y(n_279)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_279),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_208),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_280),
.B(n_293),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_201),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_281),
.B(n_285),
.Y(n_344)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_143),
.Y(n_282)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_282),
.Y(n_338)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_144),
.Y(n_284)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_284),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_169),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_231),
.Y(n_286)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_286),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_186),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_287),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_188),
.B(n_5),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_212),
.B(n_14),
.C(n_15),
.Y(n_290)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_149),
.Y(n_293)
);

INVx11_ASAP7_75t_L g296 ( 
.A(n_147),
.Y(n_296)
);

BUFx12f_ASAP7_75t_L g318 ( 
.A(n_296),
.Y(n_318)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_149),
.Y(n_297)
);

INVx13_ASAP7_75t_L g372 ( 
.A(n_297),
.Y(n_372)
);

INVx3_ASAP7_75t_SL g298 ( 
.A(n_219),
.Y(n_298)
);

CKINVDCx10_ASAP7_75t_R g333 ( 
.A(n_298),
.Y(n_333)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_213),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_299),
.B(n_305),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_192),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_177),
.A2(n_18),
.B1(n_7),
.B2(n_8),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_L g303 ( 
.A1(n_200),
.A2(n_216),
.B1(n_194),
.B2(n_155),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_162),
.B(n_6),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_304),
.B(n_306),
.Y(n_331)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_164),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_205),
.B(n_6),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_168),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_308),
.Y(n_359)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_168),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_203),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_309),
.B(n_310),
.Y(n_361)
);

INVx3_ASAP7_75t_SL g310 ( 
.A(n_198),
.Y(n_310)
);

INVx11_ASAP7_75t_L g312 ( 
.A(n_147),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_203),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_313),
.B(n_314),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_217),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_208),
.A2(n_146),
.B(n_211),
.C(n_198),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_L g353 ( 
.A1(n_315),
.A2(n_180),
.B(n_147),
.C(n_230),
.Y(n_353)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_217),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_316),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_317),
.A2(n_366),
.B1(n_368),
.B2(n_291),
.Y(n_399)
);

AND2x2_ASAP7_75t_SL g320 ( 
.A(n_238),
.B(n_156),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_320),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_264),
.A2(n_136),
.B1(n_135),
.B2(n_155),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_321),
.A2(n_355),
.B1(n_366),
.B2(n_368),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_329),
.B(n_283),
.Y(n_404)
);

OA22x2_ASAP7_75t_L g330 ( 
.A1(n_273),
.A2(n_194),
.B1(n_135),
.B2(n_136),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_330),
.B(n_284),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_235),
.B(n_230),
.C(n_146),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_334),
.B(n_240),
.C(n_280),
.Y(n_386)
);

OAI21xp33_ASAP7_75t_L g340 ( 
.A1(n_268),
.A2(n_18),
.B(n_146),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_340),
.B(n_370),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_288),
.A2(n_236),
.B(n_315),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_345),
.A2(n_351),
.B(n_325),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_289),
.A2(n_176),
.B1(n_223),
.B2(n_214),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_347),
.A2(n_283),
.B1(n_255),
.B2(n_260),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_303),
.A2(n_157),
.B1(n_196),
.B2(n_159),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_348),
.A2(n_364),
.B1(n_317),
.B2(n_321),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_262),
.B(n_161),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_350),
.B(n_376),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_351),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_353),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_276),
.A2(n_242),
.B1(n_294),
.B2(n_304),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_360),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_306),
.A2(n_173),
.B1(n_144),
.B2(n_158),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_301),
.A2(n_158),
.B1(n_209),
.B2(n_171),
.Y(n_366)
);

O2A1O1Ixp33_ASAP7_75t_SL g367 ( 
.A1(n_276),
.A2(n_171),
.B(n_204),
.C(n_190),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_367),
.A2(n_375),
.B1(n_283),
.B2(n_240),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_232),
.A2(n_209),
.B1(n_204),
.B2(n_190),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_249),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_278),
.A2(n_190),
.B1(n_7),
.B2(n_8),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_251),
.B(n_6),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_261),
.A2(n_7),
.B1(n_8),
.B2(n_267),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_377),
.A2(n_255),
.B1(n_277),
.B2(n_311),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_331),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_380),
.B(n_382),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_345),
.A2(n_254),
.B1(n_271),
.B2(n_292),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_381),
.A2(n_384),
.B1(n_390),
.B2(n_397),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_239),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_325),
.A2(n_275),
.B1(n_282),
.B2(n_245),
.Y(n_384)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_378),
.Y(n_385)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_385),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_386),
.B(n_404),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_388),
.A2(n_402),
.B(n_408),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_371),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_392),
.B(n_422),
.Y(n_462)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_369),
.Y(n_393)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_393),
.Y(n_430)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_365),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_394),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_395),
.Y(n_444)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_396),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_352),
.A2(n_253),
.B1(n_258),
.B2(n_248),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_370),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_398),
.B(n_410),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_399),
.A2(n_343),
.B1(n_330),
.B2(n_362),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_331),
.B(n_290),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_400),
.B(n_407),
.Y(n_452)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_363),
.Y(n_403)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_403),
.Y(n_435)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_363),
.Y(n_406)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_406),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_322),
.B(n_295),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_367),
.A2(n_233),
.B1(n_283),
.B2(n_312),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_322),
.B(n_358),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_409),
.B(n_412),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_336),
.B(n_269),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_336),
.B(n_285),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_411),
.B(n_426),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_358),
.B(n_295),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_365),
.Y(n_413)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_413),
.Y(n_450)
);

OAI22xp33_ASAP7_75t_L g471 ( 
.A1(n_414),
.A2(n_233),
.B1(n_296),
.B2(n_333),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_348),
.A2(n_327),
.B1(n_360),
.B2(n_329),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_415),
.A2(n_419),
.B1(n_425),
.B2(n_353),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_334),
.B(n_263),
.C(n_243),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_416),
.B(n_429),
.Y(n_448)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_339),
.Y(n_417)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_417),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_327),
.A2(n_266),
.B1(n_256),
.B2(n_237),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_355),
.B(n_295),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_420),
.B(n_421),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_243),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_354),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_342),
.Y(n_423)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_423),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_424),
.B(n_428),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_356),
.A2(n_246),
.B1(n_258),
.B2(n_253),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_326),
.B(n_252),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_427),
.B(n_323),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_352),
.B(n_248),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_320),
.B(n_263),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_438),
.A2(n_451),
.B1(n_456),
.B2(n_458),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_426),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_440),
.B(n_442),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_410),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_389),
.A2(n_320),
.B1(n_364),
.B2(n_367),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_445),
.A2(n_464),
.B1(n_419),
.B2(n_421),
.Y(n_496)
);

OA21x2_ASAP7_75t_L g447 ( 
.A1(n_395),
.A2(n_330),
.B(n_344),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_468),
.Y(n_478)
);

AOI32xp33_ASAP7_75t_L g449 ( 
.A1(n_391),
.A2(n_332),
.A3(n_361),
.B1(n_343),
.B2(n_333),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_449),
.B(n_401),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_389),
.A2(n_341),
.B1(n_328),
.B2(n_319),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_454),
.A2(n_455),
.B(n_466),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_388),
.A2(n_328),
.B(n_319),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_415),
.A2(n_330),
.B1(n_326),
.B2(n_376),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_398),
.Y(n_457)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_457),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_384),
.A2(n_362),
.B1(n_338),
.B2(n_335),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_418),
.A2(n_338),
.B1(n_335),
.B2(n_374),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_459),
.A2(n_349),
.B1(n_337),
.B2(n_378),
.Y(n_502)
);

OA22x2_ASAP7_75t_L g461 ( 
.A1(n_399),
.A2(n_374),
.B1(n_342),
.B2(n_323),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_461),
.B(n_451),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_418),
.A2(n_335),
.B1(n_349),
.B2(n_277),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_387),
.A2(n_354),
.B(n_357),
.Y(n_466)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_467),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_411),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_412),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_380),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_471),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_463),
.B(n_404),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_472),
.B(n_453),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_463),
.B(n_404),
.C(n_416),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_473),
.B(n_476),
.C(n_483),
.Y(n_514)
);

AOI32xp33_ASAP7_75t_L g474 ( 
.A1(n_470),
.A2(n_387),
.A3(n_420),
.B1(n_407),
.B2(n_392),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_474),
.B(n_509),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_386),
.C(n_409),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_455),
.A2(n_402),
.B(n_401),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_477),
.A2(n_480),
.B(n_466),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_481),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_432),
.A2(n_408),
.B(n_395),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_482),
.A2(n_493),
.B(n_495),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_448),
.B(n_429),
.C(n_428),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_438),
.A2(n_383),
.B1(n_390),
.B2(n_395),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_484),
.A2(n_458),
.B1(n_433),
.B2(n_459),
.Y(n_534)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_430),
.Y(n_486)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_486),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_436),
.A2(n_383),
.B1(n_400),
.B2(n_382),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_487),
.A2(n_496),
.B1(n_443),
.B2(n_460),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_457),
.B(n_405),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_488),
.B(n_506),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_452),
.B(n_381),
.C(n_397),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_489),
.B(n_494),
.C(n_503),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_467),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_490),
.A2(n_502),
.B1(n_505),
.B2(n_507),
.Y(n_530)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_446),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_491),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_432),
.A2(n_425),
.B(n_396),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_452),
.B(n_423),
.C(n_403),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_449),
.A2(n_393),
.B(n_406),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_445),
.A2(n_405),
.B1(n_424),
.B2(n_413),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_497),
.A2(n_498),
.B1(n_500),
.B2(n_469),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_436),
.A2(n_385),
.B1(n_414),
.B2(n_394),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_430),
.Y(n_499)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_499),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_456),
.A2(n_385),
.B1(n_417),
.B2(n_427),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_431),
.Y(n_501)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_501),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_453),
.B(n_359),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_431),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_441),
.B(n_379),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_433),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_435),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_508),
.B(n_511),
.Y(n_524)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_446),
.Y(n_509)
);

AOI21x1_ASAP7_75t_L g515 ( 
.A1(n_495),
.A2(n_477),
.B(n_478),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_515),
.A2(n_527),
.B(n_547),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_516),
.A2(n_521),
.B1(n_523),
.B2(n_531),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_479),
.Y(n_517)
);

INVx13_ASAP7_75t_L g572 ( 
.A(n_517),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_519),
.B(n_522),
.C(n_543),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_473),
.B(n_441),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_520),
.B(n_483),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_484),
.A2(n_444),
.B1(n_447),
.B2(n_468),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_476),
.B(n_454),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_492),
.A2(n_444),
.B1(n_447),
.B2(n_443),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_507),
.B(n_434),
.Y(n_525)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_525),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_489),
.B(n_462),
.Y(n_526)
);

CKINVDCx14_ASAP7_75t_R g560 ( 
.A(n_526),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_479),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_528),
.B(n_539),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_487),
.A2(n_444),
.B1(n_447),
.B2(n_460),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_511),
.A2(n_444),
.B1(n_440),
.B2(n_442),
.Y(n_532)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_532),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_481),
.B(n_462),
.Y(n_533)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_533),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_534),
.A2(n_537),
.B1(n_544),
.B2(n_510),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_478),
.A2(n_464),
.B1(n_434),
.B2(n_435),
.Y(n_535)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_535),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_482),
.A2(n_437),
.B1(n_469),
.B2(n_461),
.Y(n_538)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_538),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_479),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_494),
.B(n_437),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_540),
.B(n_541),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_490),
.B(n_485),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_493),
.A2(n_461),
.B1(n_450),
.B2(n_465),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_542),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_472),
.B(n_450),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_497),
.A2(n_496),
.B1(n_498),
.B2(n_500),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_503),
.B(n_379),
.Y(n_548)
);

CKINVDCx14_ASAP7_75t_R g564 ( 
.A(n_548),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_485),
.B(n_461),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_549),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_546),
.B(n_474),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g608 ( 
.A(n_553),
.Y(n_608)
);

CKINVDCx16_ASAP7_75t_R g557 ( 
.A(n_541),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_557),
.B(n_563),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_546),
.B(n_512),
.Y(n_558)
);

CKINVDCx16_ASAP7_75t_R g611 ( 
.A(n_558),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_559),
.B(n_578),
.Y(n_587)
);

A2O1A1Ixp33_ASAP7_75t_SL g561 ( 
.A1(n_549),
.A2(n_504),
.B(n_510),
.C(n_475),
.Y(n_561)
);

A2O1A1Ixp33_ASAP7_75t_L g599 ( 
.A1(n_561),
.A2(n_524),
.B(n_513),
.C(n_544),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_525),
.Y(n_563)
);

BUFx24_ASAP7_75t_SL g565 ( 
.A(n_520),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_565),
.B(n_297),
.Y(n_610)
);

INVx2_ASAP7_75t_R g568 ( 
.A(n_517),
.Y(n_568)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_568),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_514),
.B(n_475),
.C(n_504),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_569),
.B(n_573),
.C(n_576),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_570),
.A2(n_521),
.B(n_532),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_518),
.B(n_337),
.Y(n_571)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_571),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_514),
.B(n_508),
.C(n_505),
.Y(n_573)
);

CKINVDCx14_ASAP7_75t_R g574 ( 
.A(n_533),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_574),
.A2(n_513),
.B1(n_530),
.B2(n_535),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_575),
.A2(n_550),
.B1(n_545),
.B2(n_529),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_522),
.B(n_499),
.C(n_486),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_519),
.B(n_543),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_540),
.B(n_527),
.C(n_539),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_579),
.B(n_580),
.C(n_515),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_528),
.B(n_501),
.C(n_465),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_516),
.B(n_461),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_582),
.B(n_583),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_531),
.B(n_354),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_536),
.Y(n_585)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_585),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_SL g589 ( 
.A(n_578),
.B(n_547),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_SL g628 ( 
.A(n_589),
.B(n_602),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_590),
.B(n_612),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_SL g625 ( 
.A1(n_591),
.A2(n_566),
.B(n_552),
.Y(n_625)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_593),
.Y(n_615)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_585),
.Y(n_595)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_595),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_559),
.B(n_523),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g637 ( 
.A(n_596),
.B(n_607),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_573),
.B(n_538),
.C(n_537),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_597),
.B(n_603),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_599),
.B(n_606),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_577),
.B(n_524),
.Y(n_601)
);

CKINVDCx14_ASAP7_75t_R g632 ( 
.A(n_601),
.Y(n_632)
);

XNOR2x1_ASAP7_75t_L g602 ( 
.A(n_579),
.B(n_542),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_569),
.B(n_534),
.C(n_545),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_567),
.B(n_550),
.C(n_536),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_604),
.B(n_551),
.C(n_556),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_605),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_555),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_567),
.B(n_529),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_SL g609 ( 
.A(n_576),
.B(n_491),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_SL g635 ( 
.A(n_609),
.B(n_554),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_610),
.B(n_580),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_570),
.B(n_555),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_584),
.A2(n_509),
.B1(n_439),
.B2(n_346),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g618 ( 
.A1(n_613),
.A2(n_566),
.B1(n_581),
.B2(n_551),
.Y(n_618)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_614),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_611),
.B(n_560),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_616),
.B(n_620),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_618),
.A2(n_346),
.B1(n_324),
.B2(n_293),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_608),
.B(n_564),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_604),
.B(n_554),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_621),
.A2(n_630),
.B(n_311),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_623),
.B(n_624),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_607),
.B(n_584),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_625),
.A2(n_561),
.B(n_605),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_587),
.B(n_556),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_L g650 ( 
.A(n_626),
.B(n_600),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_586),
.B(n_587),
.C(n_596),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_627),
.B(n_629),
.C(n_633),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_586),
.B(n_552),
.C(n_581),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_591),
.A2(n_562),
.B(n_568),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_603),
.B(n_583),
.C(n_582),
.Y(n_633)
);

MAJx2_ASAP7_75t_L g639 ( 
.A(n_635),
.B(n_589),
.C(n_590),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_588),
.B(n_561),
.Y(n_636)
);

OAI321xp33_ASAP7_75t_L g644 ( 
.A1(n_636),
.A2(n_572),
.A3(n_561),
.B1(n_598),
.B2(n_602),
.C(n_594),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_SL g638 ( 
.A1(n_615),
.A2(n_592),
.B1(n_601),
.B2(n_599),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_638),
.A2(n_644),
.B1(n_647),
.B2(n_651),
.Y(n_668)
);

XOR2xp5_ASAP7_75t_L g659 ( 
.A(n_639),
.B(n_650),
.Y(n_659)
);

XOR2xp5_ASAP7_75t_L g640 ( 
.A(n_637),
.B(n_597),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_L g665 ( 
.A(n_640),
.B(n_645),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_642),
.B(n_649),
.Y(n_660)
);

XOR2xp5_ASAP7_75t_L g645 ( 
.A(n_637),
.B(n_609),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_SL g647 ( 
.A1(n_632),
.A2(n_634),
.B1(n_613),
.B2(n_617),
.Y(n_647)
);

FAx1_ASAP7_75t_SL g649 ( 
.A(n_629),
.B(n_612),
.CI(n_572),
.CON(n_649),
.SN(n_649)
);

OAI22xp5_ASAP7_75t_SL g651 ( 
.A1(n_617),
.A2(n_598),
.B1(n_600),
.B2(n_439),
.Y(n_651)
);

MAJx2_ASAP7_75t_L g652 ( 
.A(n_628),
.B(n_439),
.C(n_324),
.Y(n_652)
);

FAx1_ASAP7_75t_SL g674 ( 
.A(n_652),
.B(n_318),
.CI(n_372),
.CON(n_674),
.SN(n_674)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_627),
.B(n_439),
.C(n_346),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_653),
.B(n_656),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g654 ( 
.A(n_624),
.B(n_274),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g669 ( 
.A(n_654),
.B(n_635),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_SL g670 ( 
.A1(n_655),
.A2(n_631),
.B1(n_652),
.B2(n_649),
.Y(n_670)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_622),
.B(n_324),
.C(n_270),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_657),
.B(n_653),
.Y(n_671)
);

AO21x1_ASAP7_75t_L g658 ( 
.A1(n_642),
.A2(n_630),
.B(n_636),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_658),
.B(n_674),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_SL g661 ( 
.A(n_646),
.B(n_619),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_661),
.Y(n_679)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_648),
.B(n_623),
.C(n_619),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_662),
.B(n_663),
.C(n_666),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_648),
.B(n_633),
.C(n_618),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_641),
.Y(n_664)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_664),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_641),
.B(n_626),
.C(n_625),
.Y(n_666)
);

XNOR2xp5_ASAP7_75t_L g683 ( 
.A(n_669),
.B(n_671),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_670),
.A2(n_673),
.B1(n_638),
.B2(n_654),
.Y(n_676)
);

NOR2xp67_ASAP7_75t_SL g672 ( 
.A(n_640),
.B(n_628),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_672),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_643),
.B(n_318),
.Y(n_673)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_676),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_660),
.A2(n_649),
.B(n_639),
.Y(n_678)
);

AOI21xp33_ASAP7_75t_L g693 ( 
.A1(n_678),
.A2(n_680),
.B(n_659),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_SL g680 ( 
.A1(n_660),
.A2(n_655),
.B(n_645),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_668),
.A2(n_657),
.B1(n_650),
.B2(n_310),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_684),
.B(n_685),
.Y(n_688)
);

MAJIxp5_ASAP7_75t_L g685 ( 
.A(n_662),
.B(n_298),
.C(n_372),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_663),
.B(n_666),
.Y(n_686)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_686),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_681),
.A2(n_682),
.B(n_658),
.Y(n_689)
);

AO21x1_ASAP7_75t_L g696 ( 
.A1(n_689),
.A2(n_681),
.B(n_679),
.Y(n_696)
);

CKINVDCx16_ASAP7_75t_R g690 ( 
.A(n_682),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_690),
.A2(n_692),
.B1(n_675),
.B2(n_677),
.Y(n_697)
);

XOR2xp5_ASAP7_75t_L g691 ( 
.A(n_683),
.B(n_665),
.Y(n_691)
);

XNOR2xp5_ASAP7_75t_L g698 ( 
.A(n_691),
.B(n_694),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_677),
.B(n_667),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_693),
.A2(n_659),
.B(n_685),
.Y(n_700)
);

XOR2xp5_ASAP7_75t_L g694 ( 
.A(n_683),
.B(n_665),
.Y(n_694)
);

AOI21x1_ASAP7_75t_L g702 ( 
.A1(n_696),
.A2(n_700),
.B(n_689),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_697),
.B(n_699),
.Y(n_701)
);

MAJIxp5_ASAP7_75t_L g699 ( 
.A(n_695),
.B(n_694),
.C(n_691),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_702),
.A2(n_703),
.B(n_698),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_SL g703 ( 
.A1(n_696),
.A2(n_687),
.B(n_674),
.C(n_669),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_704),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_701),
.B(n_688),
.Y(n_705)
);

MAJIxp5_ASAP7_75t_L g707 ( 
.A(n_706),
.B(n_705),
.C(n_318),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_707),
.B(n_318),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_708),
.B(n_252),
.Y(n_709)
);

AO21x1_ASAP7_75t_L g710 ( 
.A1(n_709),
.A2(n_291),
.B(n_7),
.Y(n_710)
);


endmodule