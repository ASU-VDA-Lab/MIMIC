module real_jpeg_9000_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_244;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_2),
.A2(n_10),
.B1(n_56),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_2),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_70),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_70),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_70),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_5),
.A2(n_38),
.B(n_41),
.C(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_5),
.B(n_41),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_5),
.A2(n_9),
.B(n_25),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_6),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_6),
.A2(n_61),
.B(n_75),
.C(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_6),
.B(n_61),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_6),
.A2(n_9),
.B(n_61),
.C(n_215),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_8),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_8),
.A2(n_33),
.B1(n_61),
.B2(n_62),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_8),
.A2(n_10),
.B1(n_33),
.B2(n_56),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_9),
.A2(n_56),
.B(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_9),
.B(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_9),
.A2(n_27),
.B1(n_61),
.B2(n_62),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_9),
.A2(n_27),
.B1(n_41),
.B2(n_42),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_9),
.B(n_58),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_9),
.B(n_125),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_10),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_45),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_136),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_134),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_106),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_15),
.B(n_106),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_91),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_83),
.B2(n_84),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_50),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_20),
.B(n_36),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_29),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_21),
.B(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_22),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_23),
.A2(n_34),
.B(n_35),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_24),
.B(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_35),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_27),
.A2(n_39),
.B(n_42),
.C(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_27),
.B(n_37),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_27),
.B(n_35),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_27),
.A2(n_41),
.B(n_76),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_28),
.B(n_32),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_28),
.B(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_29),
.A2(n_35),
.B(n_94),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_30),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_34),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_34),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B(n_46),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_37),
.A2(n_88),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_38),
.B(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_38),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_38),
.B(n_98),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_40),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_46),
.B(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_48),
.B(n_187),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_71),
.B2(n_82),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_64),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_55),
.B(n_66),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_59),
.B(n_60),
.C(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_60),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_57),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_58),
.B(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_69),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_61),
.B(n_63),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_62),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_64),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_67),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_73),
.B(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_74),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_80),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_77),
.B(n_149),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_79),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_80),
.B(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_90),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_85),
.A2(n_86),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_86),
.B(n_214),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_89),
.B(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.C(n_102),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_95),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_97),
.B(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_98),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_111),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_107),
.B(n_110),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_111),
.A2(n_112),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_122),
.C(n_130),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_114),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_123),
.B1(n_130),
.B2(n_131),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_129),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_169),
.B(n_247),
.C(n_252),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_155),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_138),
.B(n_155),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_152),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_140),
.B(n_141),
.C(n_152),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_147),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_156),
.A2(n_157),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_243)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.C(n_165),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_163),
.B(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_164),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_178),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_179),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_246),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_240),
.B(n_245),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_225),
.B(n_239),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_210),
.B(n_224),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_199),
.B(n_209),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_188),
.B(n_198),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_180),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_182),
.B(n_184),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_193),
.B(n_197),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_191),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_201),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_206),
.C(n_208),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_212),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_217),
.B1(n_218),
.B2(n_223),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_213),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_214),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_219),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_222),
.C(n_223),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_226),
.B(n_227),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_232),
.B2(n_233),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_234),
.C(n_238),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_234),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_236),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_241),
.B(n_242),
.Y(n_245)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);


endmodule