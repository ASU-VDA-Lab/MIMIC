module fake_jpeg_24921_n_347 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_43),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_38),
.B(n_40),
.Y(n_79)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_45),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_0),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_24),
.Y(n_73)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_33),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_16),
.B1(n_25),
.B2(n_31),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_51),
.A2(n_35),
.B1(n_29),
.B2(n_32),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_54),
.A2(n_63),
.B1(n_68),
.B2(n_76),
.Y(n_102)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_35),
.B1(n_29),
.B2(n_32),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_71),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_32),
.B1(n_20),
.B2(n_27),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_17),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_82),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_36),
.A2(n_20),
.B1(n_18),
.B2(n_26),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_40),
.A2(n_27),
.B1(n_33),
.B2(n_31),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_33),
.B1(n_31),
.B2(n_52),
.Y(n_85)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_18),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_85),
.A2(n_72),
.B1(n_70),
.B2(n_82),
.Y(n_131)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_89),
.Y(n_128)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_91),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_18),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_96),
.C(n_113),
.Y(n_153)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_41),
.B1(n_48),
.B2(n_44),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_93),
.A2(n_103),
.B1(n_7),
.B2(n_14),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_49),
.B(n_41),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_94),
.A2(n_104),
.B(n_24),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_49),
.C(n_47),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_83),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_118),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_30),
.B1(n_42),
.B2(n_40),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_54),
.B1(n_61),
.B2(n_69),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_60),
.A2(n_16),
.B1(n_22),
.B2(n_30),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_47),
.B1(n_39),
.B2(n_42),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_121),
.B1(n_72),
.B2(n_74),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_66),
.B(n_26),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_109),
.B(n_110),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_22),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_22),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_53),
.B(n_39),
.C(n_44),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_76),
.A2(n_25),
.B1(n_43),
.B2(n_34),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_23),
.B(n_34),
.C(n_78),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_59),
.B(n_34),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_56),
.B(n_24),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_24),
.B(n_23),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_0),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_58),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_119),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_60),
.A2(n_34),
.B1(n_23),
.B2(n_10),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_145),
.B(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_127),
.B(n_130),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_SL g129 ( 
.A(n_93),
.B(n_74),
.C(n_70),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_132),
.B1(n_90),
.B2(n_89),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_104),
.B1(n_93),
.B2(n_102),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_118),
.B1(n_97),
.B2(n_100),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_138),
.A2(n_84),
.B(n_2),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_152),
.Y(n_154)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_147),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_134),
.B1(n_124),
.B2(n_151),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_93),
.B(n_0),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_97),
.A2(n_9),
.B(n_14),
.C(n_13),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_115),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_15),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_104),
.B1(n_92),
.B2(n_118),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_98),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_176),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_160),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_139),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_161),
.A2(n_172),
.B1(n_1),
.B2(n_2),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_162),
.B(n_164),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_122),
.B1(n_95),
.B2(n_111),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_163),
.A2(n_165),
.B1(n_168),
.B2(n_170),
.Y(n_215)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_166),
.B(n_169),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_122),
.B1(n_95),
.B2(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

AO21x2_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_117),
.B(n_99),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_171),
.A2(n_187),
.B1(n_125),
.B2(n_126),
.Y(n_193)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_102),
.B1(n_100),
.B2(n_92),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_175),
.B1(n_180),
.B2(n_135),
.Y(n_203)
);

OR2x2_ASAP7_75t_SL g174 ( 
.A(n_137),
.B(n_106),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_174),
.A2(n_179),
.B(n_12),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_86),
.B1(n_120),
.B2(n_114),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_101),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_87),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_181),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_91),
.Y(n_178)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_SL g179 ( 
.A(n_137),
.B(n_84),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_90),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_183),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_141),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_188),
.B(n_150),
.Y(n_191)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_4),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_146),
.A2(n_153),
.B1(n_147),
.B2(n_125),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_153),
.A2(n_1),
.B(n_2),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_171),
.A2(n_150),
.B1(n_149),
.B2(n_124),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_189),
.A2(n_190),
.B1(n_202),
.B2(n_203),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_171),
.B1(n_184),
.B2(n_156),
.Y(n_190)
);

XOR2x1_ASAP7_75t_SL g238 ( 
.A(n_191),
.B(n_162),
.Y(n_238)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_192),
.B(n_200),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_193),
.A2(n_206),
.B1(n_210),
.B2(n_161),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_126),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_194),
.B(n_197),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_136),
.C(n_130),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_127),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_199),
.B(n_217),
.Y(n_223)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_214),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_171),
.A2(n_135),
.B1(n_9),
.B2(n_11),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_1),
.B(n_2),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_204),
.A2(n_221),
.B(n_206),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_205),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_169),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_177),
.B1(n_176),
.B2(n_170),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_171),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_160),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_213),
.Y(n_228)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_181),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_216),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_154),
.B(n_9),
.Y(n_217)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_5),
.C(n_6),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_220),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_154),
.B(n_15),
.C(n_11),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_167),
.B(n_204),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_191),
.B(n_196),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_179),
.Y(n_227)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_193),
.B(n_173),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_229),
.B(n_238),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_182),
.Y(n_230)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_231),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_211),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_234),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_188),
.Y(n_235)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_203),
.A2(n_171),
.B1(n_155),
.B2(n_174),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_237),
.A2(n_250),
.B1(n_221),
.B2(n_207),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_164),
.C(n_185),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_249),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_192),
.B(n_172),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_161),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_197),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_244),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_196),
.Y(n_246)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_201),
.A2(n_222),
.B1(n_215),
.B2(n_210),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_194),
.C(n_207),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_264),
.C(n_265),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_189),
.B1(n_208),
.B2(n_195),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_254),
.A2(n_261),
.B1(n_231),
.B2(n_227),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_273),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_199),
.Y(n_263)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_263),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_220),
.C(n_219),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_217),
.C(n_230),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_233),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_238),
.B(n_237),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_246),
.Y(n_275)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_279),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_270),
.A2(n_247),
.B1(n_225),
.B2(n_226),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_270),
.B1(n_261),
.B2(n_259),
.Y(n_300)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_229),
.C(n_248),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_286),
.C(n_292),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_266),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_283),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_284),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_269),
.B(n_241),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_289),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_251),
.C(n_265),
.Y(n_286)
);

AO22x1_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_273),
.B1(n_259),
.B2(n_269),
.Y(n_301)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_290),
.Y(n_298)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_248),
.C(n_227),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_266),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_235),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_251),
.B(n_255),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_294),
.A2(n_233),
.B(n_260),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_275),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_299),
.B(n_302),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_300),
.A2(n_301),
.B1(n_262),
.B2(n_263),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_267),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_305),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_271),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_286),
.C(n_281),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_308),
.A2(n_309),
.B(n_310),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_281),
.C(n_282),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_274),
.C(n_291),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_291),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_314),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_300),
.A2(n_287),
.B1(n_258),
.B2(n_262),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_313),
.A2(n_294),
.B1(n_304),
.B2(n_305),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_228),
.C(n_234),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_315),
.B(n_293),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_285),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_320),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_228),
.C(n_264),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_292),
.C(n_224),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_298),
.B1(n_236),
.B2(n_289),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_324),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_302),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_310),
.A2(n_298),
.B1(n_295),
.B2(n_312),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_325),
.B(n_328),
.Y(n_332)
);

XOR2x2_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_323),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_334),
.Y(n_340)
);

XOR2x2_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_329),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_333),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_326),
.A2(n_308),
.B(n_309),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_321),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_335),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_325),
.Y(n_336)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_336),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_338),
.Y(n_341)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_341),
.A2(n_342),
.B(n_338),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_339),
.A2(n_331),
.B1(n_336),
.B2(n_332),
.Y(n_342)
);

AOI21x1_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_340),
.B(n_322),
.Y(n_344)
);

BUFx24_ASAP7_75t_SL g345 ( 
.A(n_344),
.Y(n_345)
);

AOI321xp33_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_337),
.A3(n_249),
.B1(n_311),
.B2(n_224),
.C(n_256),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_256),
.Y(n_347)
);


endmodule