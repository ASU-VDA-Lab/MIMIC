module fake_jpeg_15762_n_79 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_79);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx2_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_24),
.B(n_27),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_13),
.B(n_1),
.Y(n_27)
);

INVxp33_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_18),
.A2(n_16),
.B1(n_15),
.B2(n_19),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_16),
.B1(n_15),
.B2(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_22),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_3),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_39),
.B1(n_40),
.B2(n_30),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_19),
.B1(n_3),
.B2(n_17),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_44),
.B1(n_34),
.B2(n_45),
.Y(n_53)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_17),
.B1(n_22),
.B2(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_25),
.A2(n_22),
.B1(n_14),
.B2(n_9),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_42),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_14),
.C(n_8),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_49),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_7),
.C(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_53),
.B1(n_39),
.B2(n_44),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_58),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_35),
.B(n_41),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_53),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_41),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_64),
.C(n_65),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_65),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_55),
.Y(n_70)
);

MAJx2_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_48),
.C(n_49),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_37),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_58),
.C(n_50),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_38),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_73)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_59),
.C(n_66),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_75),
.C(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_77),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_75),
.Y(n_79)
);


endmodule