module real_jpeg_29199_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_292;
wire n_215;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_293;
wire n_200;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_167;
wire n_216;
wire n_213;
wire n_128;
wire n_179;
wire n_202;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_127;
wire n_53;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_0),
.A2(n_74),
.B1(n_75),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_0),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_125),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_125),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_0),
.A2(n_45),
.B1(n_48),
.B2(n_125),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_1),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_1),
.B(n_70),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_1),
.B(n_27),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g216 ( 
.A1(n_1),
.A2(n_27),
.B(n_212),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_170),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_1),
.A2(n_45),
.B(n_49),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_1),
.B(n_119),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_1),
.A2(n_87),
.B1(n_115),
.B2(n_260),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_2),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_3),
.A2(n_38),
.B1(n_45),
.B2(n_48),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_7),
.A2(n_74),
.B1(n_75),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_7),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_172),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_172),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_7),
.A2(n_45),
.B1(n_48),
.B2(n_172),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_8),
.A2(n_74),
.B1(n_75),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_8),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_151),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_151),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_8),
.A2(n_45),
.B1(n_48),
.B2(n_151),
.Y(n_252)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_10),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_10),
.A2(n_42),
.B1(n_74),
.B2(n_75),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_42),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_11),
.A2(n_55),
.B1(n_74),
.B2(n_75),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_11),
.A2(n_45),
.B1(n_48),
.B2(n_55),
.Y(n_112)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_13),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_13),
.Y(n_211)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_14),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_15),
.A2(n_36),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_15),
.A2(n_36),
.B1(n_45),
.B2(n_48),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_100),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_19),
.B(n_100),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_84),
.B2(n_85),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_56),
.B2(n_57),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_23),
.A2(n_24),
.B(n_39),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_25),
.B(n_67),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_25),
.A2(n_31),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_25),
.A2(n_31),
.B1(n_166),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_25),
.A2(n_31),
.B1(n_195),
.B2(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_27),
.A2(n_28),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_27),
.B(n_71),
.Y(n_184)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_28),
.A2(n_79),
.B1(n_169),
.B2(n_184),
.Y(n_183)
);

AOI32xp33_ASAP7_75t_L g208 ( 
.A1(n_28),
.A2(n_32),
.A3(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_31),
.B(n_147),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_33),
.B1(n_47),
.B2(n_49),
.Y(n_53)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g213 ( 
.A(n_33),
.B(n_210),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_33),
.A2(n_47),
.B(n_170),
.C(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_35),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_50),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_40),
.A2(n_52),
.B(n_220),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_43),
.B(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_52),
.B(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_44),
.A2(n_52),
.B1(n_95),
.B2(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_44),
.A2(n_50),
.B(n_117),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_44),
.A2(n_52),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_44),
.A2(n_52),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_44),
.A2(n_52),
.B1(n_219),
.B2(n_237),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_44),
.B(n_170),
.Y(n_258)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_48),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_52),
.A2(n_61),
.B(n_96),
.Y(n_163)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_68),
.B1(n_82),
.B2(n_83),
.Y(n_57)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_64),
.A2(n_66),
.B(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_64),
.A2(n_180),
.B(n_181),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B(n_77),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_81),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_69),
.A2(n_123),
.B1(n_124),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_69),
.A2(n_123),
.B1(n_150),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_71),
.B(n_75),
.C(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_70),
.B(n_98),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_70),
.A2(n_78),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_75),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g169 ( 
.A(n_75),
.B(n_170),
.CON(n_169),
.SN(n_169)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_93),
.B(n_97),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_97),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_86),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_86),
.A2(n_94),
.B1(n_104),
.B2(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_90),
.B(n_91),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_87),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_87),
.A2(n_115),
.B1(n_141),
.B2(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_87),
.A2(n_113),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_87),
.A2(n_199),
.B1(n_252),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_88),
.A2(n_92),
.B(n_143),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_88),
.A2(n_114),
.B1(n_251),
.B2(n_253),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_112),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_94),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_97),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.C(n_106),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_101),
.B(n_105),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_106),
.A2(n_107),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_118),
.C(n_121),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_116),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_109),
.B(n_116),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_110),
.A2(n_186),
.B(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_121),
.B1(n_122),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B(n_126),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_155),
.B(n_303),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_152),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_131),
.B(n_152),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.C(n_138),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_132),
.A2(n_133),
.B1(n_136),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_136),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_138),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.C(n_148),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_139),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_144),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_145),
.A2(n_148),
.B1(n_149),
.B2(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_145),
.Y(n_293)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_297),
.B(n_302),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_200),
.B(n_283),
.C(n_296),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_187),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_158),
.B(n_187),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_173),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_160),
.B(n_161),
.C(n_173),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_168),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_168),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_170),
.B(n_199),
.Y(n_264)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_182),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_175),
.B(n_179),
.C(n_182),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.C(n_193),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_188),
.A2(n_189),
.B1(n_278),
.B2(n_280),
.Y(n_277)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_193),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.C(n_198),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_198),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_282),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_275),
.B(n_281),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_230),
.B(n_274),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_221),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_204),
.B(n_221),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_214),
.C(n_217),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_205),
.A2(n_206),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_208),
.Y(n_228)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_228),
.C(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_268),
.B(n_273),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_248),
.B(n_267),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_233),
.B(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_234),
.A2(n_235),
.B1(n_238),
.B2(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_246),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_247),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_256),
.B(n_266),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_254),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_261),
.B(n_265),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_259),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_276),
.B(n_277),
.Y(n_281)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_285),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_294),
.B2(n_295),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_291),
.C(n_295),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);


endmodule