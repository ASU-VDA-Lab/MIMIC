module fake_jpeg_26395_n_247 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_39),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_34),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_30),
.B1(n_23),
.B2(n_26),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_60),
.B1(n_63),
.B2(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_43),
.Y(n_70)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_56),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_64),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_28),
.C(n_33),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_28),
.C(n_33),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_25),
.B1(n_30),
.B2(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_17),
.B1(n_29),
.B2(n_22),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_41),
.B1(n_22),
.B2(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_34),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_69),
.B(n_76),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_75),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_43),
.B1(n_32),
.B2(n_28),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_58),
.B1(n_33),
.B2(n_32),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_82),
.Y(n_120)
);

AND2x4_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_43),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_96),
.B(n_58),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_81),
.B(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_17),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_84),
.B(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_17),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_35),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_77),
.Y(n_116)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_29),
.B1(n_31),
.B2(n_18),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_29),
.B1(n_51),
.B2(n_57),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_94),
.C(n_68),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_32),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_35),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_33),
.Y(n_101)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_100),
.Y(n_124)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_101),
.B(n_103),
.Y(n_144)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_31),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_18),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_104),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_1),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_SL g139 ( 
.A(n_105),
.B(n_106),
.C(n_96),
.Y(n_139)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_16),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_108),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_112),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_93),
.B(n_95),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_46),
.C(n_58),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_79),
.B1(n_88),
.B2(n_87),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_94),
.Y(n_137)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_71),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_81),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_139),
.B1(n_102),
.B2(n_114),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_79),
.B(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_137),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_79),
.B1(n_89),
.B2(n_72),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_142),
.B1(n_132),
.B2(n_126),
.Y(n_171)
);

AND2x6_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_76),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_136),
.B(n_138),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_85),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_73),
.B(n_72),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_142),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_118),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_84),
.B(n_86),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_117),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_32),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_146),
.B(n_113),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_112),
.A2(n_95),
.B1(n_93),
.B2(n_3),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_121),
.B1(n_107),
.B2(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_150),
.Y(n_191)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_144),
.B(n_109),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_153),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_120),
.C(n_119),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_135),
.C(n_131),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_121),
.A3(n_120),
.B1(n_109),
.B2(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_157),
.A2(n_134),
.B1(n_127),
.B2(n_137),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_158),
.B(n_133),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_171),
.B1(n_127),
.B2(n_137),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_160),
.B(n_162),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_161),
.B(n_164),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_114),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_102),
.A3(n_100),
.B1(n_98),
.B2(n_4),
.Y(n_163)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_16),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_166),
.Y(n_179)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_129),
.B(n_1),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_172),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_167),
.A2(n_147),
.B1(n_139),
.B2(n_140),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_174),
.A2(n_185),
.B1(n_168),
.B2(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_183),
.Y(n_201)
);

NOR2xp67_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_125),
.Y(n_181)
);

OAI322xp33_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_169),
.A3(n_150),
.B1(n_15),
.B2(n_14),
.C1(n_7),
.C2(n_8),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_188),
.C(n_156),
.Y(n_195)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_187),
.B(n_190),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_131),
.C(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_15),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_155),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_194),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_197),
.C(n_186),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_172),
.C(n_155),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_176),
.B1(n_180),
.B2(n_187),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_166),
.B(n_165),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_199),
.A2(n_179),
.B(n_184),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_169),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_203),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_6),
.C(n_7),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_2),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_205),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_2),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_175),
.B1(n_183),
.B2(n_189),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_215),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_213),
.Y(n_221)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_191),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_219),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_217),
.B(n_218),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_175),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_182),
.A3(n_190),
.B1(n_173),
.B2(n_9),
.C1(n_10),
.C2(n_6),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_220),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_213),
.A2(n_198),
.B1(n_194),
.B2(n_193),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_223),
.B1(n_221),
.B2(n_224),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_199),
.B1(n_207),
.B2(n_197),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_196),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_214),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_216),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_232),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_208),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_230),
.B(n_231),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_227),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_235),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_210),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_225),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_208),
.B(n_8),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_230),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_243),
.B(n_12),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_7),
.C(n_9),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_241),
.A2(n_237),
.B(n_11),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_245),
.B1(n_12),
.B2(n_242),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g247 ( 
.A(n_246),
.Y(n_247)
);


endmodule