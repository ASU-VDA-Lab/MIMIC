module fake_jpeg_3886_n_259 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_259);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_259;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_8),
.B(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_20),
.B1(n_23),
.B2(n_25),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_20),
.B1(n_33),
.B2(n_34),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_20),
.B(n_19),
.C(n_17),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_19),
.B(n_15),
.C(n_25),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_49),
.Y(n_68)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_55),
.Y(n_64)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_61),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_14),
.B1(n_24),
.B2(n_17),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_30),
.B1(n_15),
.B2(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_25),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_15),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_62),
.B(n_15),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_75),
.B(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_15),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_78),
.B(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_32),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_39),
.B(n_14),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_36),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_57),
.B1(n_59),
.B2(n_49),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_86),
.B1(n_73),
.B2(n_65),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_71),
.B(n_69),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_85),
.B(n_92),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_87),
.B(n_75),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_57),
.B(n_62),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_51),
.B1(n_47),
.B2(n_62),
.Y(n_86)
);

XOR2x2_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_62),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_53),
.C(n_39),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_89),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_36),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_93),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_14),
.Y(n_96)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_64),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_103),
.B(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_91),
.B1(n_88),
.B2(n_95),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_113),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_110),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_72),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_72),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_64),
.B1(n_80),
.B2(n_78),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_117),
.B1(n_84),
.B2(n_85),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_78),
.B1(n_75),
.B2(n_60),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_83),
.B(n_92),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_136),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_109),
.A2(n_87),
.B1(n_83),
.B2(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_124),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_114),
.B1(n_115),
.B2(n_95),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_125),
.B(n_113),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_116),
.A2(n_90),
.B1(n_88),
.B2(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

AOI22x1_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_92),
.B1(n_84),
.B2(n_85),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_111),
.B1(n_106),
.B2(n_100),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_118),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_133),
.C(n_122),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_89),
.C(n_90),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_106),
.B1(n_105),
.B2(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_76),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_135),
.B(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_89),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_96),
.B1(n_58),
.B2(n_60),
.Y(n_137)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_153),
.C(n_154),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_126),
.B1(n_134),
.B2(n_52),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_112),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_158),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_152),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_112),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_151),
.A2(n_125),
.B(n_130),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_79),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_37),
.C(n_32),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_37),
.C(n_27),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_76),
.B(n_12),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_137),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_37),
.C(n_28),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_121),
.C(n_128),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_37),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_131),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_159),
.A2(n_131),
.B(n_126),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_18),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_145),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_153),
.C(n_26),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_58),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_18),
.B(n_13),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_46),
.B(n_41),
.C(n_21),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_37),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_173),
.C(n_31),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_179),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_52),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_50),
.B1(n_48),
.B2(n_24),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_28),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_178),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_158),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_50),
.B1(n_22),
.B2(n_21),
.Y(n_179)
);

NAND2x1_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_151),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_183),
.B(n_188),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_163),
.A2(n_139),
.B1(n_157),
.B2(n_152),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_186),
.Y(n_201)
);

FAx1_ASAP7_75t_SL g186 ( 
.A(n_170),
.B(n_141),
.CI(n_154),
.CON(n_186),
.SN(n_186)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_167),
.C(n_161),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_0),
.B(n_1),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_195),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_18),
.Y(n_192)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_0),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_197),
.C(n_188),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_1),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_164),
.B(n_13),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_202),
.C(n_207),
.Y(n_216)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_161),
.C(n_167),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_178),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_208),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_205),
.A2(n_13),
.B(n_21),
.Y(n_227)
);

AO221x1_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_46),
.B1(n_41),
.B2(n_177),
.C(n_13),
.Y(n_206)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_46),
.C(n_41),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_183),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_181),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_21),
.B1(n_22),
.B2(n_13),
.Y(n_211)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_198),
.B1(n_190),
.B2(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

AO21x1_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_201),
.B(n_209),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_215),
.A2(n_220),
.B(n_222),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_203),
.B(n_191),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_12),
.C(n_26),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_197),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_226),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_194),
.B(n_186),
.Y(n_222)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_1),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_219),
.B(n_186),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_216),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_230),
.B(n_233),
.Y(n_245)
);

NOR2xp67_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_31),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_235),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_18),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_234),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_18),
.Y(n_235)
);

INVx11_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_216),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_18),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_239),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_240),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_244),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_218),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_247),
.B(n_2),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_237),
.B1(n_233),
.B2(n_231),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_227),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_245),
.A2(n_2),
.B(n_5),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_252),
.C(n_253),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_246),
.A2(n_11),
.B(n_6),
.Y(n_253)
);

AOI321xp33_ASAP7_75t_L g255 ( 
.A1(n_249),
.A2(n_247),
.A3(n_248),
.B1(n_242),
.B2(n_8),
.C(n_5),
.Y(n_255)
);

OAI321xp33_ASAP7_75t_L g257 ( 
.A1(n_255),
.A2(n_256),
.A3(n_7),
.B1(n_9),
.B2(n_10),
.C(n_254),
.Y(n_257)
);

NOR2x1_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_5),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_257),
.A2(n_9),
.B(n_10),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_258),
.Y(n_259)
);


endmodule