module fake_netlist_1_11508_n_687 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_687);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_687;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_490;
wire n_247;
wire n_613;
wire n_393;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_582;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_2), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_14), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_54), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_21), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_22), .Y(n_84) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_63), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_5), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_3), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_78), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_66), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_30), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_70), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_64), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_77), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_57), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_28), .Y(n_95) );
BUFx6f_ASAP7_75t_L g96 ( .A(n_20), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_32), .Y(n_97) );
BUFx2_ASAP7_75t_L g98 ( .A(n_76), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_29), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_73), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_45), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_8), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_38), .Y(n_103) );
CKINVDCx14_ASAP7_75t_R g104 ( .A(n_25), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_5), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_47), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_61), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_41), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_50), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_1), .Y(n_110) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_26), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_17), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_72), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_67), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_18), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_9), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_74), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_44), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_48), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_68), .Y(n_121) );
BUFx5_ASAP7_75t_L g122 ( .A(n_53), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_14), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_71), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_123), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_92), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_124), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_92), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_123), .B(n_0), .Y(n_129) );
INVx2_ASAP7_75t_SL g130 ( .A(n_98), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_93), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_93), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_98), .B(n_4), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_96), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_124), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_120), .B(n_4), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_124), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_117), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_96), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_122), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_117), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g142 ( .A1(n_80), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_122), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_120), .B(n_6), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_96), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_122), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_96), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_80), .B(n_7), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_102), .B(n_9), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_83), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_102), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_96), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_122), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_99), .Y(n_155) );
BUFx8_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_108), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_108), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_91), .B(n_10), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_122), .B(n_10), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_110), .B(n_11), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_108), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_91), .B(n_11), .Y(n_163) );
INVx1_ASAP7_75t_SL g164 ( .A(n_144), .Y(n_164) );
OR2x2_ASAP7_75t_L g165 ( .A(n_130), .B(n_86), .Y(n_165) );
AND2x6_ASAP7_75t_L g166 ( .A(n_133), .B(n_107), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_130), .B(n_106), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_148), .Y(n_168) );
OR2x2_ASAP7_75t_L g169 ( .A(n_129), .B(n_86), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_156), .B(n_85), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_150), .B(n_82), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_133), .B(n_107), .Y(n_173) );
INVx5_ASAP7_75t_L g174 ( .A(n_159), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_129), .B(n_111), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_150), .B(n_109), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_154), .B(n_112), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_127), .B(n_126), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_154), .B(n_103), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_155), .B(n_113), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_148), .Y(n_183) );
OR2x6_ASAP7_75t_L g184 ( .A(n_133), .B(n_81), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_138), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_127), .B(n_89), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
INVx1_ASAP7_75t_SL g192 ( .A(n_133), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_127), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_149), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_159), .A2(n_87), .B1(n_116), .B2(n_105), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_159), .A2(n_94), .B1(n_121), .B2(n_90), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_151), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_126), .B(n_128), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_128), .B(n_89), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_138), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_155), .B(n_100), .Y(n_202) );
INVxp67_ASAP7_75t_L g203 ( .A(n_136), .Y(n_203) );
OR2x2_ASAP7_75t_L g204 ( .A(n_161), .B(n_84), .Y(n_204) );
NAND3xp33_ASAP7_75t_L g205 ( .A(n_156), .B(n_84), .C(n_121), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_131), .B(n_101), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_156), .Y(n_207) );
BUFx10_ASAP7_75t_L g208 ( .A(n_163), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_151), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_131), .B(n_119), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_177), .B(n_132), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_187), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_164), .B(n_132), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_188), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_180), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_168), .A2(n_163), .B(n_140), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_164), .B(n_156), .Y(n_217) );
NOR2xp33_ASAP7_75t_SL g218 ( .A(n_207), .B(n_88), .Y(n_218) );
NAND2x1p5_ASAP7_75t_L g219 ( .A(n_170), .B(n_163), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_176), .B(n_151), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_184), .B(n_163), .Y(n_221) );
AND2x6_ASAP7_75t_SL g222 ( .A(n_167), .B(n_125), .Y(n_222) );
INVx8_ASAP7_75t_L g223 ( .A(n_184), .Y(n_223) );
BUFx5_ASAP7_75t_L g224 ( .A(n_166), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_201), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_180), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_192), .B(n_143), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_203), .B(n_141), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_204), .B(n_141), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_199), .Y(n_230) );
NAND2xp33_ASAP7_75t_SL g231 ( .A(n_196), .B(n_88), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_171), .B(n_90), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_172), .A2(n_137), .B1(n_135), .B2(n_146), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_199), .B(n_97), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_184), .A2(n_125), .B1(n_142), .B2(n_160), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_192), .B(n_97), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_190), .B(n_118), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_190), .Y(n_238) );
OAI22xp5_ASAP7_75t_SL g239 ( .A1(n_197), .A2(n_115), .B1(n_118), .B2(n_104), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_169), .A2(n_137), .B(n_135), .C(n_140), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_198), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_193), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_165), .B(n_115), .Y(n_243) );
INVx1_ASAP7_75t_SL g244 ( .A(n_189), .Y(n_244) );
BUFx2_ASAP7_75t_L g245 ( .A(n_166), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_209), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_166), .B(n_153), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_166), .B(n_153), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_166), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_173), .B(n_143), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_183), .A2(n_146), .B(n_101), .Y(n_251) );
AND2x4_ASAP7_75t_SL g252 ( .A(n_208), .B(n_114), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_185), .A2(n_114), .B1(n_122), .B2(n_108), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_208), .B(n_122), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_173), .B(n_108), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_191), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_191), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_173), .B(n_162), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_174), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_173), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_186), .A2(n_162), .B1(n_158), .B2(n_157), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_173), .B(n_162), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_194), .B(n_162), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_195), .B(n_162), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_174), .B(n_158), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_189), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g267 ( .A1(n_200), .A2(n_12), .B(n_13), .C(n_15), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_243), .B(n_205), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_216), .A2(n_174), .B(n_206), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_256), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_223), .Y(n_271) );
BUFx6f_ASAP7_75t_SL g272 ( .A(n_221), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_243), .B(n_232), .Y(n_273) );
NAND2x1p5_ASAP7_75t_L g274 ( .A(n_221), .B(n_174), .Y(n_274) );
AOI21x1_ASAP7_75t_SL g275 ( .A1(n_255), .A2(n_206), .B(n_200), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_211), .B(n_202), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_256), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_227), .A2(n_210), .B(n_182), .Y(n_278) );
INVx4_ASAP7_75t_L g279 ( .A(n_223), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_230), .A2(n_181), .B(n_179), .C(n_178), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_215), .A2(n_147), .B1(n_158), .B2(n_157), .Y(n_281) );
NOR3xp33_ASAP7_75t_SL g282 ( .A(n_239), .B(n_231), .C(n_228), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_223), .A2(n_147), .B1(n_158), .B2(n_157), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_244), .Y(n_284) );
AOI21x1_ASAP7_75t_L g285 ( .A1(n_258), .A2(n_175), .B(n_158), .Y(n_285) );
O2A1O1Ixp5_ASAP7_75t_L g286 ( .A1(n_254), .A2(n_175), .B(n_49), .C(n_51), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_222), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_238), .Y(n_288) );
AOI21x1_ASAP7_75t_L g289 ( .A1(n_262), .A2(n_175), .B(n_157), .Y(n_289) );
BUFx12f_ASAP7_75t_L g290 ( .A(n_219), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g291 ( .A1(n_213), .A2(n_12), .B(n_13), .C(n_15), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_249), .Y(n_292) );
OAI22x1_ASAP7_75t_L g293 ( .A1(n_235), .A2(n_16), .B1(n_19), .B2(n_23), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_257), .Y(n_294) );
OR2x6_ASAP7_75t_L g295 ( .A(n_249), .B(n_157), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_238), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_266), .B(n_152), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_228), .B(n_24), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_241), .Y(n_299) );
NAND2xp33_ASAP7_75t_SL g300 ( .A(n_245), .B(n_152), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_226), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_242), .Y(n_302) );
OR2x6_ASAP7_75t_SL g303 ( .A(n_217), .B(n_27), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_229), .B(n_152), .Y(n_304) );
AND2x6_ASAP7_75t_L g305 ( .A(n_260), .B(n_152), .Y(n_305) );
OR2x6_ASAP7_75t_L g306 ( .A(n_260), .B(n_152), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_252), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_229), .B(n_147), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_241), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_234), .A2(n_147), .B1(n_145), .B2(n_139), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_233), .A2(n_147), .B1(n_145), .B2(n_139), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_220), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_246), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_252), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_246), .B(n_145), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_242), .B(n_31), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_224), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_227), .A2(n_145), .B(n_139), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_299), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_275), .A2(n_251), .B(n_264), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_301), .Y(n_321) );
OA21x2_ASAP7_75t_L g322 ( .A1(n_318), .A2(n_253), .B(n_265), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_297), .A2(n_254), .B(n_248), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_284), .B(n_236), .Y(n_324) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_279), .B(n_259), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_309), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_297), .A2(n_247), .B(n_250), .Y(n_327) );
OAI22xp33_ASAP7_75t_L g328 ( .A1(n_303), .A2(n_219), .B1(n_218), .B2(n_237), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_280), .A2(n_240), .B(n_267), .C(n_253), .Y(n_329) );
O2A1O1Ixp5_ASAP7_75t_L g330 ( .A1(n_311), .A2(n_263), .B(n_259), .C(n_212), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_312), .B(n_233), .Y(n_331) );
BUFx12f_ASAP7_75t_L g332 ( .A(n_279), .Y(n_332) );
AO31x2_ASAP7_75t_L g333 ( .A1(n_293), .A2(n_263), .A3(n_214), .B(n_225), .Y(n_333) );
NAND3x1_ASAP7_75t_L g334 ( .A(n_268), .B(n_224), .C(n_34), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_273), .B(n_224), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_276), .B(n_224), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_SL g337 ( .A1(n_304), .A2(n_225), .B(n_214), .C(n_212), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_272), .B(n_224), .Y(n_338) );
A2O1A1Ixp33_ASAP7_75t_L g339 ( .A1(n_278), .A2(n_261), .B(n_224), .C(n_145), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_290), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g341 ( .A1(n_269), .A2(n_261), .B(n_139), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_SL g342 ( .A1(n_304), .A2(n_33), .B(n_35), .C(n_36), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_318), .A2(n_139), .B(n_134), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_287), .A2(n_134), .B1(n_39), .B2(n_40), .C(n_42), .Y(n_344) );
INVxp67_ASAP7_75t_SL g345 ( .A(n_313), .Y(n_345) );
AOI21x1_ASAP7_75t_L g346 ( .A1(n_285), .A2(n_134), .B(n_43), .Y(n_346) );
OAI221xp5_ASAP7_75t_L g347 ( .A1(n_282), .A2(n_134), .B1(n_46), .B2(n_52), .C(n_55), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_298), .A2(n_37), .B(n_56), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_314), .B(n_58), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_315), .A2(n_59), .B(n_60), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_308), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_271), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_294), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_326), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_337), .A2(n_315), .B(n_311), .Y(n_356) );
OAI21xp5_ASAP7_75t_L g357 ( .A1(n_329), .A2(n_291), .B(n_316), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_345), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_353), .Y(n_359) );
OAI221xp5_ASAP7_75t_L g360 ( .A1(n_324), .A2(n_314), .B1(n_307), .B2(n_310), .C(n_274), .Y(n_360) );
INVx4_ASAP7_75t_L g361 ( .A(n_332), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_321), .B(n_307), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_340), .Y(n_363) );
A2O1A1Ixp33_ASAP7_75t_L g364 ( .A1(n_336), .A2(n_316), .B(n_286), .C(n_270), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_320), .Y(n_365) );
OA21x2_ASAP7_75t_L g366 ( .A1(n_330), .A2(n_289), .B(n_281), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_346), .A2(n_281), .B(n_283), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_337), .A2(n_345), .B(n_336), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_328), .B(n_272), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_328), .B(n_302), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_331), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_351), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_335), .A2(n_288), .B1(n_296), .B2(n_277), .Y(n_373) );
AO21x2_ASAP7_75t_L g374 ( .A1(n_339), .A2(n_317), .B(n_300), .Y(n_374) );
OR2x6_ASAP7_75t_L g375 ( .A(n_325), .B(n_306), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_325), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_352), .B(n_296), .Y(n_377) );
AOI21x1_ASAP7_75t_L g378 ( .A1(n_343), .A2(n_306), .B(n_295), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_322), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_323), .A2(n_317), .B(n_306), .Y(n_380) );
OA21x2_ASAP7_75t_L g381 ( .A1(n_330), .A2(n_305), .B(n_295), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_334), .A2(n_274), .B(n_305), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_379), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_358), .B(n_333), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_363), .B(n_338), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_381), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_379), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_363), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_381), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_354), .B(n_333), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_354), .B(n_333), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_365), .Y(n_392) );
AOI21x1_ASAP7_75t_L g393 ( .A1(n_368), .A2(n_348), .B(n_350), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_358), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_369), .B(n_338), .Y(n_395) );
OR2x6_ASAP7_75t_L g396 ( .A(n_375), .B(n_295), .Y(n_396) );
INVx5_ASAP7_75t_SL g397 ( .A(n_375), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_359), .B(n_335), .Y(n_398) );
AO21x2_ASAP7_75t_L g399 ( .A1(n_356), .A2(n_347), .B(n_341), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_365), .Y(n_400) );
AOI21x1_ASAP7_75t_L g401 ( .A1(n_381), .A2(n_349), .B(n_322), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_375), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_355), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_371), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_355), .Y(n_405) );
AO21x2_ASAP7_75t_L g406 ( .A1(n_357), .A2(n_342), .B(n_327), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_372), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_366), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_366), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_370), .A2(n_344), .B1(n_322), .B2(n_292), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_372), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_376), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_376), .B(n_333), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_370), .B(n_292), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_404), .B(n_377), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_385), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_404), .B(n_362), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_383), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_386), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_397), .A2(n_360), .B1(n_375), .B2(n_373), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_383), .B(n_374), .Y(n_421) );
INVx5_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
NOR2xp33_ASAP7_75t_R g423 ( .A(n_388), .B(n_361), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_383), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_387), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_387), .Y(n_427) );
INVx4_ASAP7_75t_L g428 ( .A(n_396), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_394), .B(n_374), .Y(n_429) );
INVx5_ASAP7_75t_L g430 ( .A(n_396), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_394), .B(n_374), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_403), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_405), .B(n_366), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_405), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_407), .B(n_361), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_403), .B(n_361), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_402), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_403), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_384), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_392), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_384), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_384), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_384), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_407), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_413), .B(n_382), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_392), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_390), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_411), .B(n_382), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_392), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_411), .B(n_364), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_390), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_391), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_386), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_391), .Y(n_454) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_386), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_400), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_413), .B(n_367), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_400), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_427), .Y(n_459) );
AO31x2_ASAP7_75t_L g460 ( .A1(n_427), .A2(n_408), .A3(n_409), .B(n_400), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_447), .B(n_408), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_439), .B(n_409), .Y(n_462) );
BUFx2_ASAP7_75t_L g463 ( .A(n_428), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_436), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_434), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_458), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_434), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_458), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_447), .B(n_409), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_418), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_451), .B(n_408), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_418), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_458), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_451), .B(n_414), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_424), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_452), .B(n_414), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_452), .B(n_389), .Y(n_477) );
INVx4_ASAP7_75t_L g478 ( .A(n_422), .Y(n_478) );
NOR2xp67_ASAP7_75t_L g479 ( .A(n_422), .B(n_389), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_454), .B(n_389), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_424), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_439), .B(n_389), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_454), .B(n_389), .Y(n_483) );
INVx1_ASAP7_75t_SL g484 ( .A(n_423), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_441), .B(n_389), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_419), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_415), .B(n_412), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_441), .B(n_386), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_425), .B(n_412), .Y(n_489) );
INVxp67_ASAP7_75t_L g490 ( .A(n_436), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_425), .B(n_397), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_444), .B(n_398), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_426), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_442), .B(n_386), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_417), .B(n_395), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_426), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_416), .A2(n_402), .B1(n_397), .B2(n_396), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_442), .B(n_386), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_432), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_428), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_432), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_443), .B(n_397), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_443), .B(n_401), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_438), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_457), .B(n_401), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_435), .B(n_402), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_448), .Y(n_507) );
BUFx3_ASAP7_75t_L g508 ( .A(n_437), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_440), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_437), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_438), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_422), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_457), .B(n_431), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_429), .B(n_397), .Y(n_514) );
NAND2x1p5_ASAP7_75t_L g515 ( .A(n_422), .B(n_396), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_429), .B(n_431), .Y(n_516) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_484), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_464), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_495), .A2(n_428), .B1(n_420), .B2(n_430), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_516), .B(n_433), .Y(n_520) );
OAI211xp5_ASAP7_75t_L g521 ( .A1(n_497), .A2(n_428), .B(n_422), .C(n_430), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_513), .B(n_456), .Y(n_522) );
OAI211xp5_ASAP7_75t_L g523 ( .A1(n_463), .A2(n_422), .B(n_430), .C(n_448), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_465), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_516), .B(n_433), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_465), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_513), .B(n_445), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_467), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_467), .B(n_421), .Y(n_529) );
NAND2x1_ASAP7_75t_L g530 ( .A(n_478), .B(n_445), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_474), .B(n_445), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_490), .B(n_456), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_470), .B(n_421), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_474), .B(n_476), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_470), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_472), .Y(n_536) );
INVxp67_ASAP7_75t_SL g537 ( .A(n_466), .Y(n_537) );
BUFx3_ASAP7_75t_L g538 ( .A(n_508), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_463), .B(n_445), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_472), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_476), .B(n_446), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_475), .B(n_450), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_481), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_508), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_503), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_507), .B(n_430), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_478), .B(n_430), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_475), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_496), .B(n_450), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_505), .B(n_430), .Y(n_550) );
INVx3_ASAP7_75t_SL g551 ( .A(n_478), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_496), .B(n_440), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_505), .B(n_419), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_500), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_461), .B(n_449), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_492), .B(n_449), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_489), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_510), .B(n_453), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_489), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_514), .B(n_453), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_481), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_493), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_514), .B(n_471), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_469), .B(n_446), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_461), .B(n_453), .Y(n_565) );
NAND2xp33_ASAP7_75t_L g566 ( .A(n_515), .B(n_410), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_477), .B(n_453), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_471), .B(n_419), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_500), .B(n_419), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_477), .B(n_455), .Y(n_570) );
NOR2x1_ASAP7_75t_L g571 ( .A(n_479), .B(n_406), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_493), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_466), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_503), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_517), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_551), .B(n_479), .Y(n_576) );
NAND2x1_ASAP7_75t_L g577 ( .A(n_547), .B(n_512), .Y(n_577) );
AOI21xp33_ASAP7_75t_L g578 ( .A1(n_566), .A2(n_487), .B(n_512), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_557), .B(n_483), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_556), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_527), .B(n_483), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_534), .B(n_480), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_573), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_524), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_526), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_559), .B(n_480), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_518), .B(n_506), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_528), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_535), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_536), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_540), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_545), .B(n_469), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_519), .A2(n_515), .B1(n_502), .B2(n_491), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_545), .B(n_486), .Y(n_594) );
NAND2x1p5_ASAP7_75t_L g595 ( .A(n_547), .B(n_491), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_520), .B(n_511), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_574), .B(n_494), .Y(n_597) );
AOI32xp33_ASAP7_75t_L g598 ( .A1(n_554), .A2(n_494), .A3(n_485), .B1(n_498), .B2(n_486), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_574), .B(n_486), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_563), .B(n_498), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_548), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_531), .B(n_485), .Y(n_602) );
AOI31xp33_ASAP7_75t_L g603 ( .A1(n_521), .A2(n_515), .A3(n_502), .B(n_504), .Y(n_603) );
INVxp67_ASAP7_75t_L g604 ( .A(n_573), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_538), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_542), .B(n_462), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_551), .Y(n_607) );
A2O1A1Ixp33_ASAP7_75t_L g608 ( .A1(n_523), .A2(n_511), .B(n_499), .C(n_504), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_530), .A2(n_501), .B1(n_499), .B2(n_459), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_520), .B(n_488), .Y(n_610) );
INVxp33_ASAP7_75t_L g611 ( .A(n_569), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_525), .B(n_488), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_550), .A2(n_488), .B1(n_482), .B2(n_462), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_525), .B(n_482), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_553), .B(n_482), .Y(n_615) );
INVx2_ASAP7_75t_SL g616 ( .A(n_544), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_560), .B(n_462), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_522), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_580), .B(n_549), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_587), .A2(n_539), .B1(n_567), .B2(n_546), .Y(n_620) );
OAI211xp5_ASAP7_75t_L g621 ( .A1(n_607), .A2(n_521), .B(n_523), .C(n_542), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_596), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_615), .B(n_539), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_603), .A2(n_541), .B1(n_537), .B2(n_532), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_592), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_578), .A2(n_549), .B1(n_529), .B2(n_533), .C(n_555), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_610), .B(n_568), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_579), .B(n_586), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_597), .B(n_555), .Y(n_629) );
OAI211xp5_ASAP7_75t_SL g630 ( .A1(n_598), .A2(n_571), .B(n_529), .C(n_533), .Y(n_630) );
OAI221xp5_ASAP7_75t_L g631 ( .A1(n_593), .A2(n_558), .B1(n_564), .B2(n_552), .C(n_561), .Y(n_631) );
INVx2_ASAP7_75t_SL g632 ( .A(n_605), .Y(n_632) );
OAI21xp5_ASAP7_75t_SL g633 ( .A1(n_576), .A2(n_567), .B(n_565), .Y(n_633) );
INVx2_ASAP7_75t_SL g634 ( .A(n_575), .Y(n_634) );
AOI31xp33_ASAP7_75t_L g635 ( .A1(n_576), .A2(n_537), .A3(n_552), .B(n_572), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_616), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_587), .A2(n_562), .B1(n_543), .B2(n_570), .C(n_501), .Y(n_637) );
NAND4xp75_ASAP7_75t_L g638 ( .A(n_594), .B(n_459), .C(n_509), .D(n_473), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_577), .A2(n_570), .B1(n_509), .B2(n_473), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_611), .B(n_468), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_584), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_585), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_618), .B(n_468), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_594), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_614), .B(n_455), .Y(n_645) );
OAI22xp33_ASAP7_75t_L g646 ( .A1(n_635), .A2(n_595), .B1(n_613), .B2(n_609), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_630), .A2(n_612), .B1(n_599), .B2(n_604), .C(n_609), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_635), .A2(n_608), .B(n_604), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_643), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_629), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_644), .A2(n_599), .B1(n_612), .B2(n_593), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_624), .A2(n_608), .B(n_595), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_641), .Y(n_653) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_624), .A2(n_606), .B(n_590), .C(n_601), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_631), .A2(n_588), .B1(n_591), .B2(n_589), .C(n_582), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_633), .A2(n_583), .B(n_617), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_642), .Y(n_657) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_636), .A2(n_602), .B(n_581), .C(n_600), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_L g659 ( .A1(n_634), .A2(n_406), .B(n_399), .C(n_380), .Y(n_659) );
AOI21xp33_ASAP7_75t_SL g660 ( .A1(n_633), .A2(n_62), .B(n_65), .Y(n_660) );
OAI21xp33_ASAP7_75t_SL g661 ( .A1(n_632), .A2(n_367), .B(n_460), .Y(n_661) );
NAND4xp25_ASAP7_75t_SL g662 ( .A(n_652), .B(n_621), .C(n_620), .D(n_626), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_646), .A2(n_637), .B1(n_625), .B2(n_640), .C(n_619), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_649), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_651), .B(n_622), .Y(n_665) );
OAI211xp5_ASAP7_75t_L g666 ( .A1(n_652), .A2(n_639), .B(n_623), .C(n_628), .Y(n_666) );
NAND2xp33_ASAP7_75t_SL g667 ( .A(n_654), .B(n_627), .Y(n_667) );
NAND2xp33_ASAP7_75t_R g668 ( .A(n_660), .B(n_638), .Y(n_668) );
NAND5xp2_ASAP7_75t_L g669 ( .A(n_647), .B(n_393), .C(n_645), .D(n_378), .E(n_69), .Y(n_669) );
AOI211xp5_ASAP7_75t_L g670 ( .A1(n_648), .A2(n_455), .B(n_292), .C(n_393), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_662), .B(n_661), .C(n_655), .Y(n_671) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_663), .B(n_659), .C(n_657), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_667), .B(n_656), .Y(n_673) );
NAND5xp2_ASAP7_75t_L g674 ( .A(n_666), .B(n_658), .C(n_650), .D(n_653), .E(n_378), .Y(n_674) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_670), .B(n_455), .C(n_79), .Y(n_675) );
AND4x1_ASAP7_75t_L g676 ( .A(n_671), .B(n_665), .C(n_668), .D(n_669), .Y(n_676) );
NAND4xp25_ASAP7_75t_SL g677 ( .A(n_672), .B(n_664), .C(n_406), .D(n_399), .Y(n_677) );
NOR2x1p5_ASAP7_75t_L g678 ( .A(n_675), .B(n_455), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_678), .Y(n_679) );
OAI22xp5_ASAP7_75t_SL g680 ( .A1(n_676), .A2(n_674), .B1(n_673), .B2(n_455), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_679), .Y(n_681) );
INVx3_ASAP7_75t_SL g682 ( .A(n_680), .Y(n_682) );
NOR2x1_ASAP7_75t_L g683 ( .A(n_681), .B(n_677), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_683), .A2(n_682), .B(n_305), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_684), .B(n_75), .C(n_305), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_685), .A2(n_399), .B1(n_460), .B2(n_682), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_686), .A2(n_399), .B1(n_460), .B2(n_671), .Y(n_687) );
endmodule