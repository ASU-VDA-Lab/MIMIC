module fake_jpeg_7960_n_272 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_43),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_58),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_20),
.B1(n_29),
.B2(n_27),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_56),
.B1(n_61),
.B2(n_65),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_31),
.Y(n_74)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_20),
.B1(n_29),
.B2(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_20),
.B1(n_29),
.B2(n_18),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_23),
.B1(n_31),
.B2(n_19),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_28),
.B1(n_32),
.B2(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_63),
.Y(n_92)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_35),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_34),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_68),
.A2(n_78),
.B1(n_81),
.B2(n_90),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_30),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_70),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_60),
.B(n_48),
.C(n_62),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_0),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_73),
.B(n_74),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_75),
.B(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_96),
.B1(n_101),
.B2(n_34),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_0),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_23),
.B1(n_19),
.B2(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_30),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_80),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_59),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_45),
.A2(n_19),
.B1(n_22),
.B2(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_45),
.B(n_12),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_44),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_49),
.B(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_89),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_30),
.C(n_34),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_94),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_50),
.B(n_11),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_24),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_97),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_21),
.B1(n_10),
.B2(n_16),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_10),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_44),
.B(n_8),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_30),
.C(n_34),
.Y(n_101)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_104),
.Y(n_153)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_106),
.B(n_113),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_67),
.A2(n_34),
.B1(n_47),
.B2(n_8),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_108),
.A2(n_92),
.B1(n_101),
.B2(n_12),
.Y(n_151)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_109),
.Y(n_133)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_125),
.B1(n_91),
.B2(n_71),
.Y(n_137)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_82),
.B1(n_99),
.B2(n_100),
.Y(n_132)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_72),
.B(n_0),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_126),
.A2(n_72),
.B1(n_77),
.B2(n_94),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_141),
.B(n_144),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_69),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_135),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_110),
.B(n_74),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_118),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_134),
.B1(n_143),
.B2(n_148),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_121),
.B1(n_102),
.B2(n_106),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_97),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_72),
.B(n_77),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_145),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_71),
.B1(n_75),
.B2(n_86),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_77),
.B1(n_73),
.B2(n_70),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_155),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_95),
.C(n_89),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_107),
.C(n_117),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_91),
.B1(n_85),
.B2(n_84),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_79),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_1),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_70),
.B1(n_76),
.B2(n_87),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_157),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_92),
.B(n_2),
.C(n_3),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_116),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_122),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_108),
.A2(n_6),
.B1(n_15),
.B2(n_14),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_162),
.C(n_174),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_161),
.B(n_166),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_168),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_125),
.B1(n_104),
.B2(n_118),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_165),
.A2(n_181),
.B1(n_152),
.B2(n_139),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_107),
.B(n_103),
.C(n_15),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_1),
.B(n_2),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_172),
.A2(n_175),
.B(n_154),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_177),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_7),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_137),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_131),
.B(n_120),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_1),
.Y(n_179)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_129),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_180),
.B(n_135),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_112),
.B1(n_109),
.B2(n_105),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_6),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_150),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_192),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_175),
.A2(n_154),
.B1(n_148),
.B2(n_144),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_156),
.B1(n_135),
.B2(n_152),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_203),
.B1(n_205),
.B2(n_164),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_176),
.B1(n_169),
.B2(n_173),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_180),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_184),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_165),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_155),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_199),
.C(n_159),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_158),
.A2(n_139),
.B1(n_136),
.B2(n_133),
.Y(n_203)
);

NAND2xp33_ASAP7_75t_SL g204 ( 
.A(n_163),
.B(n_13),
.Y(n_204)
);

OAI321xp33_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_172),
.A3(n_166),
.B1(n_182),
.B2(n_176),
.C(n_181),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_183),
.A2(n_136),
.B1(n_133),
.B2(n_140),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_140),
.B(n_3),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_206),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_222),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_203),
.A2(n_160),
.B1(n_177),
.B2(n_158),
.Y(n_211)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_212),
.B(n_213),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_219),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_220),
.C(n_221),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_174),
.C(n_169),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_202),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_179),
.C(n_105),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_198),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_193),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_207),
.C(n_220),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_234),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_195),
.B1(n_189),
.B2(n_186),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_232),
.A2(n_236),
.B1(n_205),
.B2(n_196),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_206),
.B(n_190),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_217),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_238),
.B(n_227),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_237),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_188),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_224),
.B(n_211),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_247),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_218),
.B1(n_210),
.B2(n_196),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_242),
.A2(n_245),
.B(n_248),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_233),
.A2(n_194),
.B1(n_188),
.B2(n_192),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_249),
.A2(n_252),
.B(n_253),
.Y(n_259)
);

XNOR2x1_ASAP7_75t_SL g250 ( 
.A(n_244),
.B(n_228),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_229),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_194),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_254),
.B(n_256),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_243),
.Y(n_257)
);

NAND3xp33_ASAP7_75t_SL g265 ( 
.A(n_257),
.B(n_258),
.C(n_249),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_251),
.A2(n_236),
.B(n_248),
.Y(n_258)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_262),
.B(n_261),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_242),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_247),
.C(n_215),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_263),
.A2(n_264),
.B(n_265),
.C(n_266),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_238),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_226),
.C(n_249),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_267),
.A3(n_221),
.B1(n_7),
.B2(n_5),
.C1(n_13),
.C2(n_16),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_267),
.B(n_5),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_7),
.B1(n_13),
.B2(n_4),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_2),
.Y(n_272)
);


endmodule