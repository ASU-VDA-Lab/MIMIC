module fake_netlist_5_2416_n_91 (n_16, n_0, n_12, n_9, n_18, n_22, n_1, n_8, n_10, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_13, n_3, n_6, n_91);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_91;

wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_69;
wire n_58;
wire n_42;
wire n_45;
wire n_46;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_85;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_8),
.B(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_2),
.Y(n_34)
);

OAI22x1_ASAP7_75t_SL g35 ( 
.A1(n_12),
.A2(n_1),
.B1(n_3),
.B2(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

AOI221xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.C(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

O2A1O1Ixp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_22),
.B(n_31),
.C(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_25),
.Y(n_45)
);

NOR2xp67_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_26),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_36),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_45),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_36),
.B(n_30),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_32),
.B1(n_23),
.B2(n_37),
.Y(n_51)
);

AO31x2_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_35),
.A3(n_33),
.B(n_24),
.Y(n_52)
);

OAI21x1_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_24),
.B(n_33),
.Y(n_53)
);

OAI21x1_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_33),
.B(n_28),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_28),
.Y(n_55)
);

OA21x2_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_43),
.B(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

OAI21x1_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_47),
.B(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx2_ASAP7_75t_SL g68 ( 
.A(n_59),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_69),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_57),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_68),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

NAND4xp25_ASAP7_75t_SL g79 ( 
.A(n_76),
.B(n_72),
.C(n_71),
.D(n_73),
.Y(n_79)
);

NOR2xp67_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_75),
.Y(n_81)
);

NOR2xp67_ASAP7_75t_SL g82 ( 
.A(n_79),
.B(n_58),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_62),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

OAI22x1_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_50),
.B1(n_62),
.B2(n_66),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_87),
.A2(n_41),
.B1(n_67),
.B2(n_86),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_85),
.B(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_88),
.Y(n_91)
);


endmodule