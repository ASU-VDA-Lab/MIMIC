module fake_jpeg_17406_n_95 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_95);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_95;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx10_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_5),
.B(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_12),
.B(n_19),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_10),
.C(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_41),
.Y(n_49)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_45),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_17),
.B1(n_16),
.B2(n_18),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_42),
.B1(n_46),
.B2(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_17),
.B1(n_12),
.B2(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_56),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_36),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_54),
.B1(n_12),
.B2(n_27),
.Y(n_65)
);

CKINVDCx11_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_47),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_36),
.B1(n_21),
.B2(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_20),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_42),
.C(n_39),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_61),
.C(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_15),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_31),
.C(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_16),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_1),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_51),
.B1(n_50),
.B2(n_19),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_22),
.B1(n_25),
.B2(n_31),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_11),
.B(n_10),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_72),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_10),
.B(n_32),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_10),
.B(n_3),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_22),
.B1(n_5),
.B2(n_7),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_78),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_SL g80 ( 
.A(n_76),
.B(n_70),
.C(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_25),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_74),
.B1(n_77),
.B2(n_9),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_85),
.B(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_83),
.B(n_9),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_81),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_26),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_88),
.A2(n_82),
.B(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_91),
.Y(n_93)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_85),
.C(n_26),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_93),
.Y(n_95)
);


endmodule