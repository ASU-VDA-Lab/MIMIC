module fake_jpeg_4943_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_33),
.Y(n_38)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_39),
.B(n_41),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_16),
.B(n_14),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_44),
.B(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_13),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_48),
.Y(n_64)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_53),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_0),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_37),
.Y(n_83)
);

CKINVDCx9p33_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_62),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_30),
.B1(n_21),
.B2(n_28),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_59),
.A2(n_34),
.B1(n_37),
.B2(n_36),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_93),
.Y(n_110)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_46),
.B1(n_30),
.B2(n_52),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_65),
.A2(n_90),
.B1(n_26),
.B2(n_27),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_30),
.B1(n_20),
.B2(n_19),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_77),
.B1(n_80),
.B2(n_24),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_29),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_67),
.Y(n_118)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_84),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_83),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_19),
.B1(n_17),
.B2(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_79),
.B(n_81),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_38),
.A2(n_20),
.B1(n_19),
.B2(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_86),
.Y(n_114)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_22),
.B(n_23),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_26),
.A3(n_27),
.B1(n_31),
.B2(n_35),
.Y(n_106)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_89),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_25),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_31),
.B1(n_25),
.B2(n_26),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

CKINVDCx12_ASAP7_75t_R g96 ( 
.A(n_51),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_98),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_25),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_43),
.A2(n_22),
.B1(n_23),
.B2(n_15),
.Y(n_99)
);

AO22x1_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_54),
.B1(n_47),
.B2(n_15),
.Y(n_133)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_37),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_57),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_31),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_107),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_106),
.A2(n_109),
.B(n_123),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_72),
.B(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_50),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_117),
.Y(n_148)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_50),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

OR2x4_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_51),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_57),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_130),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_135),
.B1(n_101),
.B2(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_24),
.Y(n_130)
);

OA21x2_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_92),
.B(n_54),
.Y(n_152)
);

OR2x2_ASAP7_75t_SL g136 ( 
.A(n_73),
.B(n_12),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_24),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_34),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_99),
.B1(n_84),
.B2(n_94),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_138),
.A2(n_167),
.B1(n_5),
.B2(n_7),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_139),
.A2(n_140),
.B1(n_152),
.B2(n_157),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_99),
.B1(n_73),
.B2(n_94),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_122),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_141),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_99),
.B1(n_78),
.B2(n_75),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_144),
.B1(n_164),
.B2(n_171),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_78),
.B1(n_75),
.B2(n_92),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_147),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_86),
.C(n_70),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_150),
.C(n_111),
.Y(n_181)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_107),
.A2(n_93),
.A3(n_91),
.B1(n_70),
.B2(n_36),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_111),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_103),
.C(n_62),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_153),
.B(n_155),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_74),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_170),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_110),
.B1(n_132),
.B2(n_135),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_110),
.A2(n_88),
.B1(n_100),
.B2(n_104),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_158),
.A2(n_163),
.B1(n_165),
.B2(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_161),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_54),
.B1(n_36),
.B2(n_34),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_120),
.B1(n_137),
.B2(n_131),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_97),
.B1(n_95),
.B2(n_15),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_124),
.A2(n_23),
.B1(n_35),
.B2(n_58),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_169),
.B(n_127),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_74),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_118),
.A2(n_35),
.B1(n_23),
.B2(n_10),
.Y(n_171)
);

AOI22x1_ASAP7_75t_L g172 ( 
.A1(n_114),
.A2(n_85),
.B1(n_74),
.B2(n_60),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_60),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_173),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_126),
.A2(n_74),
.B(n_2),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_174),
.A2(n_10),
.B(n_12),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_136),
.B(n_118),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_178),
.A2(n_190),
.B(n_192),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_179),
.B(n_197),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_187),
.C(n_188),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_172),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_186),
.Y(n_227)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_116),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_SL g222 ( 
.A(n_184),
.B(n_142),
.C(n_154),
.Y(n_222)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_128),
.C(n_116),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_128),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_134),
.B(n_2),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_0),
.B(n_2),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g193 ( 
.A(n_142),
.B(n_0),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_204),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_8),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_202),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_0),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_206),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_150),
.B(n_127),
.C(n_119),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_141),
.B(n_8),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_149),
.B(n_8),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_138),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_209),
.B1(n_165),
.B2(n_162),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_145),
.B(n_3),
.C(n_4),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_151),
.B(n_3),
.C(n_5),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_12),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_163),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_229),
.B1(n_212),
.B2(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_213),
.B(n_214),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_159),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_217),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_193),
.B(n_153),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_203),
.A2(n_152),
.B1(n_167),
.B2(n_142),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_190),
.B(n_178),
.Y(n_243)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

AO221x1_ASAP7_75t_L g241 ( 
.A1(n_223),
.A2(n_224),
.B1(n_230),
.B2(n_236),
.C(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_203),
.A2(n_152),
.B1(n_169),
.B2(n_155),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_174),
.B1(n_147),
.B2(n_166),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_189),
.A2(n_168),
.B1(n_161),
.B2(n_7),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_180),
.B(n_13),
.Y(n_232)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_193),
.B(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_176),
.Y(n_235)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_181),
.C(n_188),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_240),
.C(n_245),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_187),
.C(n_200),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_223),
.B1(n_234),
.B2(n_183),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_208),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_191),
.C(n_207),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_228),
.B1(n_225),
.B2(n_229),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_194),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_250),
.C(n_254),
.Y(n_263)
);

OAI322xp33_ASAP7_75t_L g249 ( 
.A1(n_225),
.A2(n_212),
.A3(n_222),
.B1(n_230),
.B2(n_215),
.C1(n_232),
.C2(n_211),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_220),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_191),
.C(n_197),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_206),
.C(n_209),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_192),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_215),
.C(n_236),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_259),
.B(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_219),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_213),
.Y(n_266)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_272),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_268),
.A2(n_270),
.B(n_273),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_271),
.C(n_274),
.Y(n_285)
);

AOI22x1_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_183),
.B1(n_225),
.B2(n_231),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_226),
.C(n_224),
.Y(n_271)
);

BUFx12f_ASAP7_75t_SL g273 ( 
.A(n_258),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_219),
.C(n_205),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_242),
.A2(n_210),
.B1(n_182),
.B2(n_201),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_275),
.A2(n_251),
.B1(n_237),
.B2(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_276),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_256),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_263),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_286),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_237),
.B1(n_242),
.B2(n_250),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_287),
.B(n_254),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_248),
.C(n_245),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_262),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_272),
.A2(n_243),
.B1(n_239),
.B2(n_247),
.Y(n_289)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_289),
.Y(n_295)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_267),
.B(n_269),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_292),
.B(n_286),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_283),
.B(n_239),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_298),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_288),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_274),
.B1(n_263),
.B2(n_247),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_285),
.B1(n_276),
.B2(n_279),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_201),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_182),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_299),
.B(n_301),
.Y(n_305)
);

AO21x1_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_295),
.B(n_300),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_306),
.C(n_307),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_285),
.C(n_284),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_290),
.B(n_289),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_310),
.B(n_295),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_281),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_301),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_312),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_304),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_294),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_316),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_317),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_281),
.B(n_309),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_SL g320 ( 
.A(n_315),
.B(n_302),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_310),
.C(n_319),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_311),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_323),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_318),
.Y(n_325)
);


endmodule