module fake_netlist_1_12052_n_37 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
AND2x4_ASAP7_75t_L g15 ( .A(n_3), .B(n_2), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_2), .B(n_5), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_12), .B(n_0), .Y(n_18) );
OAI22xp33_ASAP7_75t_L g19 ( .A1(n_12), .A2(n_0), .B1(n_1), .B2(n_4), .Y(n_19) );
AOI22xp5_ASAP7_75t_L g20 ( .A1(n_15), .A2(n_1), .B1(n_4), .B2(n_5), .Y(n_20) );
BUFx6f_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g22 ( .A(n_18), .B(n_13), .Y(n_22) );
INVxp67_ASAP7_75t_SL g23 ( .A(n_20), .Y(n_23) );
AO31x2_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_13), .A3(n_14), .B(n_15), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_19), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_24), .B(n_23), .Y(n_26) );
NAND2xp33_ASAP7_75t_L g27 ( .A(n_25), .B(n_16), .Y(n_27) );
OAI31xp33_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_15), .A3(n_16), .B(n_14), .Y(n_28) );
AOI21xp5_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_15), .B(n_13), .Y(n_29) );
OAI221xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_14), .B1(n_17), .B2(n_24), .C(n_21), .Y(n_30) );
OAI21xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_6), .B(n_7), .Y(n_31) );
AND2x4_ASAP7_75t_L g32 ( .A(n_31), .B(n_6), .Y(n_32) );
OAI22xp5_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_17), .B1(n_21), .B2(n_9), .Y(n_33) );
OA22x2_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_7), .B1(n_8), .B2(n_11), .Y(n_34) );
OAI22xp5_ASAP7_75t_SL g35 ( .A1(n_33), .A2(n_17), .B1(n_8), .B2(n_11), .Y(n_35) );
HB1xp67_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
NAND2xp5_ASAP7_75t_L g37 ( .A(n_36), .B(n_35), .Y(n_37) );
endmodule