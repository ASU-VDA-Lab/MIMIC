module fake_jpeg_1845_n_571 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_571);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_571;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_55),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_9),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_56),
.B(n_66),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_58),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_61),
.Y(n_127)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_65),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_18),
.B(n_8),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_73),
.Y(n_112)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g121 ( 
.A(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_26),
.B(n_10),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_96),
.Y(n_125)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_52),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_76),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_79),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_31),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_85),
.Y(n_163)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_34),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_102),
.Y(n_142)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_25),
.B(n_1),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_26),
.B(n_10),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_100),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_44),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_103),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_25),
.B(n_1),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_34),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_44),
.B(n_1),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_107),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_47),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_41),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_27),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_109),
.B(n_23),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_27),
.B1(n_41),
.B2(n_43),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_116),
.A2(n_133),
.B1(n_144),
.B2(n_99),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_105),
.A2(n_27),
.B1(n_33),
.B2(n_50),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_120),
.A2(n_128),
.B1(n_138),
.B2(n_143),
.Y(n_232)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_76),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_100),
.A2(n_53),
.B1(n_39),
.B2(n_40),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_83),
.A2(n_33),
.B1(n_104),
.B2(n_60),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_54),
.B(n_43),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_140),
.B(n_150),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_72),
.A2(n_33),
.B1(n_51),
.B2(n_50),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_101),
.A2(n_107),
.B1(n_106),
.B2(n_89),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_95),
.A2(n_23),
.B1(n_51),
.B2(n_50),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_147),
.A2(n_151),
.B1(n_157),
.B2(n_173),
.Y(n_239)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_103),
.B(n_35),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_95),
.A2(n_21),
.B1(n_51),
.B2(n_46),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_59),
.B(n_53),
.C(n_40),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_153),
.B(n_49),
.C(n_30),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_97),
.A2(n_19),
.B1(n_46),
.B2(n_21),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_103),
.A2(n_35),
.B1(n_46),
.B2(n_37),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_28),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_61),
.B(n_39),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_169),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_62),
.B(n_32),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_86),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_171),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_97),
.A2(n_19),
.B1(n_37),
.B2(n_32),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_87),
.A2(n_19),
.B1(n_37),
.B2(n_32),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_178),
.B1(n_90),
.B2(n_79),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_65),
.B(n_23),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_74),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_177),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_88),
.A2(n_21),
.B1(n_28),
.B2(n_49),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_179),
.B(n_208),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_180),
.Y(n_255)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_91),
.B1(n_71),
.B2(n_84),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_182),
.A2(n_185),
.B1(n_212),
.B2(n_216),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_125),
.B(n_93),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_183),
.B(n_197),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_135),
.A2(n_67),
.B1(n_85),
.B2(n_80),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_184),
.A2(n_236),
.B1(n_163),
.B2(n_158),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_133),
.B(n_64),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_187),
.B(n_209),
.Y(n_245)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_189),
.Y(n_274)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_190),
.Y(n_275)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_191),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_110),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_192),
.B(n_199),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_193),
.B(n_206),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_195),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_134),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_196),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_123),
.B(n_109),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_198),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_112),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_200),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_201),
.Y(n_263)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_202),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_203),
.Y(n_294)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_205),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_117),
.B(n_69),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_63),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_207),
.B(n_214),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_152),
.B(n_1),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_141),
.Y(n_211)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_211),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_165),
.A2(n_152),
.B1(n_159),
.B2(n_77),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_152),
.B(n_1),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_227),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_139),
.B(n_114),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_175),
.B(n_82),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g279 ( 
.A1(n_215),
.A2(n_237),
.B(n_30),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_159),
.A2(n_78),
.B1(n_82),
.B2(n_49),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_118),
.B(n_74),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_217),
.B(n_219),
.Y(n_304)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_177),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_149),
.Y(n_221)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_221),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_81),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_222),
.Y(n_291)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_146),
.Y(n_224)
);

INVx5_ASAP7_75t_SL g249 ( 
.A(n_224),
.Y(n_249)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_154),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_225),
.B(n_228),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_128),
.A2(n_81),
.B(n_70),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_226),
.A2(n_229),
.B(n_235),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_132),
.B(n_3),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_166),
.A2(n_94),
.B(n_30),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_121),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_230),
.Y(n_261)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_231),
.A2(n_234),
.B1(n_113),
.B2(n_129),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_132),
.B(n_3),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_5),
.Y(n_257)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_161),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_128),
.A2(n_24),
.B(n_49),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_159),
.A2(n_164),
.B1(n_145),
.B2(n_162),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_121),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_155),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_30),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_241),
.C(n_113),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_155),
.B(n_4),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_164),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_242),
.Y(n_289)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_163),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_244),
.Y(n_292)
);

AO21x1_ASAP7_75t_SL g246 ( 
.A1(n_226),
.A2(n_128),
.B(n_121),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_246),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_185),
.A2(n_115),
.B1(n_122),
.B2(n_149),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_253),
.A2(n_260),
.B1(n_270),
.B2(n_276),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_256),
.B(n_283),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_257),
.B(n_295),
.Y(n_309)
);

AO22x1_ASAP7_75t_L g258 ( 
.A1(n_210),
.A2(n_124),
.B1(n_137),
.B2(n_167),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_258),
.B(n_286),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_187),
.A2(n_115),
.B1(n_122),
.B2(n_158),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_265),
.A2(n_191),
.B1(n_189),
.B2(n_196),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_130),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_268),
.B(n_277),
.C(n_278),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_235),
.A2(n_130),
.B1(n_124),
.B2(n_137),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_271),
.A2(n_281),
.B1(n_244),
.B2(n_196),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_232),
.A2(n_146),
.B1(n_172),
.B2(n_119),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_210),
.B(n_172),
.C(n_119),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_188),
.B(n_119),
.C(n_111),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_279),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_299),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_184),
.A2(n_49),
.B1(n_126),
.B2(n_30),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_222),
.B(n_111),
.C(n_126),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_227),
.B(n_5),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_12),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_222),
.B(n_111),
.C(n_126),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_179),
.A2(n_49),
.B1(n_111),
.B2(n_126),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_287),
.A2(n_288),
.B1(n_221),
.B2(n_198),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_239),
.A2(n_24),
.B1(n_6),
.B2(n_7),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_209),
.B(n_5),
.C(n_6),
.Y(n_295)
);

O2A1O1Ixp33_ASAP7_75t_SL g297 ( 
.A1(n_243),
.A2(n_7),
.B(n_10),
.C(n_11),
.Y(n_297)
);

A2O1A1O1Ixp25_ASAP7_75t_L g341 ( 
.A1(n_297),
.A2(n_12),
.B(n_13),
.C(n_14),
.D(n_15),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_243),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_213),
.A2(n_10),
.B(n_11),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_300),
.A2(n_229),
.B(n_241),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_220),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_307),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_308),
.A2(n_314),
.B(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_310),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_252),
.B(n_186),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_311),
.B(n_317),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_302),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_313),
.B(n_326),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_266),
.A2(n_233),
.B(n_241),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_304),
.B(n_236),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_315),
.B(n_339),
.Y(n_373)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_316),
.Y(n_363)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_247),
.B(n_181),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_319),
.B(n_324),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_320),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_321),
.A2(n_344),
.B1(n_347),
.B2(n_349),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_266),
.A2(n_202),
.B(n_231),
.Y(n_322)
);

OAI22x1_ASAP7_75t_L g323 ( 
.A1(n_246),
.A2(n_228),
.B1(n_218),
.B2(n_201),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_323),
.A2(n_249),
.B1(n_274),
.B2(n_290),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_247),
.B(n_190),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_302),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_328),
.A2(n_342),
.B1(n_345),
.B2(n_348),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_282),
.B(n_269),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_331),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_257),
.B(n_242),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_296),
.A2(n_234),
.B(n_194),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_343),
.B(n_350),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_245),
.B(n_225),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_333),
.B(n_334),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_248),
.B(n_195),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_302),
.Y(n_335)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_261),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_346),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_294),
.B(n_223),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_337),
.B(n_338),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_284),
.B(n_211),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_180),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_245),
.B(n_200),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_340),
.B(n_351),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_352),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_276),
.A2(n_296),
.B1(n_287),
.B2(n_288),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_296),
.A2(n_204),
.B(n_224),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_271),
.A2(n_200),
.B1(n_14),
.B2(n_15),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_292),
.A2(n_13),
.B1(n_15),
.B2(n_251),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_294),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_270),
.A2(n_13),
.B1(n_281),
.B2(n_291),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_256),
.A2(n_13),
.B1(n_277),
.B2(n_278),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_280),
.A2(n_300),
.B1(n_258),
.B2(n_273),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_297),
.A2(n_258),
.B(n_283),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_295),
.B(n_289),
.Y(n_351)
);

AOI22x1_ASAP7_75t_SL g352 ( 
.A1(n_254),
.A2(n_250),
.B1(n_286),
.B2(n_273),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_353),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_293),
.B(n_254),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_355),
.B(n_275),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_327),
.A2(n_303),
.B1(n_255),
.B2(n_264),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_356),
.A2(n_358),
.B1(n_375),
.B2(n_384),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_327),
.A2(n_303),
.B1(n_255),
.B2(n_264),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_312),
.B(n_267),
.C(n_272),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_364),
.C(n_367),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_310),
.Y(n_362)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_362),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_312),
.B(n_250),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_305),
.B(n_249),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_365),
.B(n_385),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_262),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_322),
.A2(n_263),
.B(n_274),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_376),
.A2(n_323),
.B(n_341),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_355),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_378),
.B(n_389),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_325),
.B(n_290),
.Y(n_381)
);

MAJx2_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_330),
.C(n_351),
.Y(n_407)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_383),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_306),
.A2(n_285),
.B1(n_262),
.B2(n_275),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_306),
.A2(n_285),
.B1(n_263),
.B2(n_259),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_386),
.A2(n_321),
.B1(n_335),
.B2(n_352),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_354),
.A2(n_259),
.B(n_305),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_388),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_311),
.B(n_307),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_339),
.B(n_348),
.C(n_354),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_391),
.B(n_338),
.C(n_308),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_337),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_315),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_329),
.B(n_334),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_394),
.B(n_346),
.Y(n_400)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_316),
.Y(n_395)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_395),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_314),
.A2(n_333),
.B1(n_330),
.B2(n_328),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_397),
.A2(n_347),
.B1(n_332),
.B2(n_343),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_400),
.B(n_423),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_349),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_401),
.A2(n_412),
.B1(n_414),
.B2(n_417),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_369),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_404),
.B(n_429),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_396),
.A2(n_350),
.B1(n_330),
.B2(n_340),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_406),
.A2(n_377),
.B1(n_392),
.B2(n_393),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_407),
.B(n_428),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_360),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_408),
.B(n_415),
.Y(n_455)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_410),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_324),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_413),
.B(n_428),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_309),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_359),
.Y(n_416)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_416),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_397),
.A2(n_323),
.B1(n_344),
.B2(n_319),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_359),
.Y(n_419)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_419),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_381),
.B(n_309),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_424),
.C(n_373),
.Y(n_435)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_363),
.Y(n_421)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_421),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_396),
.A2(n_352),
.B1(n_313),
.B2(n_326),
.Y(n_422)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_379),
.B(n_331),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_425),
.A2(n_376),
.B(n_366),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_368),
.A2(n_318),
.B1(n_317),
.B2(n_341),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_427),
.A2(n_375),
.B1(n_371),
.B2(n_390),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_364),
.B(n_391),
.Y(n_428)
);

FAx1_ASAP7_75t_SL g429 ( 
.A(n_357),
.B(n_366),
.CI(n_361),
.CON(n_429),
.SN(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_363),
.Y(n_430)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_430),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_365),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_434),
.Y(n_462)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_370),
.Y(n_432)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_432),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_371),
.B(n_374),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_433),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_365),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_437),
.C(n_451),
.Y(n_468)
);

XNOR2x1_ASAP7_75t_L g488 ( 
.A(n_436),
.B(n_419),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_403),
.B(n_357),
.C(n_378),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_410),
.Y(n_440)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_440),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_418),
.A2(n_377),
.B1(n_390),
.B2(n_398),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_444),
.B(n_445),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_418),
.A2(n_377),
.B(n_380),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_448),
.A2(n_432),
.B(n_430),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_387),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_449),
.B(n_461),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_403),
.B(n_380),
.C(n_372),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_411),
.Y(n_452)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_452),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_407),
.B(n_372),
.C(n_387),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_402),
.C(n_427),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_426),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_463),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_457),
.A2(n_416),
.B1(n_399),
.B2(n_426),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_424),
.B(n_393),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_412),
.A2(n_401),
.B1(n_417),
.B2(n_431),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_464),
.B(n_434),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_404),
.B(n_362),
.Y(n_465)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_465),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_455),
.B(n_409),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_466),
.B(n_473),
.Y(n_496)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_470),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_413),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_476),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_SL g472 ( 
.A(n_439),
.B(n_406),
.C(n_429),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_436),
.C(n_444),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_438),
.B(n_409),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_454),
.B(n_429),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_477),
.B(n_435),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_456),
.Y(n_479)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_479),
.Y(n_511)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_457),
.Y(n_499)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_446),
.B(n_402),
.C(n_399),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_482),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_SL g482 ( 
.A(n_439),
.B(n_425),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_462),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_483),
.B(n_485),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_484),
.A2(n_443),
.B(n_362),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_451),
.B(n_453),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_437),
.B(n_421),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_486),
.B(n_450),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_411),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_490),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_488),
.B(n_459),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_489),
.A2(n_464),
.B1(n_441),
.B2(n_460),
.Y(n_494)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_442),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_492),
.B(n_501),
.Y(n_526)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_494),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_480),
.A2(n_447),
.B1(n_463),
.B2(n_448),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_495),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_504),
.Y(n_519)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_499),
.Y(n_523)
);

XOR2x2_ASAP7_75t_L g501 ( 
.A(n_477),
.B(n_449),
.Y(n_501)
);

AO22x1_ASAP7_75t_L g502 ( 
.A1(n_475),
.A2(n_445),
.B1(n_405),
.B2(n_452),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_502),
.B(n_509),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_479),
.B(n_443),
.Y(n_503)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_503),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_458),
.Y(n_507)
);

CKINVDCx14_ASAP7_75t_R g524 ( 
.A(n_507),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_508),
.B(n_474),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_467),
.A2(n_356),
.B1(n_358),
.B2(n_442),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_510),
.A2(n_484),
.B(n_470),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_370),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_512),
.B(n_513),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_468),
.B(n_395),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_515),
.A2(n_510),
.B(n_493),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_497),
.B(n_468),
.C(n_469),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_516),
.B(n_517),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_497),
.B(n_469),
.C(n_471),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_498),
.B(n_472),
.C(n_491),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_520),
.B(n_501),
.C(n_504),
.Y(n_536)
);

FAx1_ASAP7_75t_SL g522 ( 
.A(n_492),
.B(n_488),
.CI(n_489),
.CON(n_522),
.SN(n_522)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_522),
.B(n_525),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_491),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_527),
.B(n_525),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_503),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_528),
.B(n_531),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_496),
.B(n_467),
.Y(n_531)
);

NOR2xp67_ASAP7_75t_L g532 ( 
.A(n_529),
.B(n_505),
.Y(n_532)
);

NOR3xp33_ASAP7_75t_L g550 ( 
.A(n_532),
.B(n_534),
.C(n_542),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_533),
.B(n_539),
.Y(n_548)
);

XOR2x1_ASAP7_75t_SL g534 ( 
.A(n_527),
.B(n_491),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_518),
.A2(n_493),
.B1(n_502),
.B2(n_475),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_535),
.A2(n_511),
.B1(n_521),
.B2(n_502),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_536),
.B(n_543),
.Y(n_547)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_530),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_541),
.A2(n_545),
.B(n_522),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_516),
.B(n_500),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_517),
.B(n_514),
.C(n_520),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_524),
.B(n_506),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_544),
.B(n_523),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_515),
.A2(n_495),
.B(n_499),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_546),
.B(n_549),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_540),
.A2(n_526),
.B(n_521),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_537),
.B(n_543),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_551),
.B(n_552),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_538),
.B(n_494),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_553),
.B(n_554),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_535),
.A2(n_511),
.B1(n_478),
.B2(n_522),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_555),
.A2(n_540),
.B(n_545),
.Y(n_557)
);

XNOR2x1_ASAP7_75t_L g556 ( 
.A(n_548),
.B(n_536),
.Y(n_556)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_556),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_557),
.B(n_558),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_547),
.B(n_546),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_559),
.B(n_550),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_563),
.A2(n_562),
.B(n_565),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_560),
.B(n_541),
.C(n_534),
.Y(n_564)
);

AOI21x1_ASAP7_75t_L g566 ( 
.A1(n_564),
.A2(n_561),
.B(n_519),
.Y(n_566)
);

NAND4xp25_ASAP7_75t_L g568 ( 
.A(n_566),
.B(n_567),
.C(n_561),
.D(n_519),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_382),
.C(n_383),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_382),
.B(n_386),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_570),
.B(n_384),
.Y(n_571)
);


endmodule