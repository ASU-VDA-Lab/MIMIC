module fake_jpeg_2794_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_6),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_4),
.B(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

AOI32xp33_ASAP7_75t_L g16 ( 
.A1(n_13),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_14),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_9),
.B1(n_8),
.B2(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_24),
.C(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_26),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_12),
.B1(n_8),
.B2(n_7),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_27),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_17),
.A2(n_19),
.B1(n_16),
.B2(n_22),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_23),
.B(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_32),
.B(n_30),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_29),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_39),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_37),
.B1(n_38),
.B2(n_29),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_41),
.B1(n_40),
.B2(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_38),
.Y(n_47)
);


endmodule