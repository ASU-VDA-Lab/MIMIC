module fake_aes_9883_n_1014 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1014);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1014;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_918;
wire n_770;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_529;
wire n_312;
wire n_1011;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_274;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_935;
wire n_460;
wire n_478;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_805;
wire n_699;
wire n_729;
wire n_693;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_703;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_716;
wire n_653;
wire n_899;
wire n_806;
wire n_881;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_429;
wire n_488;
wire n_763;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_912;
wire n_620;
wire n_841;
wire n_924;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_859;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_120), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_216), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_77), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_110), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_225), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_97), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_235), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_40), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_269), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_154), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_167), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_87), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_150), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_70), .Y(n_283) );
BUFx2_ASAP7_75t_SL g284 ( .A(n_55), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_52), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_21), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_265), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_133), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_64), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_243), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_219), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_68), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_132), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_183), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_12), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_224), .Y(n_296) );
BUFx2_ASAP7_75t_SL g297 ( .A(n_220), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_36), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_147), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_145), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_244), .B(n_184), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_149), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_4), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_82), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_20), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_91), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_79), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_227), .Y(n_308) );
INVxp67_ASAP7_75t_SL g309 ( .A(n_6), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_236), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_107), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_81), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_23), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_61), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_234), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_189), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_123), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_112), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_232), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_127), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_38), .Y(n_321) );
INVx1_ASAP7_75t_SL g322 ( .A(n_177), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_139), .Y(n_323) );
INVxp67_ASAP7_75t_L g324 ( .A(n_7), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_247), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_20), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_138), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_163), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_146), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_80), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_56), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_258), .Y(n_332) );
BUFx2_ASAP7_75t_SL g333 ( .A(n_41), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_45), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_245), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_267), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_136), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_214), .Y(n_338) );
INVxp67_ASAP7_75t_SL g339 ( .A(n_32), .Y(n_339) );
BUFx5_ASAP7_75t_L g340 ( .A(n_54), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_59), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_57), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_42), .Y(n_343) );
BUFx10_ASAP7_75t_L g344 ( .A(n_206), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_90), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_246), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_129), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_212), .Y(n_348) );
CKINVDCx16_ASAP7_75t_R g349 ( .A(n_179), .Y(n_349) );
CKINVDCx16_ASAP7_75t_R g350 ( .A(n_142), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_11), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_239), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_63), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_203), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_255), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_23), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_30), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_173), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_125), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_230), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_88), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_94), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_126), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_84), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_164), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_16), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_134), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_217), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_121), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_152), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_28), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_95), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_135), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_187), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_86), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_108), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_21), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_250), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_8), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_43), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_259), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_175), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_124), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_12), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_155), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_160), .Y(n_386) );
INVx2_ASAP7_75t_SL g387 ( .A(n_196), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_83), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_223), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_193), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_102), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_118), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_256), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_172), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_89), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_192), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_171), .Y(n_397) );
INVxp67_ASAP7_75t_L g398 ( .A(n_176), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_202), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_174), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_211), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_14), .Y(n_402) );
INVx1_ASAP7_75t_SL g403 ( .A(n_27), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_109), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_252), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_384), .B(n_0), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_349), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_350), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_340), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_274), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_340), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_305), .B(n_1), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_340), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_302), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_362), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_340), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_405), .Y(n_417) );
INVx5_ASAP7_75t_L g418 ( .A(n_306), .Y(n_418) );
OAI21x1_ASAP7_75t_L g419 ( .A1(n_317), .A2(n_31), .B(n_29), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_306), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_351), .Y(n_421) );
AOI22xp5_ASAP7_75t_SL g422 ( .A1(n_366), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_340), .B(n_3), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_326), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_344), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_320), .Y(n_426) );
INVx3_ASAP7_75t_L g427 ( .A(n_344), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_276), .B(n_5), .Y(n_428) );
OAI21x1_ASAP7_75t_L g429 ( .A1(n_329), .A2(n_34), .B(n_33), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_381), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_330), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_295), .B(n_8), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_286), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_356), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_379), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_394), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_432), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_425), .B(n_335), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_432), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_409), .B(n_401), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_425), .B(n_427), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_432), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_410), .Y(n_443) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_420), .Y(n_444) );
INVx2_ASAP7_75t_SL g445 ( .A(n_425), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_409), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_410), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_427), .B(n_387), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_411), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_413), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_413), .B(n_404), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_416), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_416), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_426), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_408), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_426), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
AOI21x1_ASAP7_75t_L g459 ( .A1(n_419), .A2(n_275), .B(n_271), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_408), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_420), .Y(n_461) );
INVx4_ASAP7_75t_L g462 ( .A(n_428), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_420), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_420), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_421), .B(n_324), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_462), .B(n_428), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_462), .B(n_428), .Y(n_467) );
NAND2xp33_ASAP7_75t_L g468 ( .A(n_439), .B(n_301), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_462), .B(n_414), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_441), .B(n_415), .Y(n_470) );
INVx3_ASAP7_75t_L g471 ( .A(n_449), .Y(n_471) );
NAND2xp33_ASAP7_75t_SL g472 ( .A(n_456), .B(n_323), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_445), .B(n_427), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_445), .B(n_417), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_437), .B(n_430), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_437), .B(n_434), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_437), .B(n_406), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_465), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_442), .B(n_435), .Y(n_479) );
NOR2x2_ASAP7_75t_L g480 ( .A(n_443), .B(n_422), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_448), .B(n_412), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_442), .B(n_431), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_442), .B(n_431), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_438), .B(n_436), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_454), .A2(n_423), .B1(n_436), .B2(n_407), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_455), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_460), .B(n_270), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_446), .A2(n_423), .B1(n_286), .B2(n_303), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_447), .Y(n_489) );
NAND2x1p5_ASAP7_75t_L g490 ( .A(n_440), .B(n_419), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_449), .B(n_272), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_440), .A2(n_328), .B1(n_369), .B2(n_325), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_449), .B(n_446), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_450), .B(n_273), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_457), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_452), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_450), .B(n_374), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_451), .A2(n_286), .B1(n_303), .B2(n_309), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_451), .B(n_398), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_453), .B(n_398), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_471), .Y(n_501) );
OR2x6_ASAP7_75t_L g502 ( .A(n_489), .B(n_284), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_466), .A2(n_453), .B(n_429), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_490), .A2(n_459), .B(n_429), .Y(n_504) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_471), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_477), .A2(n_339), .B(n_281), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_476), .A2(n_282), .B(n_279), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_470), .A2(n_392), .B1(n_424), .B2(n_443), .Y(n_508) );
BUFx4f_ASAP7_75t_L g509 ( .A(n_467), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_478), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_481), .A2(n_283), .B(n_288), .C(n_287), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_495), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_469), .B(n_313), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_469), .B(n_377), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_492), .A2(n_402), .B1(n_396), .B2(n_322), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_479), .A2(n_296), .B(n_294), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_468), .B(n_310), .C(n_298), .Y(n_517) );
NOR3xp33_ASAP7_75t_L g518 ( .A(n_472), .B(n_396), .C(n_322), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_468), .A2(n_311), .B(n_318), .C(n_314), .Y(n_519) );
OAI21xp33_ASAP7_75t_SL g520 ( .A1(n_495), .A2(n_321), .B(n_319), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_482), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_467), .B(n_403), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_474), .B(n_403), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_483), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_475), .A2(n_486), .B(n_499), .C(n_497), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_493), .A2(n_337), .B(n_334), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_485), .B(n_277), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_472), .A2(n_346), .B1(n_347), .B2(n_345), .Y(n_528) );
INVx3_ASAP7_75t_SL g529 ( .A(n_480), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_487), .B(n_278), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_490), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_484), .A2(n_352), .B1(n_353), .B2(n_348), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_500), .B(n_285), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_496), .A2(n_355), .B(n_354), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_473), .A2(n_360), .B(n_359), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_490), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_498), .Y(n_537) );
AO31x2_ASAP7_75t_L g538 ( .A1(n_531), .A2(n_364), .A3(n_365), .B(n_363), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_510), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_503), .A2(n_494), .B(n_491), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_512), .Y(n_541) );
AOI21x1_ASAP7_75t_L g542 ( .A1(n_504), .A2(n_370), .B(n_368), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_509), .B(n_488), .Y(n_543) );
AO21x1_ASAP7_75t_L g544 ( .A1(n_525), .A2(n_373), .B(n_372), .Y(n_544) );
BUFx12f_ASAP7_75t_L g545 ( .A(n_502), .Y(n_545) );
NAND2x1_ASAP7_75t_L g546 ( .A(n_505), .B(n_306), .Y(n_546) );
AO31x2_ASAP7_75t_L g547 ( .A1(n_536), .A2(n_385), .A3(n_391), .B(n_376), .Y(n_547) );
OAI21x1_ASAP7_75t_L g548 ( .A1(n_501), .A2(n_399), .B(n_397), .Y(n_548) );
CKINVDCx8_ASAP7_75t_R g549 ( .A(n_502), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_SL g550 ( .A1(n_511), .A2(n_400), .B(n_464), .C(n_463), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_521), .A2(n_461), .B(n_458), .Y(n_551) );
CKINVDCx11_ASAP7_75t_R g552 ( .A(n_529), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_524), .A2(n_464), .B(n_463), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_502), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_SL g555 ( .A1(n_519), .A2(n_433), .B(n_333), .C(n_297), .Y(n_555) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_526), .A2(n_433), .B(n_342), .Y(n_556) );
BUFx2_ASAP7_75t_L g557 ( .A(n_509), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_537), .B(n_280), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_508), .B(n_480), .Y(n_559) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_507), .A2(n_433), .B(n_342), .Y(n_560) );
AO31x2_ASAP7_75t_L g561 ( .A1(n_532), .A2(n_342), .A3(n_332), .B(n_371), .Y(n_561) );
OAI21xp5_ASAP7_75t_L g562 ( .A1(n_516), .A2(n_290), .B(n_289), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g563 ( .A1(n_520), .A2(n_336), .B(n_393), .C(n_316), .Y(n_563) );
OAI21x1_ASAP7_75t_L g564 ( .A1(n_534), .A2(n_371), .B(n_332), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_527), .A2(n_292), .B(n_291), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_523), .B(n_303), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_513), .B(n_9), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_505), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_520), .A2(n_332), .B(n_371), .C(n_390), .Y(n_569) );
AOI21xp5_ASAP7_75t_SL g570 ( .A1(n_505), .A2(n_390), .B(n_299), .Y(n_570) );
OAI21xp5_ASAP7_75t_SL g571 ( .A1(n_517), .A2(n_390), .B(n_9), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_528), .B(n_418), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_522), .B(n_293), .Y(n_573) );
A2O1A1Ixp33_ASAP7_75t_L g574 ( .A1(n_506), .A2(n_358), .B(n_304), .C(n_395), .Y(n_574) );
OAI21x1_ASAP7_75t_L g575 ( .A1(n_535), .A2(n_37), .B(n_35), .Y(n_575) );
AO21x1_ASAP7_75t_L g576 ( .A1(n_518), .A2(n_44), .B(n_39), .Y(n_576) );
AOI221xp5_ASAP7_75t_SL g577 ( .A1(n_515), .A2(n_444), .B1(n_11), .B2(n_13), .C(n_14), .Y(n_577) );
BUFx2_ASAP7_75t_L g578 ( .A(n_514), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_530), .B(n_10), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_533), .A2(n_307), .B(n_300), .Y(n_580) );
OA21x2_ASAP7_75t_L g581 ( .A1(n_542), .A2(n_312), .B(n_308), .Y(n_581) );
AOI21xp5_ASAP7_75t_SL g582 ( .A1(n_569), .A2(n_327), .B(n_315), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_539), .B(n_10), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_540), .A2(n_444), .B(n_418), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_541), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_541), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_578), .B(n_13), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_545), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_567), .B(n_558), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_566), .Y(n_590) );
OAI21x1_ASAP7_75t_L g591 ( .A1(n_560), .A2(n_444), .B(n_418), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_561), .Y(n_592) );
OAI21x1_ASAP7_75t_L g593 ( .A1(n_556), .A2(n_418), .B(n_47), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_538), .Y(n_594) );
OAI21xp5_ASAP7_75t_L g595 ( .A1(n_563), .A2(n_418), .B(n_338), .Y(n_595) );
INVx3_ASAP7_75t_L g596 ( .A(n_549), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_555), .A2(n_341), .B(n_331), .Y(n_597) );
BUFx12f_ASAP7_75t_L g598 ( .A(n_552), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_558), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_561), .Y(n_600) );
AO21x2_ASAP7_75t_L g601 ( .A1(n_544), .A2(n_48), .B(n_46), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_579), .B(n_15), .Y(n_602) );
AO21x2_ASAP7_75t_L g603 ( .A1(n_571), .A2(n_50), .B(n_49), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_538), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_561), .Y(n_605) );
BUFx2_ASAP7_75t_L g606 ( .A(n_557), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_538), .Y(n_607) );
OAI21x1_ASAP7_75t_L g608 ( .A1(n_564), .A2(n_53), .B(n_51), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_550), .A2(n_357), .B(n_343), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_551), .A2(n_367), .B(n_361), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_559), .A2(n_389), .B1(n_388), .B2(n_386), .Y(n_611) );
OR2x6_ASAP7_75t_L g612 ( .A(n_570), .B(n_15), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_547), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_547), .Y(n_614) );
OAI21xp5_ASAP7_75t_L g615 ( .A1(n_577), .A2(n_383), .B(n_382), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_553), .A2(n_380), .B(n_378), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_547), .Y(n_617) );
AO21x2_ASAP7_75t_L g618 ( .A1(n_571), .A2(n_162), .B(n_268), .Y(n_618) );
OA21x2_ASAP7_75t_L g619 ( .A1(n_548), .A2(n_375), .B(n_161), .Y(n_619) );
OAI21x1_ASAP7_75t_L g620 ( .A1(n_575), .A2(n_159), .B(n_264), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_554), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_573), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_622) );
AO21x2_ASAP7_75t_L g623 ( .A1(n_576), .A2(n_158), .B(n_263), .Y(n_623) );
NOR2x1_ASAP7_75t_SL g624 ( .A(n_568), .B(n_17), .Y(n_624) );
BUFx2_ASAP7_75t_L g625 ( .A(n_572), .Y(n_625) );
OAI21x1_ASAP7_75t_L g626 ( .A1(n_546), .A2(n_165), .B(n_262), .Y(n_626) );
AOI21xp5_ASAP7_75t_SL g627 ( .A1(n_574), .A2(n_157), .B(n_261), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_543), .Y(n_628) );
BUFx3_ASAP7_75t_L g629 ( .A(n_565), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_562), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_580), .A2(n_156), .B(n_260), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_539), .B(n_18), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_569), .A2(n_19), .B(n_22), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_541), .Y(n_634) );
NAND2x1p5_ASAP7_75t_L g635 ( .A(n_557), .B(n_19), .Y(n_635) );
BUFx8_ASAP7_75t_L g636 ( .A(n_545), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_541), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_540), .A2(n_166), .B(n_257), .Y(n_638) );
BUFx8_ASAP7_75t_L g639 ( .A(n_545), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_541), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_637), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_628), .B(n_22), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_585), .B(n_24), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_640), .B(n_25), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_586), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_634), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_625), .Y(n_647) );
BUFx2_ASAP7_75t_L g648 ( .A(n_606), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_632), .B(n_26), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_587), .B(n_26), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_600), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_635), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_589), .B(n_58), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_635), .Y(n_654) );
INVx1_ASAP7_75t_SL g655 ( .A(n_588), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_583), .Y(n_656) );
OA21x2_ASAP7_75t_L g657 ( .A1(n_605), .A2(n_60), .B(n_62), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_599), .B(n_65), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_624), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_589), .B(n_621), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_594), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_602), .Y(n_662) );
INVxp67_ASAP7_75t_SL g663 ( .A(n_594), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_630), .B(n_66), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_602), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_596), .B(n_266), .Y(n_666) );
AO21x2_ASAP7_75t_L g667 ( .A1(n_604), .A2(n_67), .B(n_69), .Y(n_667) );
AO21x1_ASAP7_75t_SL g668 ( .A1(n_633), .A2(n_71), .B(n_72), .Y(n_668) );
BUFx3_ASAP7_75t_L g669 ( .A(n_636), .Y(n_669) );
OR2x6_ASAP7_75t_L g670 ( .A(n_612), .B(n_73), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_622), .Y(n_671) );
INVx4_ASAP7_75t_L g672 ( .A(n_612), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_607), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_613), .Y(n_674) );
AO21x2_ASAP7_75t_L g675 ( .A1(n_614), .A2(n_74), .B(n_75), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_617), .Y(n_676) );
BUFx2_ASAP7_75t_L g677 ( .A(n_596), .Y(n_677) );
BUFx3_ASAP7_75t_L g678 ( .A(n_636), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_612), .B(n_76), .Y(n_679) );
AO21x2_ASAP7_75t_L g680 ( .A1(n_615), .A2(n_78), .B(n_85), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_620), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_590), .A2(n_92), .B1(n_93), .B2(n_96), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_591), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_633), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_593), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_603), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_629), .B(n_98), .Y(n_687) );
BUFx2_ASAP7_75t_L g688 ( .A(n_639), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_615), .B(n_99), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_603), .B(n_100), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_608), .Y(n_691) );
INVxp67_ASAP7_75t_L g692 ( .A(n_618), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_611), .B(n_595), .Y(n_693) );
INVx3_ASAP7_75t_L g694 ( .A(n_618), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_595), .B(n_101), .Y(n_695) );
AO21x2_ASAP7_75t_L g696 ( .A1(n_584), .A2(n_103), .B(n_104), .Y(n_696) );
INVx3_ASAP7_75t_L g697 ( .A(n_626), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_581), .B(n_610), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_619), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_619), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_601), .Y(n_701) );
AO21x2_ASAP7_75t_L g702 ( .A1(n_584), .A2(n_601), .B(n_623), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_623), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_638), .B(n_105), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_598), .B(n_106), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_631), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_631), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_639), .Y(n_708) );
INVx3_ASAP7_75t_L g709 ( .A(n_582), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_627), .Y(n_710) );
OA21x2_ASAP7_75t_L g711 ( .A1(n_638), .A2(n_111), .B(n_113), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_610), .B(n_114), .Y(n_712) );
AO21x2_ASAP7_75t_L g713 ( .A1(n_597), .A2(n_115), .B(n_116), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_609), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_609), .Y(n_715) );
CKINVDCx5p33_ASAP7_75t_R g716 ( .A(n_616), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_616), .Y(n_717) );
AO21x2_ASAP7_75t_L g718 ( .A1(n_592), .A2(n_117), .B(n_119), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_587), .B(n_122), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_628), .B(n_128), .Y(n_720) );
AO21x2_ASAP7_75t_L g721 ( .A1(n_592), .A2(n_130), .B(n_131), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_637), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_637), .Y(n_723) );
INVx5_ASAP7_75t_SL g724 ( .A(n_612), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_637), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_637), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_637), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_594), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_628), .A2(n_137), .B1(n_140), .B2(n_141), .Y(n_729) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_585), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_641), .Y(n_731) );
CKINVDCx5p33_ASAP7_75t_R g732 ( .A(n_669), .Y(n_732) );
AND2x4_ASAP7_75t_L g733 ( .A(n_672), .B(n_143), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_722), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_660), .B(n_144), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_723), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_656), .B(n_148), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_643), .B(n_151), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_648), .B(n_153), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_662), .B(n_168), .Y(n_740) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_730), .Y(n_741) );
BUFx3_ASAP7_75t_L g742 ( .A(n_669), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_665), .B(n_169), .Y(n_743) );
INVx2_ASAP7_75t_SL g744 ( .A(n_678), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_725), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_645), .Y(n_746) );
AND2x4_ASAP7_75t_L g747 ( .A(n_672), .B(n_170), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_726), .Y(n_748) );
INVx3_ASAP7_75t_L g749 ( .A(n_672), .Y(n_749) );
BUFx3_ASAP7_75t_L g750 ( .A(n_678), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_646), .B(n_178), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_727), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_643), .B(n_180), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_673), .Y(n_754) );
INVxp67_ASAP7_75t_SL g755 ( .A(n_663), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_674), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_676), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_684), .B(n_181), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_644), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_671), .A2(n_182), .B1(n_185), .B2(n_186), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_730), .Y(n_761) );
AND2x4_ASAP7_75t_L g762 ( .A(n_670), .B(n_188), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_647), .B(n_190), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_652), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_655), .B(n_191), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_708), .B(n_254), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_654), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_647), .B(n_194), .Y(n_768) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_663), .Y(n_769) );
NOR3xp33_ASAP7_75t_L g770 ( .A(n_659), .B(n_195), .C(n_197), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_661), .B(n_198), .Y(n_771) );
OR2x2_ASAP7_75t_L g772 ( .A(n_649), .B(n_199), .Y(n_772) );
AND2x4_ASAP7_75t_L g773 ( .A(n_670), .B(n_200), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_661), .B(n_201), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_677), .B(n_204), .Y(n_775) );
INVx3_ASAP7_75t_L g776 ( .A(n_670), .Y(n_776) );
AND2x4_ASAP7_75t_L g777 ( .A(n_728), .B(n_205), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_728), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_719), .B(n_207), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_650), .B(n_208), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_724), .B(n_209), .Y(n_781) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_724), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_642), .Y(n_783) );
AND2x4_ASAP7_75t_L g784 ( .A(n_679), .B(n_210), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_716), .B(n_213), .Y(n_785) );
AND2x4_ASAP7_75t_L g786 ( .A(n_687), .B(n_215), .Y(n_786) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_724), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_705), .B(n_218), .Y(n_788) );
OR2x2_ASAP7_75t_L g789 ( .A(n_688), .B(n_221), .Y(n_789) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_687), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_716), .B(n_253), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_653), .B(n_222), .Y(n_792) );
INVx5_ASAP7_75t_SL g793 ( .A(n_687), .Y(n_793) );
OR2x2_ASAP7_75t_L g794 ( .A(n_651), .B(n_251), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_666), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_653), .B(n_226), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_664), .Y(n_797) );
NOR2x1_ASAP7_75t_L g798 ( .A(n_667), .B(n_228), .Y(n_798) );
OR2x2_ASAP7_75t_L g799 ( .A(n_698), .B(n_229), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_720), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_658), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_714), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_712), .B(n_231), .Y(n_803) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_689), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_715), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_712), .B(n_233), .Y(n_806) );
INVxp67_ASAP7_75t_L g807 ( .A(n_668), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_689), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_693), .B(n_237), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_717), .B(n_238), .Y(n_810) );
OR2x2_ASAP7_75t_L g811 ( .A(n_706), .B(n_249), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_667), .Y(n_812) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_683), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_695), .B(n_240), .Y(n_814) );
NOR2x1_ASAP7_75t_L g815 ( .A(n_675), .B(n_710), .Y(n_815) );
BUFx3_ASAP7_75t_L g816 ( .A(n_709), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_657), .Y(n_817) );
OR2x2_ASAP7_75t_L g818 ( .A(n_707), .B(n_248), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_709), .B(n_241), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_657), .Y(n_820) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_690), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_709), .B(n_242), .Y(n_822) );
INVx3_ASAP7_75t_L g823 ( .A(n_690), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_746), .B(n_704), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_731), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_764), .B(n_686), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_752), .B(n_704), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_776), .A2(n_680), .B1(n_686), .B2(n_710), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_767), .B(n_692), .Y(n_829) );
NAND2x1p5_ASAP7_75t_L g830 ( .A(n_762), .B(n_711), .Y(n_830) );
OR2x2_ASAP7_75t_L g831 ( .A(n_778), .B(n_692), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_734), .B(n_696), .Y(n_832) );
BUFx2_ASAP7_75t_L g833 ( .A(n_742), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_736), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_754), .B(n_694), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_756), .B(n_757), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_802), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_745), .B(n_694), .Y(n_838) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_755), .Y(n_839) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_755), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_748), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_805), .B(n_694), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_769), .Y(n_843) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_769), .Y(n_844) );
AND2x4_ASAP7_75t_L g845 ( .A(n_823), .B(n_697), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_813), .Y(n_846) );
AND2x4_ASAP7_75t_L g847 ( .A(n_790), .B(n_697), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_808), .B(n_701), .Y(n_848) );
NAND2xp5_ASAP7_75t_SL g849 ( .A(n_793), .B(n_697), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_776), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_783), .B(n_680), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_813), .Y(n_852) );
INVx2_ASAP7_75t_L g853 ( .A(n_817), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_795), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_793), .B(n_696), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_759), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_797), .B(n_702), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_793), .B(n_702), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_821), .B(n_699), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_820), .Y(n_860) );
INVx4_ASAP7_75t_L g861 ( .A(n_786), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_804), .B(n_721), .Y(n_862) );
INVx3_ASAP7_75t_L g863 ( .A(n_790), .Y(n_863) );
AND2x4_ASAP7_75t_SL g864 ( .A(n_762), .B(n_729), .Y(n_864) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_741), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_801), .B(n_700), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_800), .B(n_729), .Y(n_867) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_790), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_735), .B(n_721), .Y(n_869) );
HB1xp67_ASAP7_75t_SL g870 ( .A(n_750), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_761), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_771), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_777), .B(n_718), .Y(n_873) );
OR2x2_ASAP7_75t_L g874 ( .A(n_744), .B(n_683), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_777), .B(n_718), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_771), .Y(n_876) );
NAND2xp5_ASAP7_75t_SL g877 ( .A(n_807), .B(n_681), .Y(n_877) );
OR2x2_ASAP7_75t_L g878 ( .A(n_739), .B(n_703), .Y(n_878) );
BUFx2_ASAP7_75t_L g879 ( .A(n_782), .Y(n_879) );
INVx3_ASAP7_75t_L g880 ( .A(n_816), .Y(n_880) );
INVx1_ASAP7_75t_SL g881 ( .A(n_732), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_774), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_815), .B(n_685), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_774), .Y(n_884) );
INVx3_ASAP7_75t_L g885 ( .A(n_749), .Y(n_885) );
NAND2x1_ASAP7_75t_L g886 ( .A(n_786), .B(n_773), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_738), .B(n_713), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_753), .B(n_787), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_794), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_836), .B(n_773), .Y(n_890) );
OR2x2_ASAP7_75t_L g891 ( .A(n_839), .B(n_799), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_836), .B(n_807), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_854), .B(n_785), .Y(n_893) );
NAND2x1p5_ASAP7_75t_L g894 ( .A(n_861), .B(n_747), .Y(n_894) );
OR2x2_ASAP7_75t_L g895 ( .A(n_839), .B(n_785), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_856), .B(n_791), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_835), .B(n_812), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_825), .B(n_809), .Y(n_898) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_840), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_835), .B(n_815), .Y(n_900) );
OR2x2_ASAP7_75t_L g901 ( .A(n_840), .B(n_789), .Y(n_901) );
OR2x2_ASAP7_75t_L g902 ( .A(n_844), .B(n_751), .Y(n_902) );
AND2x2_ASAP7_75t_L g903 ( .A(n_888), .B(n_784), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_833), .B(n_784), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_834), .B(n_809), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_841), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_844), .B(n_775), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_843), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_872), .B(n_737), .Y(n_909) );
BUFx2_ASAP7_75t_L g910 ( .A(n_861), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_850), .B(n_822), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_837), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_842), .B(n_810), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_837), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_866), .Y(n_915) );
INVxp67_ASAP7_75t_SL g916 ( .A(n_865), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_876), .B(n_747), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_879), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_865), .B(n_819), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_882), .B(n_772), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_831), .Y(n_921) );
INVx2_ASAP7_75t_L g922 ( .A(n_853), .Y(n_922) );
AND2x4_ASAP7_75t_L g923 ( .A(n_845), .B(n_733), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_884), .A2(n_766), .B1(n_765), .B2(n_780), .C(n_740), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_829), .B(n_826), .Y(n_925) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_867), .B(n_733), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_827), .B(n_803), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_842), .B(n_798), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_824), .B(n_889), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_838), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_861), .B(n_806), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_848), .B(n_743), .Y(n_932) );
AND2x2_ASAP7_75t_L g933 ( .A(n_859), .B(n_798), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_859), .B(n_691), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_832), .B(n_691), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_874), .B(n_818), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_930), .B(n_857), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_925), .B(n_868), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_900), .B(n_862), .Y(n_939) );
INVxp67_ASAP7_75t_L g940 ( .A(n_899), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_926), .A2(n_886), .B1(n_864), .B2(n_870), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_915), .B(n_848), .Y(n_942) );
INVxp67_ASAP7_75t_L g943 ( .A(n_899), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_906), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_892), .B(n_868), .Y(n_945) );
NAND2xp5_ASAP7_75t_SL g946 ( .A(n_910), .B(n_830), .Y(n_946) );
AOI21xp33_ASAP7_75t_L g947 ( .A1(n_918), .A2(n_851), .B(n_788), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_894), .A2(n_864), .B1(n_830), .B2(n_880), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_908), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_921), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_890), .B(n_858), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_929), .B(n_852), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_903), .B(n_855), .Y(n_953) );
NOR2x1p5_ASAP7_75t_L g954 ( .A(n_916), .B(n_880), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_913), .B(n_875), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_912), .Y(n_956) );
AOI22xp5_ASAP7_75t_SL g957 ( .A1(n_904), .A2(n_881), .B1(n_880), .B2(n_885), .Y(n_957) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_896), .B(n_877), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_893), .B(n_846), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_914), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_916), .Y(n_961) );
INVx2_ASAP7_75t_L g962 ( .A(n_922), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_922), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_895), .Y(n_964) );
NOR2x1_ASAP7_75t_L g965 ( .A(n_954), .B(n_885), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_964), .B(n_900), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_952), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_959), .Y(n_968) );
AOI21xp33_ASAP7_75t_L g969 ( .A1(n_958), .A2(n_920), .B(n_901), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_937), .B(n_920), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_944), .Y(n_971) );
A2O1A1Ixp33_ASAP7_75t_L g972 ( .A1(n_957), .A2(n_926), .B(n_923), .C(n_924), .Y(n_972) );
NAND2xp33_ASAP7_75t_L g973 ( .A(n_941), .B(n_894), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_950), .B(n_897), .Y(n_974) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_948), .A2(n_931), .B1(n_885), .B2(n_891), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_946), .A2(n_923), .B1(n_927), .B2(n_917), .Y(n_976) );
AND2x4_ASAP7_75t_L g977 ( .A(n_946), .B(n_938), .Y(n_977) );
OAI21xp5_ASAP7_75t_L g978 ( .A1(n_940), .A2(n_770), .B(n_877), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_961), .B(n_935), .Y(n_979) );
AOI221xp5_ASAP7_75t_L g980 ( .A1(n_947), .A2(n_898), .B1(n_905), .B2(n_909), .C(n_932), .Y(n_980) );
O2A1O1Ixp5_ASAP7_75t_L g981 ( .A1(n_972), .A2(n_949), .B(n_942), .C(n_960), .Y(n_981) );
OAI22xp33_ASAP7_75t_L g982 ( .A1(n_976), .A2(n_940), .B1(n_943), .B2(n_923), .Y(n_982) );
OAI22xp33_ASAP7_75t_L g983 ( .A1(n_975), .A2(n_943), .B1(n_902), .B2(n_936), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_980), .B(n_939), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_973), .A2(n_945), .B1(n_953), .B2(n_907), .Y(n_985) );
OAI22xp33_ASAP7_75t_L g986 ( .A1(n_965), .A2(n_849), .B1(n_956), .B2(n_955), .Y(n_986) );
OAI221xp5_ASAP7_75t_L g987 ( .A1(n_969), .A2(n_939), .B1(n_849), .B2(n_951), .C(n_828), .Y(n_987) );
AO21x1_ASAP7_75t_L g988 ( .A1(n_977), .A2(n_770), .B(n_781), .Y(n_988) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_970), .A2(n_963), .B1(n_962), .B2(n_933), .C(n_928), .Y(n_989) );
OAI22xp33_ASAP7_75t_L g990 ( .A1(n_977), .A2(n_962), .B1(n_919), .B2(n_933), .Y(n_990) );
NAND3xp33_ASAP7_75t_L g991 ( .A(n_978), .B(n_828), .C(n_887), .Y(n_991) );
OAI221xp5_ASAP7_75t_L g992 ( .A1(n_967), .A2(n_928), .B1(n_873), .B2(n_911), .C(n_863), .Y(n_992) );
OAI211xp5_ASAP7_75t_L g993 ( .A1(n_968), .A2(n_779), .B(n_869), .C(n_863), .Y(n_993) );
NOR3xp33_ASAP7_75t_L g994 ( .A(n_971), .B(n_743), .C(n_740), .Y(n_994) );
AOI211xp5_ASAP7_75t_L g995 ( .A1(n_966), .A2(n_845), .B(n_913), .C(n_814), .Y(n_995) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_974), .A2(n_935), .B1(n_934), .B2(n_845), .C(n_883), .Y(n_996) );
NAND4xp75_ASAP7_75t_L g997 ( .A(n_979), .B(n_768), .C(n_763), .D(n_792), .Y(n_997) );
AOI21xp33_ASAP7_75t_L g998 ( .A1(n_981), .A2(n_988), .B(n_984), .Y(n_998) );
NOR3xp33_ASAP7_75t_L g999 ( .A(n_986), .B(n_982), .C(n_987), .Y(n_999) );
NOR2xp67_ASAP7_75t_L g1000 ( .A(n_991), .B(n_993), .Y(n_1000) );
OA211x2_ASAP7_75t_L g1001 ( .A1(n_985), .A2(n_989), .B(n_996), .C(n_983), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_999), .B(n_995), .Y(n_1002) );
NAND2x1p5_ASAP7_75t_L g1003 ( .A(n_1000), .B(n_796), .Y(n_1003) );
NAND3xp33_ASAP7_75t_L g1004 ( .A(n_998), .B(n_994), .C(n_992), .Y(n_1004) );
NOR3xp33_ASAP7_75t_L g1005 ( .A(n_1002), .B(n_1001), .C(n_997), .Y(n_1005) );
NAND4xp75_ASAP7_75t_L g1006 ( .A(n_1003), .B(n_682), .C(n_711), .D(n_758), .Y(n_1006) );
INVx2_ASAP7_75t_L g1007 ( .A(n_1006), .Y(n_1007) );
OAI221xp5_ASAP7_75t_L g1008 ( .A1(n_1005), .A2(n_1004), .B1(n_760), .B2(n_811), .C(n_863), .Y(n_1008) );
HB1xp67_ASAP7_75t_L g1009 ( .A(n_1007), .Y(n_1009) );
AOI22x1_ASAP7_75t_L g1010 ( .A1(n_1009), .A2(n_1008), .B1(n_990), .B2(n_847), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_1010), .A2(n_847), .B1(n_883), .B2(n_871), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1011), .Y(n_1012) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_1012), .B(n_878), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_1013), .A2(n_934), .B1(n_860), .B2(n_853), .Y(n_1014) );
endmodule