module fake_jpeg_17940_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_28),
.Y(n_65)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_30),
.B1(n_16),
.B2(n_27),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_53),
.B1(n_16),
.B2(n_31),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_23),
.C(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_48),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_60),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_30),
.B1(n_16),
.B2(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_57),
.Y(n_75)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_18),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_76),
.Y(n_108)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_81),
.B1(n_83),
.B2(n_85),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_86),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_27),
.B1(n_19),
.B2(n_32),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_19),
.B1(n_32),
.B2(n_16),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_19),
.B1(n_32),
.B2(n_16),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_29),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_17),
.C(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_60),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_26),
.C(n_22),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_43),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_69),
.B(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_101),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_19),
.B1(n_32),
.B2(n_24),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_96),
.A2(n_105),
.B1(n_115),
.B2(n_31),
.Y(n_140)
);

FAx1_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_77),
.CI(n_53),
.CON(n_99),
.SN(n_99)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_75),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_24),
.B1(n_32),
.B2(n_53),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_87),
.B1(n_56),
.B2(n_37),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_46),
.C(n_23),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_104),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_53),
.B1(n_56),
.B2(n_41),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_31),
.B1(n_17),
.B2(n_25),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_24),
.B1(n_37),
.B2(n_41),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_44),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_21),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_18),
.B1(n_17),
.B2(n_22),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_120),
.B(n_123),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_92),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_107),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_143),
.B(n_20),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_131),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_91),
.B1(n_78),
.B2(n_73),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_90),
.B1(n_24),
.B2(n_58),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_57),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_142),
.C(n_147),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_133),
.Y(n_158)
);

BUFx24_ASAP7_75t_SL g133 ( 
.A(n_110),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_0),
.B(n_1),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_135),
.A2(n_136),
.B(n_137),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_31),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_146),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_99),
.A2(n_25),
.B1(n_18),
.B2(n_22),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_26),
.B1(n_25),
.B2(n_20),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_111),
.B1(n_109),
.B2(n_21),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_106),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_28),
.C(n_33),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_98),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_114),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_92),
.B(n_104),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_137),
.B1(n_136),
.B2(n_120),
.Y(n_186)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_153),
.B(n_155),
.Y(n_199)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_116),
.A3(n_102),
.B1(n_118),
.B2(n_114),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_160),
.C(n_165),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_103),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_112),
.C(n_105),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_169),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_23),
.B(n_28),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_172),
.B(n_1),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_174),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_134),
.A2(n_28),
.B(n_33),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_21),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_148),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_175),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

INVxp33_ASAP7_75t_SL g187 ( 
.A(n_176),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_80),
.C(n_40),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_179),
.C(n_67),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_0),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_144),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_50),
.C(n_33),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_181),
.B(n_205),
.Y(n_208)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_136),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_194),
.C(n_197),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_186),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_126),
.B1(n_135),
.B2(n_125),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_151),
.A2(n_131),
.B1(n_139),
.B2(n_122),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_67),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_196),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_168),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_159),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_178),
.B1(n_13),
.B2(n_15),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_167),
.B(n_170),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_9),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_165),
.C(n_177),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_159),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_203),
.A2(n_206),
.B1(n_173),
.B2(n_169),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_153),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_206)
);

AOI22x1_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_149),
.B1(n_152),
.B2(n_172),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_209),
.A2(n_228),
.B1(n_233),
.B2(n_7),
.Y(n_254)
);

XOR2x2_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_152),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_SL g253 ( 
.A(n_210),
.B(n_213),
.C(n_226),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_192),
.B(n_158),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_212),
.B(n_218),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_194),
.B(n_163),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_164),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_227),
.B(n_191),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_193),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_231),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_154),
.Y(n_220)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_224),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_201),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_183),
.A2(n_175),
.B1(n_176),
.B2(n_149),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_157),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_157),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_229),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_179),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_232),
.C(n_181),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_171),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_197),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_207),
.B1(n_188),
.B2(n_199),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_235),
.A2(n_239),
.B1(n_249),
.B2(n_238),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_150),
.B1(n_161),
.B2(n_166),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_243),
.C(n_244),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_200),
.C(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_209),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_217),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_209),
.A2(n_203),
.B1(n_3),
.B2(n_5),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_2),
.C(n_5),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_252),
.C(n_227),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_6),
.C(n_7),
.Y(n_252)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_254),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_213),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_268),
.Y(n_285)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_222),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_265),
.C(n_269),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_246),
.Y(n_263)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_225),
.C(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_233),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_267),
.Y(n_281)
);

XNOR2x1_ASAP7_75t_SL g268 ( 
.A(n_254),
.B(n_210),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_228),
.C(n_208),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_235),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_245),
.A2(n_229),
.B1(n_217),
.B2(n_214),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_271),
.A2(n_261),
.B1(n_256),
.B2(n_268),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_240),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_248),
.Y(n_278)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_234),
.B(n_211),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_280),
.A2(n_10),
.B(n_11),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_252),
.C(n_247),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_10),
.C(n_11),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_249),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_265),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_259),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_285),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_254),
.B(n_269),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_288),
.A2(n_291),
.B(n_299),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_218),
.B(n_237),
.Y(n_289)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_289),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_293),
.C(n_297),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_257),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_236),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_284),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_277),
.B(n_7),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_12),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_282),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_300),
.A2(n_303),
.B(n_287),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_305),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_290),
.A2(n_272),
.B1(n_279),
.B2(n_283),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_299),
.C(n_297),
.Y(n_314)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_288),
.A2(n_274),
.B(n_275),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_306),
.B(n_309),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_278),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_286),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_312),
.B(n_315),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_314),
.B1(n_316),
.B2(n_307),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_308),
.B(n_289),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_301),
.B(n_293),
.Y(n_316)
);

AOI21xp33_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_318),
.B(n_309),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_310),
.B(n_319),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_275),
.B(n_14),
.C(n_6),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_323),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_6),
.B(n_320),
.Y(n_325)
);


endmodule