module fake_jpeg_20314_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx6p67_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_48),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_31),
.B1(n_22),
.B2(n_30),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_22),
.B1(n_31),
.B2(n_39),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_22),
.B1(n_34),
.B2(n_17),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_27),
.B1(n_47),
.B2(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_67),
.B(n_28),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_25),
.B1(n_21),
.B2(n_24),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_21),
.B1(n_24),
.B2(n_29),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_90),
.B1(n_96),
.B2(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_53),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_32),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_94),
.C(n_32),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_99),
.Y(n_104)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_81),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_27),
.B1(n_21),
.B2(n_29),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

OAI32xp33_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_58),
.A3(n_64),
.B1(n_45),
.B2(n_25),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_84),
.B(n_89),
.Y(n_115)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_65),
.B1(n_57),
.B2(n_52),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_86),
.A2(n_33),
.B1(n_26),
.B2(n_23),
.Y(n_133)
);

BUFx4f_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_87),
.Y(n_122)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_28),
.B1(n_19),
.B2(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_32),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_20),
.B1(n_28),
.B2(n_19),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_93),
.A2(n_95),
.B1(n_36),
.B2(n_33),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_57),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_65),
.A2(n_42),
.B1(n_46),
.B2(n_44),
.Y(n_96)
);

AO22x2_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_48),
.B1(n_37),
.B2(n_42),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_36),
.B1(n_33),
.B2(n_26),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_17),
.B1(n_34),
.B2(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_48),
.B(n_34),
.C(n_18),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_123),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_37),
.C(n_32),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_113),
.C(n_87),
.Y(n_145)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_37),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_111),
.B(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_48),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_70),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_121),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_33),
.B1(n_26),
.B2(n_23),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_26),
.B1(n_23),
.B2(n_36),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_32),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_126),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_69),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_97),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_129),
.A2(n_131),
.B1(n_72),
.B2(n_87),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_94),
.B(n_97),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_68),
.A2(n_18),
.B1(n_10),
.B2(n_15),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_96),
.B1(n_100),
.B2(n_99),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_139),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_140),
.B1(n_151),
.B2(n_127),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_112),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_97),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_107),
.B1(n_114),
.B2(n_125),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_148),
.B1(n_140),
.B2(n_136),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_101),
.B1(n_75),
.B2(n_76),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_156),
.B1(n_161),
.B2(n_133),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_117),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_88),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_157),
.Y(n_173)
);

INVx3_ASAP7_75t_SL g147 ( 
.A(n_118),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_85),
.B1(n_82),
.B2(n_68),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_116),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_18),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_158),
.Y(n_183)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_123),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_132),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_125),
.A2(n_23),
.B1(n_18),
.B2(n_83),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_185),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_174),
.B1(n_179),
.B2(n_191),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_103),
.C(n_105),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_167),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_175),
.C(n_186),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_111),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_150),
.B(n_111),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_168),
.B(n_171),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_142),
.B(n_155),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_169),
.A2(n_170),
.B(n_172),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_127),
.B(n_126),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_146),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_130),
.B(n_110),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_145),
.B(n_110),
.Y(n_175)
);

XOR2x1_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_126),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_176),
.A2(n_170),
.B(n_190),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_130),
.B1(n_122),
.B2(n_132),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_148),
.B1(n_151),
.B2(n_137),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_130),
.B1(n_122),
.B2(n_108),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_187),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_157),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_108),
.C(n_124),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_120),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_135),
.A2(n_120),
.B(n_109),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_147),
.B(n_1),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_135),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_190),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_124),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_137),
.A2(n_122),
.B1(n_109),
.B2(n_92),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_194),
.B(n_195),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_164),
.A2(n_143),
.B1(n_156),
.B2(n_138),
.Y(n_197)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_176),
.A3(n_184),
.B1(n_175),
.B2(n_172),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_11),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_161),
.B1(n_149),
.B2(n_153),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_208),
.B1(n_219),
.B2(n_223),
.Y(n_236)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_178),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_205),
.B(n_218),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_154),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_149),
.B1(n_152),
.B2(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_180),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_215),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_212),
.A2(n_213),
.B(n_217),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_168),
.A2(n_177),
.B(n_188),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_147),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_222),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_186),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_166),
.A2(n_92),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_92),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_167),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_181),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_0),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_220),
.Y(n_227)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_165),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_232),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_183),
.C(n_14),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_240),
.C(n_241),
.Y(n_252)
);

AOI21xp33_ASAP7_75t_L g233 ( 
.A1(n_193),
.A2(n_10),
.B(n_1),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_217),
.B1(n_211),
.B2(n_210),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_203),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_224),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_10),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_0),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_0),
.C(n_2),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_249),
.C(n_248),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_245),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_207),
.A2(n_0),
.B(n_2),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_3),
.B(n_4),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_198),
.B(n_2),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_207),
.A2(n_212),
.B(n_213),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g253 ( 
.A1(n_246),
.A2(n_218),
.B1(n_244),
.B2(n_225),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_267),
.B1(n_236),
.B2(n_219),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_256),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_195),
.B1(n_197),
.B2(n_199),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_258),
.B1(n_264),
.B2(n_265),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_202),
.Y(n_259)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_259),
.Y(n_287)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_262),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_204),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_239),
.B(n_223),
.Y(n_264)
);

BUFx12_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_243),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_270),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_242),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_268),
.A2(n_247),
.B1(n_242),
.B2(n_222),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_236),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_235),
.A2(n_199),
.B(n_194),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_250),
.B(n_246),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_284),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_228),
.C(n_231),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_276),
.C(n_282),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_249),
.C(n_257),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_235),
.B(n_230),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_265),
.B(n_232),
.CI(n_241),
.CON(n_279),
.SN(n_279)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_230),
.B(n_208),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_214),
.C(n_201),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_240),
.C(n_210),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_289),
.C(n_256),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_288),
.B1(n_290),
.B2(n_251),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_253),
.A2(n_204),
.B1(n_247),
.B2(n_200),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_209),
.C(n_234),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_234),
.B1(n_5),
.B2(n_6),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_254),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_291),
.B(n_294),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_277),
.B(n_260),
.Y(n_295)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_261),
.C(n_255),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_297),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_262),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_272),
.B1(n_286),
.B2(n_287),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_265),
.Y(n_300)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_273),
.A2(n_251),
.B1(n_268),
.B2(n_260),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_288),
.B1(n_272),
.B2(n_279),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_304),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_258),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_274),
.B(n_3),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_280),
.C(n_290),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_315),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_284),
.C(n_281),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_305),
.C(n_292),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_317),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_300),
.A2(n_272),
.B1(n_278),
.B2(n_279),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_298),
.A2(n_301),
.B(n_293),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_301),
.B(n_306),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_298),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_9),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_323),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_318),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_325),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_292),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_323),
.B(n_324),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_303),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_316),
.B(n_3),
.CI(n_5),
.CON(n_327),
.SN(n_327)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_321),
.A2(n_312),
.B(n_308),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_332),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_309),
.C(n_314),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_313),
.C(n_311),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_334),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_329),
.A2(n_319),
.B(n_325),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_336),
.B(n_334),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_337),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_335),
.C(n_333),
.Y(n_340)
);

AOI322xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_330),
.A3(n_328),
.B1(n_327),
.B2(n_307),
.C1(n_9),
.C2(n_8),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_341),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_7),
.B(n_8),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_7),
.C(n_8),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_7),
.C(n_9),
.Y(n_345)
);


endmodule