module fake_netlist_1_484_n_40 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_30;
wire n_25;
wire n_26;
wire n_13;
wire n_16;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
wire n_39;
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_4), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_1), .B(n_10), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_6), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_8), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_5), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_12), .B(n_0), .Y(n_19) );
A2O1A1Ixp33_ASAP7_75t_L g20 ( .A1(n_12), .A2(n_1), .B(n_2), .C(n_3), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_12), .Y(n_21) );
NOR2xp33_ASAP7_75t_SL g22 ( .A(n_17), .B(n_3), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_18), .Y(n_23) );
NOR2xp67_ASAP7_75t_L g24 ( .A(n_17), .B(n_4), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_21), .Y(n_25) );
OAI22xp33_ASAP7_75t_L g26 ( .A1(n_22), .A2(n_18), .B1(n_14), .B2(n_11), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_21), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_23), .B(n_14), .Y(n_28) );
AOI22xp33_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_19), .B1(n_24), .B2(n_23), .Y(n_29) );
AOI22xp33_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_24), .B1(n_13), .B2(n_15), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_29), .B(n_26), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_25), .Y(n_32) );
OAI32xp33_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_25), .A3(n_27), .B1(n_16), .B2(n_13), .Y(n_33) );
NOR2xp33_ASAP7_75t_L g34 ( .A(n_32), .B(n_20), .Y(n_34) );
NOR2xp33_ASAP7_75t_R g35 ( .A(n_34), .B(n_32), .Y(n_35) );
OAI221xp5_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_27), .B1(n_6), .B2(n_7), .C(n_9), .Y(n_36) );
INVx1_ASAP7_75t_SL g37 ( .A(n_35), .Y(n_37) );
CKINVDCx12_ASAP7_75t_R g38 ( .A(n_36), .Y(n_38) );
NOR3xp33_ASAP7_75t_SL g39 ( .A(n_37), .B(n_38), .C(n_7), .Y(n_39) );
AOI22xp33_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_37), .B1(n_5), .B2(n_9), .Y(n_40) );
endmodule