module fake_jpeg_19872_n_183 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_9),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g31 ( 
.A(n_20),
.B(n_6),
.CON(n_31),
.SN(n_31)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_32),
.B1(n_18),
.B2(n_22),
.Y(n_44)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_36),
.B1(n_39),
.B2(n_14),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_15),
.B1(n_17),
.B2(n_23),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_21),
.B1(n_20),
.B2(n_23),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_23),
.B1(n_21),
.B2(n_13),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_32),
.B1(n_30),
.B2(n_26),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_12),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_14),
.B(n_22),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_29),
.B(n_26),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_54),
.B(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_32),
.B1(n_30),
.B2(n_22),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_56),
.B1(n_58),
.B2(n_40),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_60),
.Y(n_78)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_24),
.B1(n_22),
.B2(n_14),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_24),
.B1(n_12),
.B2(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_66),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_41),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_40),
.B1(n_38),
.B2(n_34),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_68),
.B1(n_74),
.B2(n_35),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_44),
.C(n_36),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_72),
.C(n_60),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_73),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_44),
.C(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_34),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_44),
.B1(n_35),
.B2(n_37),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_82),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_53),
.B1(n_60),
.B2(n_35),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_79),
.B1(n_71),
.B2(n_24),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_60),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_47),
.B(n_50),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_84),
.B(n_88),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_37),
.B(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_89),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_59),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_90),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_69),
.B(n_72),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_67),
.B1(n_68),
.B2(n_74),
.Y(n_89)
);

A2O1A1O1Ixp25_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_63),
.B(n_62),
.C(n_77),
.D(n_75),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_35),
.B1(n_37),
.B2(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_96),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_47),
.B(n_1),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_93),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_43),
.B1(n_55),
.B2(n_24),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_55),
.C(n_43),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_43),
.C(n_57),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_108),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_91),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_100),
.B(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_8),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_64),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_112),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_87),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_SL g118 ( 
.A1(n_114),
.A2(n_87),
.A3(n_89),
.B1(n_92),
.B2(n_94),
.C1(n_82),
.C2(n_83),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_71),
.C(n_64),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_11),
.C(n_9),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_130),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_92),
.B(n_84),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_102),
.B(n_128),
.Y(n_142)
);

OAI322xp33_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_94),
.A3(n_92),
.B1(n_85),
.B2(n_8),
.C1(n_10),
.C2(n_11),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_124),
.B(n_7),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_106),
.C(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_128),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_0),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_9),
.B1(n_8),
.B2(n_7),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_106),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_141),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_101),
.B(n_103),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_137),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_115),
.C(n_108),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_121),
.C(n_129),
.Y(n_144)
);

AOI31xp67_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_119),
.A3(n_131),
.B(n_3),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_110),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_107),
.B(n_126),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_151),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_143),
.A2(n_134),
.B1(n_130),
.B2(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_120),
.B1(n_133),
.B2(n_121),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_152),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_150),
.A2(n_136),
.B(n_107),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_125),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_127),
.C(n_120),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_153),
.A2(n_139),
.B(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_144),
.B(n_119),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_155),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_151),
.B(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_149),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_141),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_1),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_142),
.B(n_137),
.C(n_4),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_162),
.A2(n_148),
.B1(n_2),
.B2(n_4),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_154),
.C(n_152),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_158),
.C(n_168),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_169),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_168),
.Y(n_173)
);

NOR2x1_ASAP7_75t_R g169 ( 
.A(n_162),
.B(n_4),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_164),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_156),
.B(n_169),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_5),
.B(n_171),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_176),
.B(n_177),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_157),
.B(n_159),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_165),
.B(n_161),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_5),
.B(n_172),
.C(n_169),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_180),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_5),
.Y(n_183)
);


endmodule