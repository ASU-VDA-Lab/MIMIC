module fake_jpeg_22595_n_37 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_37);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_24),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_0),
.C(n_1),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_9),
.B(n_10),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_19),
.B1(n_18),
.B2(n_0),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_27),
.B(n_28),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_11),
.B(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_33),
.Y(n_35)
);

OAI22x1_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_31),
.B1(n_30),
.B2(n_16),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_14),
.B(n_15),
.Y(n_37)
);


endmodule