module fake_jpeg_30114_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_20),
.A2(n_0),
.B(n_1),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_33),
.C(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_45),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_35),
.B1(n_36),
.B2(n_32),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_53),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_116)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_22),
.B1(n_19),
.B2(n_28),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_64),
.B1(n_33),
.B2(n_28),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_17),
.Y(n_78)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_33),
.B1(n_22),
.B2(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_29),
.Y(n_81)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_31),
.Y(n_108)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_81),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_33),
.B1(n_30),
.B2(n_22),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_76),
.A2(n_93),
.B1(n_113),
.B2(n_21),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_77),
.A2(n_88),
.B1(n_89),
.B2(n_100),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_92),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_82),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx8_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_25),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_95),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_38),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_90),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_41),
.B1(n_40),
.B2(n_34),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_41),
.B1(n_40),
.B2(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_24),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_39),
.A3(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_47),
.C(n_44),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_30),
.B1(n_31),
.B2(n_20),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_96),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_31),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_103),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_31),
.B1(n_36),
.B2(n_20),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_112),
.B1(n_39),
.B2(n_26),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_20),
.B1(n_47),
.B2(n_30),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_56),
.B(n_11),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_54),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_105),
.B(n_110),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_58),
.Y(n_107)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_26),
.CI(n_21),
.CON(n_140),
.SN(n_140)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_111),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_31),
.B1(n_39),
.B2(n_26),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_54),
.A2(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_115),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_18),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_73),
.B1(n_39),
.B2(n_11),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_135),
.B1(n_98),
.B2(n_90),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_135),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_73),
.B1(n_10),
.B2(n_12),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_78),
.B(n_79),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_136),
.B(n_104),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_92),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_142),
.B1(n_107),
.B2(n_110),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_82),
.A2(n_0),
.B(n_1),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_147),
.B(n_105),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_1),
.B(n_2),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_91),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_87),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_149),
.A2(n_152),
.B1(n_165),
.B2(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_139),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_151),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_154),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_104),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_157),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_109),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_156),
.C(n_159),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_109),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_134),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_94),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_167),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_94),
.B(n_83),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_164),
.Y(n_192)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_107),
.B1(n_111),
.B2(n_86),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_168),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_101),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_172),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_118),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_170),
.Y(n_191)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_173),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_167),
.B1(n_170),
.B2(n_168),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_125),
.A2(n_84),
.B1(n_106),
.B2(n_115),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_176),
.A2(n_179),
.B1(n_123),
.B2(n_143),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_96),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_177),
.A2(n_121),
.B(n_75),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_136),
.B(n_16),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_178),
.A2(n_141),
.B(n_147),
.Y(n_183)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_150),
.A2(n_152),
.B1(n_163),
.B2(n_175),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_180),
.A2(n_181),
.B(n_207),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_145),
.B(n_124),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_182),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_174),
.A2(n_127),
.B1(n_124),
.B2(n_130),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_184),
.A2(n_200),
.B1(n_202),
.B2(n_198),
.Y(n_227)
);

INVx3_ASAP7_75t_SL g240 ( 
.A(n_185),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_199),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_124),
.C(n_140),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_188),
.C(n_206),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_140),
.C(n_134),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_146),
.B(n_128),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_197),
.A2(n_198),
.B(n_204),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_151),
.A2(n_146),
.B(n_128),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_151),
.A2(n_153),
.B1(n_154),
.B2(n_161),
.Y(n_200)
);

AND2x4_ASAP7_75t_SL g203 ( 
.A(n_165),
.B(n_123),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_122),
.B(n_137),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_155),
.B(n_126),
.C(n_131),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_164),
.A2(n_80),
.B(n_118),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_121),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_212),
.B(n_126),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_213),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_180),
.A2(n_211),
.B1(n_208),
.B2(n_181),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_219),
.B1(n_233),
.B2(n_202),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_178),
.Y(n_216)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_172),
.Y(n_217)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_143),
.B1(n_173),
.B2(n_169),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_206),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_171),
.Y(n_221)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_176),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_223),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_176),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_190),
.B(n_188),
.Y(n_248)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_229),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_234),
.B1(n_235),
.B2(n_185),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_190),
.B(n_197),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_228),
.A2(n_232),
.B(n_226),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_102),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_201),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_236),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_193),
.A2(n_114),
.B1(n_85),
.B2(n_75),
.Y(n_233)
);

OAI22x1_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_97),
.B1(n_114),
.B2(n_85),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_182),
.A2(n_21),
.B1(n_18),
.B2(n_97),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_201),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_200),
.B(n_14),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_238),
.B(n_239),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_194),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_196),
.B(n_18),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_222),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_205),
.C(n_186),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_252),
.C(n_265),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_227),
.B1(n_226),
.B2(n_213),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_246),
.A2(n_231),
.B1(n_225),
.B2(n_230),
.Y(n_282)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_199),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_251),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_196),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_216),
.A2(n_183),
.B1(n_203),
.B2(n_210),
.Y(n_253)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_203),
.B1(n_210),
.B2(n_184),
.Y(n_254)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_261),
.B(n_228),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_219),
.A2(n_209),
.B1(n_207),
.B2(n_204),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_260),
.A2(n_262),
.B1(n_240),
.B2(n_234),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_232),
.A2(n_212),
.B(n_195),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_214),
.A2(n_195),
.B1(n_12),
.B2(n_10),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_215),
.B(n_12),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_242),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_273),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_268),
.A2(n_276),
.B1(n_250),
.B2(n_264),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_215),
.C(n_238),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_279),
.C(n_284),
.Y(n_288)
);

HAxp5_ASAP7_75t_SL g301 ( 
.A(n_270),
.B(n_277),
.CON(n_301),
.SN(n_301)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_240),
.B(n_234),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_261),
.B(n_247),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_218),
.Y(n_273)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_240),
.B1(n_231),
.B2(n_236),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_282),
.B1(n_260),
.B2(n_245),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_243),
.B(n_223),
.Y(n_278)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_249),
.C(n_251),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_221),
.C(n_239),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_229),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_285),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_10),
.C(n_3),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_262),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_295),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_303),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_292),
.A2(n_301),
.B(n_302),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_263),
.B(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

NAND3xp33_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_263),
.C(n_255),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_294),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_250),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_3),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_298),
.A2(n_267),
.B1(n_5),
.B2(n_6),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_270),
.A2(n_281),
.B(n_282),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_2),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_269),
.C(n_279),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_304),
.B(n_311),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_298),
.A2(n_283),
.B1(n_271),
.B2(n_284),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_305),
.A2(n_312),
.B1(n_299),
.B2(n_301),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_276),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_308),
.Y(n_325)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_267),
.C(n_286),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_303),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_302),
.A2(n_3),
.B(n_5),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_292),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_310),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_321),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_327),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_297),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_323),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_291),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_326),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_289),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_307),
.B(n_295),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_313),
.B(n_309),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_328),
.A2(n_331),
.B(n_329),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_310),
.C(n_306),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_333),
.B(n_5),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_325),
.A2(n_313),
.B1(n_287),
.B2(n_315),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_325),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_336),
.C(n_337),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_332),
.A2(n_312),
.B1(n_314),
.B2(n_6),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_333),
.B(n_3),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_338),
.A2(n_339),
.B(n_330),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_340),
.B(n_334),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_341),
.B1(n_7),
.B2(n_8),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_343),
.A2(n_6),
.B(n_8),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_344),
.B(n_6),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_345),
.B(n_8),
.Y(n_346)
);


endmodule