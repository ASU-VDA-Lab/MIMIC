module fake_netlist_6_4357_n_2104 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2104);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2104;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_1159;
wire n_276;
wire n_995;
wire n_1092;
wire n_441;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_204),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_94),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_7),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_160),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_6),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_32),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_92),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_159),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_93),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_178),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_112),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_172),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_91),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_19),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_88),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_188),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_78),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_183),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_138),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_30),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_76),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_130),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_104),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_182),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_146),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_120),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_127),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_71),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_132),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_124),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_37),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_47),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_213),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_193),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_33),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_97),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_166),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_200),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_176),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_75),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_203),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_134),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_149),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_46),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_129),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_45),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_66),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_44),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_89),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_148),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_71),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_185),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_51),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_126),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_4),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_131),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_225),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_133),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_31),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_29),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_95),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_59),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_210),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_43),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_150),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_143),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_48),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_44),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_70),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_26),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_61),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_28),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_197),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_18),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_51),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_68),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_47),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_54),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_184),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_84),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_86),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_27),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_62),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_177),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_109),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_27),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_144),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_26),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_29),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_206),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_69),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_52),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_212),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_152),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_96),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_57),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_42),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_145),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_10),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_8),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_70),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_77),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_116),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_87),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_113),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_19),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_192),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_99),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_155),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_174),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_226),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_50),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_190),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_3),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_34),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_208),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_223),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_168),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_179),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_8),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_157),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_82),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_170),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_106),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_189),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_58),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_202),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_50),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_158),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_169),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_135),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_220),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_103),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_224),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_137),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_20),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_52),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_198),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_147),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_14),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_123),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_222),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_211),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_69),
.Y(n_377)
);

INVxp33_ASAP7_75t_SL g378 ( 
.A(n_45),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_101),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_171),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_139),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_54),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_22),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_201),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_167),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_196),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_80),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_136),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_63),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_161),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_153),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_2),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_49),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_180),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_23),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g396 ( 
.A(n_67),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_68),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_61),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_32),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_56),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_18),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_12),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_194),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_214),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_40),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_108),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_42),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_62),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_64),
.Y(n_409)
);

INVxp33_ASAP7_75t_R g410 ( 
.A(n_43),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_5),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_156),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_53),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_12),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_66),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_207),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_67),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_209),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_35),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_215),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_40),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_175),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_16),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_118),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_39),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_151),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_49),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_125),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_64),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_14),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_3),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_38),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_9),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_114),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_142),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_205),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_15),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_55),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_20),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_164),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_117),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_0),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_140),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_163),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_2),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_57),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_15),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_243),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_304),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_248),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_275),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_301),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_282),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_383),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_396),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_251),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_301),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_265),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_397),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_312),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_336),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_264),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_280),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_264),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_264),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_264),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_336),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_349),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_264),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_435),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_445),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_445),
.Y(n_473)
);

INVxp33_ASAP7_75t_L g474 ( 
.A(n_233),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_301),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_340),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_445),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_286),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_445),
.Y(n_479)
);

INVxp33_ASAP7_75t_L g480 ( 
.A(n_277),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_445),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_288),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_319),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_292),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_319),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_324),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_324),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_297),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_242),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_300),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_231),
.Y(n_491)
);

INVxp33_ASAP7_75t_SL g492 ( 
.A(n_231),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_281),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_284),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_293),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_379),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_295),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_303),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_305),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_259),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_307),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_379),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_316),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_321),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_329),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_302),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_234),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_333),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_334),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_310),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_322),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_325),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_285),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_345),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_361),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_330),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_228),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_271),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_372),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_237),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_370),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_234),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_244),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_400),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_401),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_332),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_347),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_240),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_239),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_402),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_408),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_272),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_240),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_417),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_353),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_359),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_334),
.Y(n_537)
);

INVxp67_ASAP7_75t_SL g538 ( 
.A(n_245),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_273),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_421),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_377),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_423),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_438),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_240),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_439),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_447),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_247),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_253),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_254),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_255),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_369),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_256),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_257),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_260),
.Y(n_554)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_262),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_373),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_377),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_419),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_382),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_419),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_429),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_263),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_244),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_262),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_276),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_269),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g567 ( 
.A(n_262),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_270),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_261),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_513),
.B(n_320),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_467),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_462),
.B(n_371),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_450),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_467),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_457),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_465),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_520),
.B(n_371),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_517),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_468),
.B(n_429),
.Y(n_579)
);

OA21x2_ASAP7_75t_L g580 ( 
.A1(n_465),
.A2(n_422),
.B(n_229),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_533),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_452),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_467),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_466),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_466),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_470),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_454),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_528),
.A2(n_309),
.B1(n_315),
.B2(n_308),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_496),
.B(n_229),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_470),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_529),
.B(n_422),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_472),
.Y(n_592)
);

BUFx8_ASAP7_75t_L g593 ( 
.A(n_522),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_472),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_473),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_473),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_477),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_518),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_457),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_461),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_538),
.B(n_436),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_477),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_448),
.A2(n_279),
.B1(n_405),
.B2(n_261),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_479),
.Y(n_604)
);

BUFx8_ASAP7_75t_L g605 ( 
.A(n_522),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_479),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_456),
.B(n_246),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_532),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_469),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_463),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_502),
.B(n_436),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_471),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_491),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_539),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_460),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_481),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_481),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_565),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_483),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_460),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_451),
.B(n_430),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_458),
.B(n_453),
.Y(n_622)
);

AND2x6_ASAP7_75t_L g623 ( 
.A(n_513),
.B(n_320),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_483),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_485),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_533),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_485),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_547),
.B(n_548),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_486),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_486),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_544),
.A2(n_555),
.B1(n_567),
.B2(n_564),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_487),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_487),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_509),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_509),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_537),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_455),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_464),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_489),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_537),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_549),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_541),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_541),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_557),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_L g645 ( 
.A(n_456),
.B(n_268),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_557),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_558),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_550),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_519),
.B(n_318),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_552),
.B(n_446),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_459),
.B(n_380),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_553),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_464),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_560),
.Y(n_654)
);

BUFx8_ASAP7_75t_L g655 ( 
.A(n_458),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_560),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_478),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_554),
.B(n_274),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_561),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_562),
.B(n_430),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_561),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_478),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_500),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_649),
.B(n_482),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_607),
.B(n_482),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_577),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_577),
.A2(n_568),
.B1(n_566),
.B2(n_446),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_641),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_592),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_585),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_585),
.Y(n_671)
);

INVxp33_ASAP7_75t_SL g672 ( 
.A(n_588),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_R g673 ( 
.A(n_653),
.B(n_484),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_577),
.B(n_484),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_585),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_591),
.A2(n_449),
.B1(n_492),
.B2(n_378),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_581),
.B(n_492),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_581),
.B(n_488),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_592),
.Y(n_679)
);

OR2x6_ASAP7_75t_L g680 ( 
.A(n_622),
.B(n_530),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_576),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_585),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_637),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_648),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_652),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_579),
.B(n_320),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_573),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_585),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_576),
.Y(n_689)
);

AO21x2_ASAP7_75t_L g690 ( 
.A1(n_589),
.A2(n_290),
.B(n_278),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_596),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_616),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_613),
.A2(n_476),
.B1(n_490),
.B2(n_488),
.Y(n_693)
);

INVxp33_ASAP7_75t_L g694 ( 
.A(n_579),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_586),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_626),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_639),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_655),
.B(n_490),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_571),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_637),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_586),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_591),
.A2(n_378),
.B1(n_523),
.B2(n_507),
.Y(n_702)
);

BUFx10_ASAP7_75t_L g703 ( 
.A(n_599),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_610),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_626),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_572),
.B(n_569),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_628),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_591),
.B(n_563),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_571),
.Y(n_709)
);

AO21x2_ASAP7_75t_L g710 ( 
.A1(n_611),
.A2(n_314),
.B(n_296),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_596),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_596),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_645),
.B(n_510),
.C(n_506),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_596),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_626),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_628),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_651),
.A2(n_506),
.B1(n_511),
.B2(n_510),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_628),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_622),
.A2(n_511),
.B1(n_516),
.B2(n_512),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_596),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_604),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_604),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_574),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_594),
.Y(n_724)
);

INVx5_ASAP7_75t_L g725 ( 
.A(n_570),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_622),
.A2(n_512),
.B1(n_526),
.B2(n_516),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_574),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_622),
.B(n_545),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_638),
.A2(n_526),
.B1(n_535),
.B2(n_527),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_583),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_583),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_584),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_658),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_655),
.B(n_527),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_575),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_594),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_655),
.B(n_535),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_604),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_584),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_601),
.B(n_536),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_601),
.B(n_493),
.Y(n_741)
);

CKINVDCx6p67_ASAP7_75t_R g742 ( 
.A(n_582),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_604),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_595),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_626),
.B(n_536),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_597),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_597),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_620),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_626),
.B(n_551),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_601),
.A2(n_495),
.B1(n_497),
.B2(n_494),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_658),
.A2(n_499),
.B1(n_501),
.B2(n_498),
.Y(n_751)
);

OR2x6_ASAP7_75t_L g752 ( 
.A(n_653),
.B(n_503),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_626),
.B(n_551),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_602),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_584),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_658),
.B(n_556),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_657),
.A2(n_556),
.B1(n_559),
.B2(n_475),
.Y(n_757)
);

BUFx10_ASAP7_75t_L g758 ( 
.A(n_639),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_590),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_602),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_650),
.A2(n_505),
.B1(n_508),
.B2(n_504),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_604),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_603),
.B(n_559),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_606),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_663),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_606),
.B(n_338),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_590),
.Y(n_767)
);

INVx4_ASAP7_75t_L g768 ( 
.A(n_570),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_662),
.B(n_474),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_590),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_617),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_617),
.B(n_418),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_650),
.Y(n_773)
);

INVx4_ASAP7_75t_L g774 ( 
.A(n_570),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_570),
.B(n_320),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_580),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_627),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_627),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_662),
.B(n_575),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_627),
.B(n_283),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_627),
.B(n_287),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_660),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_627),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_633),
.Y(n_784)
);

BUFx10_ASAP7_75t_L g785 ( 
.A(n_663),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_578),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_633),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_633),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_SL g789 ( 
.A1(n_593),
.A2(n_348),
.B1(n_389),
.B2(n_395),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_615),
.B(n_380),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_633),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_633),
.Y(n_792)
);

AND3x1_ASAP7_75t_L g793 ( 
.A(n_621),
.B(n_410),
.C(n_514),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_640),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_640),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_640),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_640),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_615),
.B(n_631),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_640),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_619),
.B(n_480),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_644),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_660),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_644),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_644),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_593),
.B(n_230),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_644),
.B(n_647),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_621),
.A2(n_580),
.B1(n_647),
.B2(n_644),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_619),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_570),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_L g810 ( 
.A(n_578),
.B(n_311),
.C(n_392),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_624),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_624),
.A2(n_399),
.B1(n_398),
.B2(n_393),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_647),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_632),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_647),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_570),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_647),
.B(n_289),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_593),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_656),
.B(n_291),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_769),
.B(n_598),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_773),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_694),
.B(n_230),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_800),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_773),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_733),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_668),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_684),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_685),
.Y(n_828)
);

BUFx6f_ASAP7_75t_SL g829 ( 
.A(n_758),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_666),
.B(n_320),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_707),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_690),
.A2(n_580),
.B1(n_431),
.B2(n_425),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_666),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_694),
.B(n_232),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_733),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_677),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_690),
.A2(n_580),
.B1(n_343),
.B2(n_331),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_776),
.B(n_656),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_752),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_674),
.B(n_740),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_687),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_776),
.B(n_331),
.Y(n_842)
);

AND2x6_ASAP7_75t_SL g843 ( 
.A(n_752),
.B(n_515),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_708),
.B(n_598),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_706),
.B(n_232),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_782),
.A2(n_802),
.B(n_756),
.C(n_741),
.Y(n_846)
);

BUFx8_ASAP7_75t_L g847 ( 
.A(n_818),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_776),
.B(n_807),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_776),
.B(n_768),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_716),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_708),
.B(n_605),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_699),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_690),
.A2(n_343),
.B1(n_331),
.B2(n_285),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_706),
.B(n_235),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_664),
.B(n_235),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_718),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_808),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_699),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_687),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_776),
.B(n_656),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_710),
.A2(n_686),
.B1(n_741),
.B2(n_689),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_772),
.B(n_656),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_811),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_709),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_717),
.B(n_665),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_709),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_814),
.B(n_661),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_757),
.B(n_605),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_723),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_724),
.B(n_744),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_683),
.B(n_605),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_746),
.B(n_661),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_683),
.B(n_236),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_747),
.B(n_661),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_700),
.B(n_236),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_723),
.Y(n_876)
);

NOR2x1p5_ASAP7_75t_L g877 ( 
.A(n_713),
.B(n_608),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_681),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_673),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_700),
.B(n_238),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_754),
.B(n_661),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_719),
.B(n_238),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_763),
.B(n_241),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_742),
.Y(n_884)
);

AOI221xp5_ASAP7_75t_L g885 ( 
.A1(n_676),
.A2(n_339),
.B1(n_268),
.B2(n_405),
.C(n_407),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_760),
.B(n_341),
.Y(n_886)
);

AO221x1_ASAP7_75t_L g887 ( 
.A1(n_812),
.A2(n_331),
.B1(n_343),
.B2(n_434),
.C(n_428),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_681),
.B(n_342),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_726),
.B(n_249),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_752),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_752),
.Y(n_891)
);

BUFx6f_ASAP7_75t_SL g892 ( 
.A(n_758),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_748),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_689),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_695),
.B(n_350),
.Y(n_895)
);

INVxp33_ASAP7_75t_L g896 ( 
.A(n_693),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_695),
.Y(n_897)
);

AO22x2_ASAP7_75t_L g898 ( 
.A1(n_798),
.A2(n_790),
.B1(n_779),
.B2(n_735),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_671),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_701),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_701),
.B(n_351),
.Y(n_901)
);

NAND2xp33_ASAP7_75t_L g902 ( 
.A(n_686),
.B(n_753),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_736),
.B(n_352),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_678),
.B(n_250),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_736),
.B(n_358),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_764),
.B(n_704),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_702),
.B(n_608),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_771),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_727),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_771),
.B(n_360),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_671),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_766),
.B(n_686),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_732),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_730),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_732),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_729),
.B(n_250),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_686),
.B(n_362),
.Y(n_917)
);

BUFx4_ASAP7_75t_L g918 ( 
.A(n_742),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_793),
.B(n_521),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_686),
.B(n_368),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_739),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_739),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_667),
.B(n_252),
.Y(n_923)
);

NAND2x1p5_ASAP7_75t_L g924 ( 
.A(n_768),
.B(n_774),
.Y(n_924)
);

AND2x6_ASAP7_75t_SL g925 ( 
.A(n_680),
.B(n_524),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_SL g926 ( 
.A(n_818),
.B(n_614),
.Y(n_926)
);

BUFx5_ASAP7_75t_L g927 ( 
.A(n_777),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_SL g928 ( 
.A(n_697),
.B(n_614),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_680),
.B(n_252),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_680),
.B(n_258),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_731),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_810),
.B(n_258),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_750),
.B(n_266),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_731),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_745),
.B(n_749),
.Y(n_935)
);

OR2x6_ASAP7_75t_SL g936 ( 
.A(n_697),
.B(n_618),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_686),
.B(n_570),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_755),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_780),
.B(n_623),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_728),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_755),
.A2(n_659),
.B(n_654),
.C(n_635),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_728),
.B(n_266),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_R g943 ( 
.A(n_765),
.B(n_618),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_759),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_768),
.B(n_331),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_710),
.A2(n_323),
.B1(n_294),
.B2(n_298),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_781),
.B(n_623),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_817),
.B(n_623),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_819),
.B(n_623),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_767),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_767),
.Y(n_951)
);

OAI22x1_ASAP7_75t_R g952 ( 
.A1(n_765),
.A2(n_587),
.B1(n_612),
.B2(n_609),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_703),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_770),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_728),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_770),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_775),
.A2(n_525),
.B(n_531),
.C(n_534),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_710),
.A2(n_343),
.B1(n_285),
.B2(n_623),
.Y(n_958)
);

OAI22xp33_ASAP7_75t_L g959 ( 
.A1(n_728),
.A2(n_414),
.B1(n_433),
.B2(n_339),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_698),
.B(n_267),
.Y(n_960)
);

INVxp33_ASAP7_75t_L g961 ( 
.A(n_789),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_788),
.B(n_623),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_788),
.B(n_623),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_788),
.B(n_625),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_791),
.B(n_625),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_816),
.B(n_404),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_669),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_L g968 ( 
.A(n_725),
.B(n_285),
.Y(n_968)
);

NOR3xp33_ASAP7_75t_L g969 ( 
.A(n_734),
.B(n_542),
.C(n_540),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_669),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_791),
.B(n_629),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_791),
.B(n_629),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_679),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_679),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_777),
.B(n_630),
.Y(n_975)
);

BUFx5_ASAP7_75t_L g976 ( 
.A(n_778),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_774),
.B(n_343),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_671),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_692),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_778),
.B(n_630),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_844),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_908),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_845),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_848),
.A2(n_860),
.B(n_838),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_831),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_850),
.Y(n_986)
);

INVx5_ASAP7_75t_L g987 ( 
.A(n_899),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_840),
.B(n_783),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_SL g989 ( 
.A1(n_961),
.A2(n_672),
.B1(n_600),
.B2(n_442),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_856),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_913),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_943),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_840),
.B(n_783),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_821),
.B(n_737),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_915),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_921),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_848),
.B(n_787),
.Y(n_997)
);

CKINVDCx6p67_ASAP7_75t_R g998 ( 
.A(n_829),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_823),
.B(n_703),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_878),
.B(n_787),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_894),
.B(n_792),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_865),
.A2(n_672),
.B1(n_797),
.B2(n_801),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_835),
.B(n_703),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_835),
.B(n_786),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_922),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_893),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_835),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_824),
.B(n_805),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_938),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_897),
.B(n_792),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_891),
.Y(n_1011)
);

NAND2xp33_ASAP7_75t_L g1012 ( 
.A(n_835),
.B(n_924),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_950),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_944),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_891),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_836),
.B(n_786),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_SL g1017 ( 
.A(n_928),
.B(n_758),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_899),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_951),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_899),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_854),
.B(n_785),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_954),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_833),
.B(n_751),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_854),
.B(n_785),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_879),
.B(n_785),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_956),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_859),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_919),
.Y(n_1028)
);

INVxp67_ASAP7_75t_SL g1029 ( 
.A(n_825),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_900),
.B(n_795),
.Y(n_1030)
);

AND2x6_ASAP7_75t_L g1031 ( 
.A(n_825),
.B(n_784),
.Y(n_1031)
);

BUFx8_ASAP7_75t_L g1032 ( 
.A(n_829),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_919),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_857),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_852),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_832),
.B(n_795),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_858),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_863),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_855),
.A2(n_797),
.B1(n_801),
.B2(n_813),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_896),
.B(n_670),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_943),
.Y(n_1041)
);

NOR2x1_ASAP7_75t_R g1042 ( 
.A(n_884),
.B(n_407),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_899),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_855),
.A2(n_794),
.B1(n_815),
.B2(n_813),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_822),
.B(n_816),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_967),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_820),
.B(n_761),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_832),
.B(n_692),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_887),
.A2(n_815),
.B1(n_794),
.B2(n_784),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_892),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_906),
.B(n_796),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_970),
.Y(n_1052)
);

O2A1O1Ixp5_ASAP7_75t_L g1053 ( 
.A1(n_945),
.A2(n_796),
.B(n_804),
.C(n_803),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_SL g1054 ( 
.A1(n_916),
.A2(n_414),
.B1(n_409),
.B2(n_411),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_973),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_864),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_940),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_861),
.B(n_799),
.Y(n_1058)
);

OA22x2_ASAP7_75t_L g1059 ( 
.A1(n_890),
.A2(n_413),
.B1(n_415),
.B2(n_427),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_866),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_847),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_822),
.B(n_834),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_842),
.A2(n_806),
.B(n_809),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_869),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_974),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_916),
.B(n_670),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_861),
.B(n_799),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_841),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_870),
.B(n_803),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_953),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_876),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_834),
.B(n_809),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_904),
.B(n_846),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_904),
.B(n_809),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_935),
.A2(n_804),
.B1(n_675),
.B2(n_738),
.Y(n_1075)
);

INVx5_ASAP7_75t_L g1076 ( 
.A(n_911),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_918),
.Y(n_1077)
);

INVx5_ASAP7_75t_L g1078 ( 
.A(n_911),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_883),
.B(n_543),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_927),
.B(n_675),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_927),
.B(n_675),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_927),
.B(n_976),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_L g1083 ( 
.A(n_883),
.B(n_406),
.C(n_404),
.Y(n_1083)
);

INVx5_ASAP7_75t_L g1084 ( 
.A(n_911),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_R g1085 ( 
.A(n_926),
.B(n_406),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_839),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_847),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_927),
.B(n_682),
.Y(n_1088)
);

OR2x2_ASAP7_75t_SL g1089 ( 
.A(n_907),
.B(n_546),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_911),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_898),
.A2(n_682),
.B1(n_712),
.B2(n_688),
.Y(n_1091)
);

NAND2xp33_ASAP7_75t_L g1092 ( 
.A(n_924),
.B(n_725),
.Y(n_1092)
);

NAND2xp33_ASAP7_75t_L g1093 ( 
.A(n_927),
.B(n_725),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_927),
.B(n_976),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_882),
.B(n_720),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_979),
.Y(n_1096)
);

INVx5_ASAP7_75t_L g1097 ( 
.A(n_978),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_955),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_853),
.A2(n_285),
.B1(n_682),
.B2(n_688),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_976),
.B(n_688),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_960),
.B(n_725),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_826),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_976),
.B(n_712),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_976),
.B(n_712),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_827),
.B(n_635),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_909),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_976),
.B(n_721),
.Y(n_1107)
);

INVx6_ASAP7_75t_L g1108 ( 
.A(n_843),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_898),
.A2(n_721),
.B1(n_738),
.B2(n_722),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_828),
.B(n_643),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_889),
.B(n_960),
.Y(n_1111)
);

AND2x6_ASAP7_75t_SL g1112 ( 
.A(n_929),
.B(n_643),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_842),
.B(n_721),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_929),
.B(n_720),
.Y(n_1114)
);

INVxp67_ASAP7_75t_L g1115 ( 
.A(n_873),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_SL g1116 ( 
.A1(n_898),
.A2(n_415),
.B1(n_409),
.B2(n_411),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_849),
.A2(n_705),
.B(n_696),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_975),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_980),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_914),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_849),
.A2(n_705),
.B(n_696),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_931),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_892),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_969),
.B(n_646),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_934),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_912),
.A2(n_722),
.B1(n_738),
.B2(n_762),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_964),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_853),
.A2(n_442),
.B1(n_437),
.B2(n_413),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_965),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_941),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_925),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_969),
.B(n_646),
.Y(n_1132)
);

OR2x6_ASAP7_75t_L g1133 ( 
.A(n_871),
.B(n_634),
.Y(n_1133)
);

NOR2x1_ASAP7_75t_R g1134 ( 
.A(n_868),
.B(n_427),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_971),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_930),
.B(n_762),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_946),
.B(n_412),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_936),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_972),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_862),
.A2(n_715),
.B(n_762),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_SL g1141 ( 
.A1(n_930),
.A2(n_432),
.B1(n_437),
.B2(n_433),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_837),
.B(n_722),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_959),
.B(n_412),
.Y(n_1143)
);

AND2x6_ASAP7_75t_SL g1144 ( 
.A(n_942),
.B(n_952),
.Y(n_1144)
);

INVx8_ASAP7_75t_L g1145 ( 
.A(n_877),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_837),
.B(n_671),
.Y(n_1146)
);

OR2x6_ASAP7_75t_L g1147 ( 
.A(n_851),
.B(n_634),
.Y(n_1147)
);

NOR2x2_ASAP7_75t_L g1148 ( 
.A(n_959),
.B(n_432),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_867),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_886),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_942),
.B(n_416),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_872),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_875),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_880),
.B(n_923),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_874),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_888),
.B(n_671),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_978),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_895),
.B(n_691),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_901),
.B(n_691),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1092),
.A2(n_947),
.B(n_939),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1062),
.A2(n_905),
.B(n_903),
.C(n_910),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_983),
.B(n_932),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1066),
.B(n_885),
.Y(n_1163)
);

O2A1O1Ixp5_ASAP7_75t_L g1164 ( 
.A1(n_1073),
.A2(n_830),
.B(n_977),
.C(n_945),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_1157),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1079),
.B(n_881),
.Y(n_1166)
);

NAND2x1p5_ASAP7_75t_L g1167 ( 
.A(n_1097),
.B(n_830),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1111),
.B(n_933),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1047),
.B(n_654),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1012),
.A2(n_1094),
.B(n_1082),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_985),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_SL g1172 ( 
.A(n_1131),
.B(n_420),
.C(n_416),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_988),
.A2(n_957),
.B(n_917),
.C(n_920),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_1157),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1021),
.B(n_966),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1082),
.A2(n_949),
.B(n_948),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_988),
.A2(n_977),
.B(n_902),
.C(n_775),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_993),
.A2(n_659),
.B(n_968),
.C(n_958),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_SL g1179 ( 
.A(n_1151),
.B(n_420),
.C(n_424),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_993),
.A2(n_958),
.B(n_962),
.C(n_963),
.Y(n_1180)
);

AOI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1101),
.A2(n_937),
.B(n_715),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1094),
.A2(n_743),
.B(n_714),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1086),
.Y(n_1183)
);

OAI21xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1146),
.A2(n_636),
.B(n_642),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_R g1185 ( 
.A(n_992),
.B(n_424),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_986),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_1068),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1026),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1116),
.A2(n_285),
.B1(n_426),
.B2(n_440),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1093),
.A2(n_743),
.B(n_714),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1035),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_1006),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1146),
.A2(n_426),
.B1(n_440),
.B2(n_441),
.Y(n_1193)
);

OA21x2_ASAP7_75t_L g1194 ( 
.A1(n_984),
.A2(n_636),
.B(n_642),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_990),
.Y(n_1195)
);

INVx1_ASAP7_75t_SL g1196 ( 
.A(n_1027),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1034),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1083),
.A2(n_441),
.B(n_443),
.C(n_444),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1024),
.B(n_443),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_SL g1200 ( 
.A(n_1085),
.B(n_326),
.C(n_317),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1038),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1023),
.B(n_299),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1023),
.A2(n_285),
.B1(n_367),
.B2(n_366),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1037),
.Y(n_1204)
);

OAI21xp33_ASAP7_75t_L g1205 ( 
.A1(n_1054),
.A2(n_1141),
.B(n_1017),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_981),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1118),
.B(n_691),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1119),
.B(n_1150),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_999),
.B(n_306),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1040),
.B(n_691),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1102),
.Y(n_1211)
);

OA22x2_ASAP7_75t_L g1212 ( 
.A1(n_1143),
.A2(n_1015),
.B1(n_1011),
.B2(n_1128),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_984),
.A2(n_374),
.B(n_313),
.Y(n_1213)
);

OAI22x1_ASAP7_75t_L g1214 ( 
.A1(n_1008),
.A2(n_327),
.B1(n_328),
.B2(n_335),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1020),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1056),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1060),
.Y(n_1217)
);

AO32x1_ASAP7_75t_L g1218 ( 
.A1(n_1130),
.A2(n_1128),
.A3(n_1013),
.B1(n_991),
.B2(n_1019),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_982),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1045),
.A2(n_743),
.B(n_714),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1072),
.A2(n_743),
.B(n_714),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1028),
.B(n_337),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1025),
.B(n_344),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1114),
.B(n_691),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1064),
.Y(n_1225)
);

OR2x6_ASAP7_75t_SL g1226 ( 
.A(n_1041),
.B(n_346),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1036),
.A2(n_285),
.B(n_1),
.C(n_4),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1156),
.A2(n_743),
.B(n_714),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1136),
.B(n_1149),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1046),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1071),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1115),
.B(n_354),
.Y(n_1232)
);

OAI21xp33_ASAP7_75t_L g1233 ( 
.A1(n_1059),
.A2(n_384),
.B(n_403),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1157),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1052),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1152),
.B(n_711),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1155),
.B(n_711),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1055),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1089),
.B(n_355),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1097),
.B(n_356),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_989),
.B(n_357),
.Y(n_1241)
);

O2A1O1Ixp5_ASAP7_75t_L g1242 ( 
.A1(n_1074),
.A2(n_711),
.B(n_394),
.C(n_391),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1058),
.A2(n_390),
.B1(n_388),
.B2(n_387),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1036),
.A2(n_0),
.B(n_1),
.C(n_5),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1139),
.B(n_363),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1156),
.A2(n_386),
.B(n_385),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1033),
.A2(n_381),
.B1(n_376),
.B2(n_375),
.Y(n_1247)
);

OAI21xp33_ASAP7_75t_L g1248 ( 
.A1(n_1059),
.A2(n_365),
.B(n_364),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1051),
.B(n_6),
.Y(n_1249)
);

AOI21x1_ASAP7_75t_L g1250 ( 
.A1(n_997),
.A2(n_227),
.B(n_221),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1098),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1002),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1097),
.B(n_219),
.Y(n_1253)
);

NOR3xp33_ASAP7_75t_L g1254 ( 
.A(n_1134),
.B(n_11),
.C(n_13),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_R g1255 ( 
.A(n_1050),
.B(n_218),
.Y(n_1255)
);

NOR2xp67_ASAP7_75t_L g1256 ( 
.A(n_1153),
.B(n_216),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1016),
.B(n_11),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1057),
.B(n_13),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1008),
.B(n_16),
.Y(n_1259)
);

BUFx8_ASAP7_75t_L g1260 ( 
.A(n_1061),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1051),
.B(n_1069),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1105),
.B(n_17),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1058),
.A2(n_199),
.B1(n_195),
.B2(n_186),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1048),
.A2(n_17),
.B(n_21),
.C(n_22),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1158),
.A2(n_165),
.B(n_154),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1158),
.A2(n_141),
.B(n_128),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_1042),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_994),
.B(n_122),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1070),
.B(n_21),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1154),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1069),
.B(n_23),
.Y(n_1271)
);

AO21x1_ASAP7_75t_L g1272 ( 
.A1(n_1067),
.A2(n_24),
.B(n_25),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1154),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1106),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1097),
.B(n_994),
.Y(n_1275)
);

OA22x2_ASAP7_75t_L g1276 ( 
.A1(n_1148),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_1276)
);

OAI21xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1142),
.A2(n_30),
.B(n_31),
.Y(n_1277)
);

NOR2x1_ASAP7_75t_L g1278 ( 
.A(n_1007),
.B(n_121),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1105),
.B(n_119),
.Y(n_1279)
);

NAND3xp33_ASAP7_75t_SL g1280 ( 
.A(n_1137),
.B(n_33),
.C(n_34),
.Y(n_1280)
);

NAND2x1_ASAP7_75t_L g1281 ( 
.A(n_1031),
.B(n_115),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1110),
.B(n_111),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1127),
.B(n_35),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1065),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1159),
.A2(n_90),
.B(n_107),
.Y(n_1285)
);

AND3x4_ASAP7_75t_L g1286 ( 
.A(n_1087),
.B(n_36),
.C(n_37),
.Y(n_1286)
);

NOR3xp33_ASAP7_75t_SL g1287 ( 
.A(n_1138),
.B(n_1123),
.C(n_1003),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1159),
.A2(n_110),
.B(n_105),
.Y(n_1288)
);

CKINVDCx10_ASAP7_75t_R g1289 ( 
.A(n_1032),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1142),
.A2(n_1063),
.B(n_1067),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1063),
.A2(n_102),
.B(n_100),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1110),
.B(n_98),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1077),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1053),
.A2(n_85),
.B(n_83),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1129),
.B(n_36),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1120),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1007),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1135),
.B(n_38),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1029),
.A2(n_81),
.B1(n_79),
.B2(n_74),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1122),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1112),
.B(n_41),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1048),
.A2(n_46),
.B1(n_48),
.B2(n_53),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1124),
.B(n_55),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1080),
.A2(n_56),
.B(n_58),
.Y(n_1304)
);

INVxp67_ASAP7_75t_L g1305 ( 
.A(n_1124),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1132),
.B(n_59),
.Y(n_1306)
);

BUFx8_ASAP7_75t_SL g1307 ( 
.A(n_1133),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1096),
.Y(n_1308)
);

NOR2x1_ASAP7_75t_L g1309 ( 
.A(n_1004),
.B(n_60),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1000),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1020),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1095),
.A2(n_60),
.B1(n_63),
.B2(n_65),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1125),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_SL g1314 ( 
.A1(n_1049),
.A2(n_65),
.B(n_72),
.C(n_73),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1170),
.A2(n_1076),
.B(n_1018),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1174),
.Y(n_1316)
);

CKINVDCx11_ASAP7_75t_R g1317 ( 
.A(n_1226),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1290),
.A2(n_1140),
.B(n_1113),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1162),
.B(n_1144),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1310),
.B(n_1000),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1169),
.B(n_1132),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1183),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1229),
.A2(n_1099),
.B1(n_1030),
.B2(n_1010),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_1206),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1182),
.A2(n_1080),
.B(n_1107),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1228),
.A2(n_1081),
.B(n_1088),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1170),
.A2(n_1078),
.B(n_1018),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1199),
.B(n_1147),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1215),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1289),
.Y(n_1330)
);

NOR2xp67_ASAP7_75t_L g1331 ( 
.A(n_1192),
.B(n_1014),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1251),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1166),
.B(n_1261),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1160),
.A2(n_1104),
.B(n_1103),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1175),
.B(n_1001),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1294),
.A2(n_1104),
.B(n_1103),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1176),
.A2(n_1100),
.B(n_1113),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1176),
.A2(n_1100),
.B(n_1121),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1260),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1215),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1171),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1181),
.A2(n_1221),
.B(n_1220),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_R g1343 ( 
.A(n_1200),
.B(n_998),
.Y(n_1343)
);

AO22x2_ASAP7_75t_L g1344 ( 
.A1(n_1280),
.A2(n_1302),
.B1(n_1312),
.B2(n_1286),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1270),
.B(n_1147),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1187),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1208),
.B(n_1108),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1305),
.B(n_1030),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1220),
.A2(n_1221),
.B(n_1190),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1190),
.A2(n_1121),
.B(n_1117),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1165),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1215),
.Y(n_1352)
);

NAND2x1p5_ASAP7_75t_L g1353 ( 
.A(n_1297),
.B(n_1084),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1186),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1195),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1205),
.A2(n_1108),
.B1(n_1147),
.B2(n_1145),
.Y(n_1356)
);

NOR4xp25_ASAP7_75t_L g1357 ( 
.A(n_1244),
.B(n_1001),
.C(n_996),
.D(n_995),
.Y(n_1357)
);

INVx6_ASAP7_75t_L g1358 ( 
.A(n_1260),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1272),
.A2(n_1117),
.A3(n_1009),
.B(n_1005),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1196),
.B(n_1078),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1241),
.A2(n_1108),
.B1(n_1145),
.B2(n_1133),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1273),
.B(n_1133),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1307),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1223),
.A2(n_1239),
.B1(n_1202),
.B2(n_1209),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1197),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1164),
.A2(n_1075),
.B(n_1109),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1210),
.A2(n_1091),
.B(n_1044),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1291),
.A2(n_1126),
.B(n_1039),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1291),
.A2(n_1090),
.B(n_1022),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1194),
.A2(n_1090),
.B(n_1031),
.Y(n_1370)
);

NAND2xp33_ASAP7_75t_L g1371 ( 
.A(n_1201),
.B(n_1020),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1194),
.A2(n_1031),
.B(n_1084),
.Y(n_1372)
);

AND3x2_ASAP7_75t_L g1373 ( 
.A(n_1254),
.B(n_1032),
.C(n_1145),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1165),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1211),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1249),
.B(n_1031),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1271),
.B(n_1043),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1168),
.A2(n_1161),
.B(n_1257),
.C(n_1259),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1161),
.A2(n_1179),
.B(n_1178),
.C(n_1189),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1177),
.A2(n_1180),
.B(n_1173),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1178),
.A2(n_987),
.B(n_1078),
.C(n_1043),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1219),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1268),
.A2(n_987),
.B1(n_1078),
.B2(n_1043),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1230),
.B(n_987),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1268),
.B(n_73),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1177),
.A2(n_1180),
.B(n_1242),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1232),
.A2(n_1292),
.B1(n_1282),
.B2(n_1279),
.Y(n_1387)
);

NOR2x1_ASAP7_75t_SL g1388 ( 
.A(n_1275),
.B(n_1253),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1306),
.B(n_1262),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1235),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_SL g1391 ( 
.A(n_1185),
.B(n_1188),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1238),
.B(n_1284),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1173),
.A2(n_1207),
.B(n_1237),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1277),
.A2(n_1285),
.B(n_1265),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1213),
.A2(n_1303),
.B(n_1252),
.C(n_1295),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1293),
.Y(n_1396)
);

AO31x2_ASAP7_75t_L g1397 ( 
.A1(n_1263),
.A2(n_1288),
.A3(n_1266),
.B(n_1265),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1287),
.Y(n_1398)
);

O2A1O1Ixp5_ASAP7_75t_L g1399 ( 
.A1(n_1246),
.A2(n_1298),
.B(n_1283),
.C(n_1240),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_SL g1400 ( 
.A1(n_1280),
.A2(n_1301),
.B(n_1203),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1167),
.A2(n_1299),
.B(n_1236),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1258),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1308),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1191),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1204),
.B(n_1217),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1234),
.B(n_1296),
.Y(n_1406)
);

AOI221xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1244),
.A2(n_1227),
.B1(n_1264),
.B2(n_1248),
.C(n_1233),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1216),
.B(n_1300),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1245),
.B(n_1269),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1225),
.B(n_1274),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1250),
.A2(n_1281),
.B(n_1278),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1297),
.A2(n_1314),
.B(n_1256),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1212),
.A2(n_1304),
.B(n_1198),
.Y(n_1413)
);

INVx4_ASAP7_75t_L g1414 ( 
.A(n_1311),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1231),
.B(n_1313),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1218),
.A2(n_1222),
.B(n_1214),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1227),
.A2(n_1309),
.B(n_1304),
.C(n_1264),
.Y(n_1417)
);

BUFx5_ASAP7_75t_L g1418 ( 
.A(n_1311),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1243),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1276),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1200),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1255),
.Y(n_1422)
);

O2A1O1Ixp5_ASAP7_75t_L g1423 ( 
.A1(n_1193),
.A2(n_1218),
.B(n_1247),
.C(n_1276),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1218),
.A2(n_1267),
.B(n_1172),
.Y(n_1424)
);

A2O1A1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1163),
.A2(n_1111),
.B(n_1151),
.C(n_1066),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_1260),
.Y(n_1426)
);

CKINVDCx16_ASAP7_75t_R g1427 ( 
.A(n_1185),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1206),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1170),
.A2(n_1092),
.B(n_1012),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1170),
.A2(n_1092),
.B(n_1012),
.Y(n_1430)
);

AO21x1_ASAP7_75t_L g1431 ( 
.A1(n_1163),
.A2(n_1073),
.B(n_1111),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1268),
.B(n_1270),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1310),
.B(n_1166),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1170),
.A2(n_1092),
.B(n_1012),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1171),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1162),
.B(n_836),
.Y(n_1436)
);

AOI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1224),
.A2(n_1181),
.B(n_1176),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1171),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1290),
.A2(n_1164),
.B(n_1184),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1310),
.B(n_1166),
.Y(n_1440)
);

AND2x2_ASAP7_75t_SL g1441 ( 
.A(n_1163),
.B(n_1017),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1169),
.B(n_823),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1169),
.B(n_823),
.Y(n_1443)
);

AND2x6_ASAP7_75t_SL g1444 ( 
.A(n_1301),
.B(n_1241),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1162),
.B(n_836),
.Y(n_1445)
);

O2A1O1Ixp5_ASAP7_75t_L g1446 ( 
.A1(n_1163),
.A2(n_1111),
.B(n_1073),
.C(n_1151),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1182),
.A2(n_984),
.B(n_1228),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1163),
.A2(n_1111),
.B(n_1151),
.C(n_1066),
.Y(n_1448)
);

AOI211x1_ASAP7_75t_L g1449 ( 
.A1(n_1205),
.A2(n_1163),
.B(n_1272),
.C(n_865),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1162),
.B(n_836),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1169),
.B(n_823),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1310),
.B(n_1166),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1310),
.B(n_1166),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1310),
.B(n_1166),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1182),
.A2(n_984),
.B(n_1228),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1290),
.A2(n_1164),
.B(n_1184),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1215),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1310),
.B(n_1166),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1183),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_L g1460 ( 
.A(n_1163),
.B(n_1111),
.C(n_1151),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1310),
.B(n_1166),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1215),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1182),
.A2(n_984),
.B(n_1228),
.Y(n_1463)
);

NAND2xp33_ASAP7_75t_L g1464 ( 
.A(n_1163),
.B(n_1205),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1305),
.B(n_1270),
.Y(n_1465)
);

AOI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1224),
.A2(n_1181),
.B(n_1176),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1182),
.A2(n_984),
.B(n_1228),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1169),
.B(n_823),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1392),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1346),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1439),
.A2(n_1456),
.B(n_1394),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1389),
.B(n_1321),
.Y(n_1472)
);

OA21x2_ASAP7_75t_L g1473 ( 
.A1(n_1439),
.A2(n_1456),
.B(n_1394),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1460),
.A2(n_1464),
.B1(n_1344),
.B2(n_1441),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1392),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1460),
.B(n_1436),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1330),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1425),
.B(n_1448),
.C(n_1364),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1432),
.B(n_1355),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1396),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1427),
.Y(n_1481)
);

AO31x2_ASAP7_75t_L g1482 ( 
.A1(n_1431),
.A2(n_1417),
.A3(n_1416),
.B(n_1395),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1375),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1447),
.A2(n_1463),
.B(n_1455),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1332),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1467),
.A2(n_1342),
.B(n_1349),
.Y(n_1486)
);

INVx4_ASAP7_75t_L g1487 ( 
.A(n_1340),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1426),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_SL g1489 ( 
.A1(n_1388),
.A2(n_1412),
.B(n_1424),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1442),
.B(n_1443),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1451),
.B(n_1468),
.Y(n_1491)
);

O2A1O1Ixp5_ASAP7_75t_L g1492 ( 
.A1(n_1446),
.A2(n_1380),
.B(n_1413),
.C(n_1379),
.Y(n_1492)
);

BUFx2_ASAP7_75t_R g1493 ( 
.A(n_1398),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1346),
.B(n_1324),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1341),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1354),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1365),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1344),
.A2(n_1409),
.B1(n_1445),
.B2(n_1450),
.Y(n_1498)
);

O2A1O1Ixp5_ASAP7_75t_L g1499 ( 
.A1(n_1380),
.A2(n_1413),
.B(n_1378),
.C(n_1423),
.Y(n_1499)
);

OA21x2_ASAP7_75t_L g1500 ( 
.A1(n_1386),
.A2(n_1318),
.B(n_1338),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1350),
.A2(n_1370),
.B(n_1334),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1382),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1322),
.B(n_1459),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1369),
.A2(n_1466),
.B(n_1437),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1390),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1420),
.A2(n_1421),
.B1(n_1335),
.B2(n_1419),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1326),
.A2(n_1336),
.B(n_1325),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1403),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1387),
.A2(n_1432),
.B1(n_1333),
.B2(n_1461),
.Y(n_1509)
);

BUFx12f_ASAP7_75t_L g1510 ( 
.A(n_1358),
.Y(n_1510)
);

O2A1O1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1400),
.A2(n_1335),
.B(n_1391),
.C(n_1319),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1318),
.A2(n_1366),
.B(n_1393),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1353),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1402),
.B(n_1385),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1435),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1337),
.A2(n_1372),
.B(n_1411),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1315),
.A2(n_1327),
.B(n_1368),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1421),
.A2(n_1333),
.B1(n_1328),
.B2(n_1385),
.Y(n_1518)
);

CKINVDCx6p67_ASAP7_75t_R g1519 ( 
.A(n_1339),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1438),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1428),
.Y(n_1521)
);

NAND2x1p5_ASAP7_75t_L g1522 ( 
.A(n_1360),
.B(n_1316),
.Y(n_1522)
);

OR2x6_ASAP7_75t_L g1523 ( 
.A(n_1449),
.B(n_1401),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1353),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_1347),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1407),
.A2(n_1399),
.B(n_1381),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1433),
.B(n_1440),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1363),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1405),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_SL g1530 ( 
.A1(n_1320),
.A2(n_1377),
.B(n_1461),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1433),
.B(n_1453),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1351),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1405),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1407),
.A2(n_1376),
.B(n_1377),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1408),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1408),
.Y(n_1536)
);

INVx4_ASAP7_75t_SL g1537 ( 
.A(n_1421),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1440),
.A2(n_1458),
.B1(n_1452),
.B2(n_1453),
.Y(n_1538)
);

OR2x6_ASAP7_75t_L g1539 ( 
.A(n_1383),
.B(n_1345),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1404),
.Y(n_1540)
);

CKINVDCx6p67_ASAP7_75t_R g1541 ( 
.A(n_1317),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1358),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1452),
.B(n_1454),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_SL g1544 ( 
.A1(n_1454),
.A2(n_1384),
.B(n_1356),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1415),
.Y(n_1545)
);

OAI211xp5_ASAP7_75t_L g1546 ( 
.A1(n_1357),
.A2(n_1361),
.B(n_1343),
.C(n_1362),
.Y(n_1546)
);

O2A1O1Ixp5_ASAP7_75t_L g1547 ( 
.A1(n_1323),
.A2(n_1383),
.B(n_1384),
.C(n_1348),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1415),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1367),
.A2(n_1410),
.B(n_1351),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1465),
.B(n_1406),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1465),
.B(n_1444),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1371),
.A2(n_1367),
.B(n_1357),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1374),
.Y(n_1553)
);

INVxp67_ASAP7_75t_SL g1554 ( 
.A(n_1331),
.Y(n_1554)
);

INVxp67_ASAP7_75t_L g1555 ( 
.A(n_1462),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1340),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1422),
.A2(n_1373),
.B1(n_1329),
.B2(n_1414),
.Y(n_1557)
);

A2O1A1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1397),
.A2(n_1359),
.B(n_1352),
.C(n_1457),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1352),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1397),
.A2(n_1418),
.B(n_1414),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1418),
.A2(n_1329),
.B(n_1352),
.Y(n_1561)
);

AO21x2_ASAP7_75t_L g1562 ( 
.A1(n_1418),
.A2(n_1457),
.B(n_1462),
.Y(n_1562)
);

AO31x2_ASAP7_75t_L g1563 ( 
.A1(n_1418),
.A2(n_1431),
.A3(n_1417),
.B(n_1416),
.Y(n_1563)
);

OA21x2_ASAP7_75t_L g1564 ( 
.A1(n_1418),
.A2(n_1456),
.B(n_1439),
.Y(n_1564)
);

NAND2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1462),
.B(n_1174),
.Y(n_1565)
);

O2A1O1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1425),
.A2(n_1448),
.B(n_1464),
.C(n_1400),
.Y(n_1566)
);

O2A1O1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1425),
.A2(n_1448),
.B(n_1464),
.C(n_1400),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1332),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1353),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1442),
.B(n_1443),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1425),
.A2(n_1448),
.B1(n_1460),
.B2(n_1436),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1332),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1442),
.B(n_1443),
.Y(n_1573)
);

AO31x2_ASAP7_75t_L g1574 ( 
.A1(n_1431),
.A2(n_1417),
.A3(n_1416),
.B(n_1425),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1392),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1439),
.A2(n_1456),
.B(n_1394),
.Y(n_1576)
);

NAND2x1p5_ASAP7_75t_L g1577 ( 
.A(n_1360),
.B(n_1174),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1439),
.A2(n_1456),
.B(n_1394),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1442),
.B(n_1443),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1392),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1430),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1460),
.B(n_1436),
.Y(n_1582)
);

OAI21x1_ASAP7_75t_L g1583 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1430),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1432),
.B(n_1355),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1442),
.B(n_1443),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1442),
.B(n_1443),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1430),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1351),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1351),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1430),
.Y(n_1590)
);

INVx3_ASAP7_75t_L g1591 ( 
.A(n_1353),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1430),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1392),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1442),
.B(n_1443),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1392),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1346),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1460),
.B(n_1436),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1355),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1355),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1355),
.Y(n_1600)
);

NAND2x1p5_ASAP7_75t_L g1601 ( 
.A(n_1360),
.B(n_1174),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1353),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1355),
.Y(n_1603)
);

OAI221xp5_ASAP7_75t_L g1604 ( 
.A1(n_1364),
.A2(n_1460),
.B1(n_1448),
.B2(n_1425),
.C(n_1400),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1432),
.B(n_1355),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1392),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1430),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1332),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1389),
.B(n_1321),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1460),
.A2(n_1464),
.B1(n_1163),
.B2(n_1111),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1460),
.A2(n_1464),
.B1(n_1163),
.B2(n_1111),
.Y(n_1611)
);

O2A1O1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1425),
.A2(n_1448),
.B(n_1464),
.C(n_1400),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1355),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_SL g1614 ( 
.A1(n_1388),
.A2(n_1272),
.B(n_1412),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_SL g1615 ( 
.A1(n_1319),
.A2(n_789),
.B1(n_672),
.B2(n_1436),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1392),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1432),
.B(n_1355),
.Y(n_1617)
);

O2A1O1Ixp33_ASAP7_75t_SL g1618 ( 
.A1(n_1425),
.A2(n_1448),
.B(n_1395),
.C(n_1252),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1392),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1330),
.Y(n_1620)
);

OA22x2_ASAP7_75t_L g1621 ( 
.A1(n_1546),
.A2(n_1571),
.B1(n_1544),
.B2(n_1615),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_SL g1622 ( 
.A1(n_1511),
.A2(n_1567),
.B(n_1566),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1527),
.B(n_1531),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1498),
.A2(n_1474),
.B1(n_1611),
.B2(n_1610),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1494),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1472),
.B(n_1609),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1498),
.A2(n_1474),
.B1(n_1610),
.B2(n_1611),
.Y(n_1627)
);

A2O1A1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1612),
.A2(n_1478),
.B(n_1597),
.C(n_1582),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_SL g1629 ( 
.A1(n_1509),
.A2(n_1582),
.B(n_1476),
.Y(n_1629)
);

OA21x2_ASAP7_75t_L g1630 ( 
.A1(n_1552),
.A2(n_1504),
.B(n_1492),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1538),
.B(n_1543),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1477),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1476),
.A2(n_1597),
.B1(n_1525),
.B2(n_1518),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1490),
.B(n_1491),
.Y(n_1634)
);

AND2x2_ASAP7_75t_SL g1635 ( 
.A(n_1471),
.B(n_1473),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1518),
.A2(n_1604),
.B1(n_1506),
.B2(n_1538),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1543),
.B(n_1570),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1554),
.A2(n_1573),
.B1(n_1594),
.B2(n_1585),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1579),
.B(n_1586),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_SL g1640 ( 
.A1(n_1471),
.A2(n_1576),
.B(n_1473),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1470),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1503),
.B(n_1596),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1479),
.B(n_1584),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1495),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1539),
.A2(n_1557),
.B1(n_1584),
.B2(n_1605),
.Y(n_1645)
);

AOI21x1_ASAP7_75t_SL g1646 ( 
.A1(n_1479),
.A2(n_1605),
.B(n_1584),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1496),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1618),
.A2(n_1499),
.B(n_1547),
.C(n_1530),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1539),
.A2(n_1617),
.B1(n_1480),
.B2(n_1551),
.Y(n_1649)
);

O2A1O1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1614),
.A2(n_1558),
.B(n_1521),
.C(n_1489),
.Y(n_1650)
);

AOI21x1_ASAP7_75t_SL g1651 ( 
.A1(n_1514),
.A2(n_1537),
.B(n_1574),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1497),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1550),
.B(n_1469),
.Y(n_1653)
);

O2A1O1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1475),
.A2(n_1580),
.B(n_1619),
.C(n_1616),
.Y(n_1654)
);

NOR2xp67_ASAP7_75t_L g1655 ( 
.A(n_1568),
.B(n_1608),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1539),
.A2(n_1551),
.B1(n_1575),
.B2(n_1606),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1485),
.B(n_1493),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1542),
.B(n_1528),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1572),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1593),
.B(n_1595),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1620),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1572),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1523),
.A2(n_1522),
.B1(n_1577),
.B2(n_1601),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1523),
.A2(n_1522),
.B1(n_1577),
.B2(n_1601),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1502),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1529),
.B(n_1533),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1620),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1535),
.B(n_1536),
.Y(n_1668)
);

O2A1O1Ixp33_ASAP7_75t_L g1669 ( 
.A1(n_1505),
.A2(n_1515),
.B(n_1520),
.C(n_1508),
.Y(n_1669)
);

OA21x2_ASAP7_75t_L g1670 ( 
.A1(n_1581),
.A2(n_1583),
.B(n_1607),
.Y(n_1670)
);

O2A1O1Ixp5_ASAP7_75t_L g1671 ( 
.A1(n_1532),
.A2(n_1613),
.B(n_1603),
.C(n_1600),
.Y(n_1671)
);

AOI21x1_ASAP7_75t_SL g1672 ( 
.A1(n_1537),
.A2(n_1574),
.B(n_1482),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1559),
.Y(n_1673)
);

AND2x2_ASAP7_75t_SL g1674 ( 
.A(n_1578),
.B(n_1526),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1598),
.B(n_1599),
.Y(n_1675)
);

AOI21x1_ASAP7_75t_SL g1676 ( 
.A1(n_1574),
.A2(n_1482),
.B(n_1563),
.Y(n_1676)
);

NAND2x1p5_ASAP7_75t_L g1677 ( 
.A(n_1560),
.B(n_1564),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1548),
.B(n_1545),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1483),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1540),
.A2(n_1553),
.B(n_1526),
.C(n_1555),
.Y(n_1680)
);

CKINVDCx16_ASAP7_75t_R g1681 ( 
.A(n_1510),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1540),
.B(n_1534),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1534),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1519),
.A2(n_1481),
.B1(n_1541),
.B2(n_1510),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1588),
.B(n_1589),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1541),
.A2(n_1602),
.B1(n_1513),
.B2(n_1524),
.Y(n_1686)
);

O2A1O1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1526),
.A2(n_1534),
.B(n_1589),
.C(n_1588),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1482),
.B(n_1563),
.Y(n_1688)
);

OA21x2_ASAP7_75t_L g1689 ( 
.A1(n_1587),
.A2(n_1592),
.B(n_1590),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1565),
.A2(n_1487),
.B(n_1512),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1513),
.B(n_1602),
.Y(n_1691)
);

CKINVDCx11_ASAP7_75t_R g1692 ( 
.A(n_1556),
.Y(n_1692)
);

AOI21x1_ASAP7_75t_SL g1693 ( 
.A1(n_1563),
.A2(n_1560),
.B(n_1517),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1562),
.B(n_1591),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1549),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1569),
.B(n_1561),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1561),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_SL g1698 ( 
.A1(n_1500),
.A2(n_1488),
.B(n_1477),
.Y(n_1698)
);

OA21x2_ASAP7_75t_L g1699 ( 
.A1(n_1507),
.A2(n_1501),
.B(n_1484),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1569),
.B(n_1500),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1516),
.B(n_1486),
.Y(n_1701)
);

AOI21x1_ASAP7_75t_SL g1702 ( 
.A1(n_1516),
.A2(n_1163),
.B(n_1335),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1527),
.B(n_1531),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1498),
.A2(n_1364),
.B1(n_1460),
.B2(n_1615),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1572),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1494),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1498),
.A2(n_1364),
.B1(n_1460),
.B2(n_1615),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1498),
.A2(n_1364),
.B1(n_1460),
.B2(n_1615),
.Y(n_1708)
);

A2O1A1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1566),
.A2(n_1111),
.B(n_1612),
.C(n_1567),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1472),
.B(n_1609),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1498),
.A2(n_1364),
.B1(n_1460),
.B2(n_1615),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1527),
.B(n_1531),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1572),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1472),
.B(n_1609),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1494),
.Y(n_1715)
);

OA21x2_ASAP7_75t_L g1716 ( 
.A1(n_1552),
.A2(n_1504),
.B(n_1492),
.Y(n_1716)
);

OA21x2_ASAP7_75t_L g1717 ( 
.A1(n_1552),
.A2(n_1504),
.B(n_1492),
.Y(n_1717)
);

BUFx3_ASAP7_75t_L g1718 ( 
.A(n_1572),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1472),
.B(n_1609),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_SL g1720 ( 
.A1(n_1511),
.A2(n_1448),
.B(n_1425),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_SL g1721 ( 
.A1(n_1511),
.A2(n_1448),
.B(n_1425),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1498),
.A2(n_1364),
.B1(n_1460),
.B2(n_1615),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1494),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1472),
.B(n_1609),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1498),
.A2(n_1364),
.B1(n_1460),
.B2(n_1615),
.Y(n_1725)
);

O2A1O1Ixp33_ASAP7_75t_L g1726 ( 
.A1(n_1571),
.A2(n_1448),
.B(n_1425),
.C(n_1464),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1527),
.B(n_1531),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1472),
.B(n_1609),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1572),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1527),
.B(n_1531),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1472),
.B(n_1609),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1527),
.B(n_1531),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1682),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1625),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1647),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1696),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1706),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1715),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1634),
.B(n_1723),
.Y(n_1739)
);

BUFx2_ASAP7_75t_L g1740 ( 
.A(n_1694),
.Y(n_1740)
);

OAI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1704),
.A2(n_1707),
.B1(n_1708),
.B2(n_1725),
.Y(n_1741)
);

INVxp67_ASAP7_75t_SL g1742 ( 
.A(n_1654),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1695),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1713),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1709),
.A2(n_1726),
.B(n_1721),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_1729),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1635),
.B(n_1674),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1697),
.B(n_1700),
.Y(n_1748)
);

OR2x6_ASAP7_75t_L g1749 ( 
.A(n_1698),
.B(n_1640),
.Y(n_1749)
);

AO21x1_ASAP7_75t_SL g1750 ( 
.A1(n_1688),
.A2(n_1631),
.B(n_1683),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1639),
.B(n_1623),
.Y(n_1751)
);

INVx2_ASAP7_75t_SL g1752 ( 
.A(n_1652),
.Y(n_1752)
);

BUFx2_ASAP7_75t_L g1753 ( 
.A(n_1677),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1703),
.B(n_1712),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1701),
.Y(n_1755)
);

AO21x2_ASAP7_75t_L g1756 ( 
.A1(n_1687),
.A2(n_1680),
.B(n_1690),
.Y(n_1756)
);

AO21x2_ASAP7_75t_L g1757 ( 
.A1(n_1687),
.A2(n_1680),
.B(n_1720),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1677),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1732),
.B(n_1727),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1665),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1699),
.Y(n_1761)
);

AO21x2_ASAP7_75t_L g1762 ( 
.A1(n_1624),
.A2(n_1627),
.B(n_1648),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1730),
.B(n_1637),
.Y(n_1763)
);

AO21x2_ASAP7_75t_L g1764 ( 
.A1(n_1648),
.A2(n_1628),
.B(n_1629),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1671),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1638),
.B(n_1653),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1669),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1633),
.B(n_1660),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1644),
.B(n_1679),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1669),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1666),
.B(n_1668),
.Y(n_1771)
);

AOI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1711),
.A2(n_1722),
.B(n_1621),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1678),
.B(n_1642),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1643),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1656),
.B(n_1630),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1675),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1643),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1654),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1691),
.Y(n_1779)
);

OA21x2_ASAP7_75t_L g1780 ( 
.A1(n_1676),
.A2(n_1636),
.B(n_1693),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1626),
.B(n_1731),
.Y(n_1781)
);

OR2x6_ASAP7_75t_L g1782 ( 
.A(n_1622),
.B(n_1726),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1649),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1710),
.B(n_1719),
.Y(n_1784)
);

OR2x6_ASAP7_75t_L g1785 ( 
.A(n_1650),
.B(n_1664),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1641),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_1632),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1716),
.Y(n_1788)
);

OR2x6_ASAP7_75t_L g1789 ( 
.A(n_1663),
.B(n_1645),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1717),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1714),
.B(n_1728),
.Y(n_1791)
);

INVx3_ASAP7_75t_SL g1792 ( 
.A(n_1621),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_SL g1793 ( 
.A1(n_1686),
.A2(n_1684),
.B(n_1718),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1685),
.Y(n_1794)
);

BUFx2_ASAP7_75t_L g1795 ( 
.A(n_1753),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1748),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1747),
.B(n_1670),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1760),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_SL g1799 ( 
.A1(n_1745),
.A2(n_1657),
.B(n_1662),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1748),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1747),
.B(n_1689),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1741),
.B(n_1705),
.Y(n_1802)
);

INVx5_ASAP7_75t_SL g1803 ( 
.A(n_1764),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1748),
.Y(n_1804)
);

CKINVDCx8_ASAP7_75t_R g1805 ( 
.A(n_1782),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1748),
.Y(n_1806)
);

INVx4_ASAP7_75t_L g1807 ( 
.A(n_1782),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_1755),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1743),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1782),
.A2(n_1724),
.B1(n_1681),
.B2(n_1673),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1735),
.Y(n_1811)
);

INVxp67_ASAP7_75t_SL g1812 ( 
.A(n_1767),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1752),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1755),
.B(n_1705),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1733),
.B(n_1705),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1740),
.B(n_1659),
.Y(n_1816)
);

AOI21xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1782),
.A2(n_1764),
.B(n_1742),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1750),
.B(n_1659),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1750),
.B(n_1672),
.Y(n_1819)
);

INVx4_ASAP7_75t_L g1820 ( 
.A(n_1782),
.Y(n_1820)
);

AND2x2_ASAP7_75t_SL g1821 ( 
.A(n_1780),
.B(n_1646),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1738),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1761),
.B(n_1655),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1761),
.B(n_1702),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1779),
.B(n_1658),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1772),
.B(n_1692),
.Y(n_1826)
);

INVx4_ASAP7_75t_L g1827 ( 
.A(n_1764),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1775),
.B(n_1651),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1809),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_R g1830 ( 
.A(n_1826),
.B(n_1661),
.Y(n_1830)
);

AOI211xp5_ASAP7_75t_SL g1831 ( 
.A1(n_1817),
.A2(n_1799),
.B(n_1793),
.C(n_1826),
.Y(n_1831)
);

INVx1_ASAP7_75t_SL g1832 ( 
.A(n_1822),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1813),
.Y(n_1833)
);

OAI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1810),
.A2(n_1772),
.B1(n_1792),
.B2(n_1768),
.C(n_1766),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1796),
.B(n_1738),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1798),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1823),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1810),
.A2(n_1792),
.B1(n_1785),
.B2(n_1789),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1807),
.A2(n_1764),
.B1(n_1762),
.B2(n_1792),
.Y(n_1839)
);

INVxp67_ASAP7_75t_L g1840 ( 
.A(n_1825),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1816),
.B(n_1736),
.Y(n_1841)
);

OAI211xp5_ASAP7_75t_L g1842 ( 
.A1(n_1827),
.A2(n_1793),
.B(n_1763),
.C(n_1739),
.Y(n_1842)
);

NAND4xp25_ASAP7_75t_SL g1843 ( 
.A(n_1818),
.B(n_1751),
.C(n_1759),
.D(n_1754),
.Y(n_1843)
);

OAI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1805),
.A2(n_1785),
.B1(n_1789),
.B2(n_1749),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1807),
.A2(n_1762),
.B1(n_1789),
.B2(n_1785),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1807),
.A2(n_1762),
.B1(n_1789),
.B2(n_1785),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_SL g1847 ( 
.A1(n_1805),
.A2(n_1802),
.B1(n_1789),
.B2(n_1785),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_R g1848 ( 
.A(n_1805),
.B(n_1667),
.Y(n_1848)
);

BUFx3_ASAP7_75t_L g1849 ( 
.A(n_1814),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1802),
.A2(n_1783),
.B1(n_1778),
.B2(n_1749),
.Y(n_1850)
);

BUFx6f_ASAP7_75t_L g1851 ( 
.A(n_1821),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1796),
.B(n_1734),
.Y(n_1852)
);

OAI211xp5_ASAP7_75t_L g1853 ( 
.A1(n_1827),
.A2(n_1770),
.B(n_1767),
.C(n_1737),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1822),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_SL g1855 ( 
.A1(n_1825),
.A2(n_1786),
.B1(n_1787),
.B2(n_1746),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1815),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1815),
.B(n_1794),
.Y(n_1857)
);

AOI211xp5_ASAP7_75t_L g1858 ( 
.A1(n_1828),
.A2(n_1773),
.B(n_1775),
.C(n_1771),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1800),
.B(n_1758),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1804),
.B(n_1765),
.Y(n_1860)
);

AOI33xp33_ASAP7_75t_L g1861 ( 
.A1(n_1819),
.A2(n_1791),
.A3(n_1784),
.B1(n_1781),
.B2(n_1769),
.B3(n_1776),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1808),
.B(n_1744),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1821),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1812),
.A2(n_1762),
.B(n_1757),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1813),
.Y(n_1865)
);

AO21x2_ASAP7_75t_L g1866 ( 
.A1(n_1824),
.A2(n_1788),
.B(n_1790),
.Y(n_1866)
);

BUFx2_ASAP7_75t_L g1867 ( 
.A(n_1795),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1806),
.B(n_1765),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1807),
.A2(n_1777),
.B1(n_1757),
.B2(n_1774),
.Y(n_1869)
);

AO21x1_ASAP7_75t_L g1870 ( 
.A1(n_1864),
.A2(n_1812),
.B(n_1828),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1829),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1837),
.B(n_1851),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1858),
.B(n_1806),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1829),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1866),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1842),
.A2(n_1757),
.B(n_1756),
.Y(n_1876)
);

INVx4_ASAP7_75t_L g1877 ( 
.A(n_1854),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1836),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1833),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1854),
.Y(n_1880)
);

BUFx2_ASAP7_75t_L g1881 ( 
.A(n_1851),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1848),
.B(n_1818),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1866),
.Y(n_1883)
);

INVx4_ASAP7_75t_SL g1884 ( 
.A(n_1847),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1840),
.B(n_1823),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1851),
.B(n_1797),
.Y(n_1886)
);

INVxp67_ASAP7_75t_SL g1887 ( 
.A(n_1865),
.Y(n_1887)
);

INVx2_ASAP7_75t_SL g1888 ( 
.A(n_1867),
.Y(n_1888)
);

INVx3_ASAP7_75t_L g1889 ( 
.A(n_1851),
.Y(n_1889)
);

NAND3xp33_ASAP7_75t_SL g1890 ( 
.A(n_1831),
.B(n_1818),
.C(n_1823),
.Y(n_1890)
);

AND2x6_ASAP7_75t_SL g1891 ( 
.A(n_1830),
.B(n_1781),
.Y(n_1891)
);

OR2x6_ASAP7_75t_L g1892 ( 
.A(n_1863),
.B(n_1820),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1863),
.B(n_1797),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1855),
.B(n_1820),
.Y(n_1894)
);

OAI21xp33_ASAP7_75t_L g1895 ( 
.A1(n_1834),
.A2(n_1821),
.B(n_1819),
.Y(n_1895)
);

HB1xp67_ASAP7_75t_L g1896 ( 
.A(n_1860),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1861),
.B(n_1820),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1843),
.B(n_1784),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1861),
.B(n_1811),
.Y(n_1899)
);

BUFx3_ASAP7_75t_L g1900 ( 
.A(n_1863),
.Y(n_1900)
);

INVx2_ASAP7_75t_SL g1901 ( 
.A(n_1862),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1835),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1881),
.B(n_1859),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1881),
.B(n_1859),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1871),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1884),
.B(n_1844),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1900),
.B(n_1819),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1884),
.B(n_1838),
.Y(n_1908)
);

INVx1_ASAP7_75t_SL g1909 ( 
.A(n_1880),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1898),
.B(n_1856),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1899),
.B(n_1832),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1872),
.B(n_1849),
.Y(n_1912)
);

INVx1_ASAP7_75t_SL g1913 ( 
.A(n_1880),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1875),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1899),
.B(n_1835),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1871),
.Y(n_1916)
);

INVx3_ASAP7_75t_L g1917 ( 
.A(n_1892),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1874),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1902),
.B(n_1852),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1872),
.B(n_1886),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1874),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1878),
.Y(n_1922)
);

NOR2x1p5_ASAP7_75t_L g1923 ( 
.A(n_1890),
.B(n_1849),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1878),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1902),
.B(n_1852),
.Y(n_1925)
);

BUFx2_ASAP7_75t_L g1926 ( 
.A(n_1891),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1873),
.B(n_1857),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1875),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1873),
.B(n_1868),
.Y(n_1929)
);

NOR2x1_ASAP7_75t_L g1930 ( 
.A(n_1894),
.B(n_1853),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1885),
.B(n_1895),
.Y(n_1931)
);

NAND3xp33_ASAP7_75t_L g1932 ( 
.A(n_1895),
.B(n_1876),
.C(n_1839),
.Y(n_1932)
);

NAND3xp33_ASAP7_75t_L g1933 ( 
.A(n_1876),
.B(n_1846),
.C(n_1845),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1893),
.B(n_1841),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1883),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1883),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1897),
.B(n_1868),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1888),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1877),
.B(n_1801),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1877),
.B(n_1801),
.Y(n_1940)
);

AOI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1884),
.A2(n_1850),
.B1(n_1803),
.B2(n_1821),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1883),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1905),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_1926),
.Y(n_1944)
);

NOR2xp67_ASAP7_75t_SL g1945 ( 
.A(n_1926),
.B(n_1880),
.Y(n_1945)
);

OAI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1932),
.A2(n_1930),
.B(n_1906),
.Y(n_1946)
);

AND2x2_ASAP7_75t_SL g1947 ( 
.A(n_1941),
.B(n_1877),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1923),
.B(n_1884),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1905),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1916),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1920),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1915),
.B(n_1896),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1909),
.B(n_1877),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1915),
.B(n_1896),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1938),
.Y(n_1955)
);

NAND2x2_ASAP7_75t_L g1956 ( 
.A(n_1923),
.B(n_1884),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1916),
.Y(n_1957)
);

INVx1_ASAP7_75t_SL g1958 ( 
.A(n_1913),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1918),
.Y(n_1959)
);

INVx2_ASAP7_75t_SL g1960 ( 
.A(n_1920),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1914),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1910),
.B(n_1891),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1918),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1914),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1903),
.B(n_1901),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1927),
.B(n_1911),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1931),
.B(n_1879),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1921),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1903),
.B(n_1904),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1914),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1929),
.B(n_1887),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1921),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1930),
.B(n_1932),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1938),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1922),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1922),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1928),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1928),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1924),
.Y(n_1979)
);

OAI21xp33_ASAP7_75t_L g1980 ( 
.A1(n_1933),
.A2(n_1890),
.B(n_1869),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1929),
.B(n_1887),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1924),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1904),
.B(n_1901),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1948),
.B(n_1907),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1960),
.B(n_1917),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1948),
.B(n_1969),
.Y(n_1986)
);

XNOR2xp5_ASAP7_75t_L g1987 ( 
.A(n_1973),
.B(n_1946),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1944),
.B(n_1919),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_1958),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1943),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1969),
.B(n_1965),
.Y(n_1991)
);

BUFx3_ASAP7_75t_L g1992 ( 
.A(n_1953),
.Y(n_1992)
);

INVx1_ASAP7_75t_SL g1993 ( 
.A(n_1955),
.Y(n_1993)
);

INVx2_ASAP7_75t_SL g1994 ( 
.A(n_1965),
.Y(n_1994)
);

INVx1_ASAP7_75t_SL g1995 ( 
.A(n_1974),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1960),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1966),
.B(n_1967),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1983),
.B(n_1907),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1983),
.B(n_1907),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1947),
.B(n_1907),
.Y(n_2000)
);

NAND3xp33_ASAP7_75t_L g2001 ( 
.A(n_1945),
.B(n_1933),
.C(n_1908),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1947),
.B(n_1945),
.Y(n_2002)
);

INVx1_ASAP7_75t_SL g2003 ( 
.A(n_1971),
.Y(n_2003)
);

AOI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1980),
.A2(n_1941),
.B1(n_1803),
.B2(n_1870),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1951),
.B(n_1912),
.Y(n_2005)
);

INVxp67_ASAP7_75t_L g2006 ( 
.A(n_1975),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1943),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1951),
.Y(n_2008)
);

INVx5_ASAP7_75t_L g2009 ( 
.A(n_1961),
.Y(n_2009)
);

INVx1_ASAP7_75t_SL g2010 ( 
.A(n_1971),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1981),
.Y(n_2011)
);

AOI22xp5_ASAP7_75t_L g2012 ( 
.A1(n_1956),
.A2(n_1803),
.B1(n_1870),
.B2(n_1882),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1961),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_2011),
.Y(n_2014)
);

INVx1_ASAP7_75t_SL g2015 ( 
.A(n_1989),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_2001),
.A2(n_1956),
.B1(n_1962),
.B2(n_1917),
.Y(n_2016)
);

AOI211xp5_ASAP7_75t_L g2017 ( 
.A1(n_2001),
.A2(n_1981),
.B(n_1917),
.C(n_1954),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2003),
.B(n_1975),
.Y(n_2018)
);

OAI21xp33_ASAP7_75t_SL g2019 ( 
.A1(n_2002),
.A2(n_1954),
.B(n_1952),
.Y(n_2019)
);

O2A1O1Ixp33_ASAP7_75t_L g2020 ( 
.A1(n_1989),
.A2(n_1952),
.B(n_1979),
.C(n_1982),
.Y(n_2020)
);

O2A1O1Ixp33_ASAP7_75t_L g2021 ( 
.A1(n_2002),
.A2(n_1982),
.B(n_1979),
.C(n_1976),
.Y(n_2021)
);

NAND2x1_ASAP7_75t_L g2022 ( 
.A(n_2000),
.B(n_1917),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1998),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1991),
.B(n_1912),
.Y(n_2024)
);

AOI222xp33_ASAP7_75t_L g2025 ( 
.A1(n_1987),
.A2(n_1976),
.B1(n_1950),
.B2(n_1949),
.C1(n_1972),
.C2(n_1959),
.Y(n_2025)
);

OAI211xp5_ASAP7_75t_L g2026 ( 
.A1(n_2004),
.A2(n_1949),
.B(n_1957),
.C(n_1972),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1990),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1998),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1999),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1985),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1990),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1985),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_1988),
.B(n_1925),
.Y(n_2033)
);

OAI22xp33_ASAP7_75t_SL g2034 ( 
.A1(n_2004),
.A2(n_2003),
.B1(n_2010),
.B2(n_1994),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_1988),
.B(n_1937),
.Y(n_2035)
);

OAI32xp33_ASAP7_75t_L g2036 ( 
.A1(n_1993),
.A2(n_1937),
.A3(n_1889),
.B1(n_1939),
.B2(n_1940),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2015),
.Y(n_2037)
);

AOI22xp33_ASAP7_75t_L g2038 ( 
.A1(n_2025),
.A2(n_1987),
.B1(n_1991),
.B2(n_2000),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_2034),
.A2(n_1986),
.B1(n_1992),
.B2(n_1997),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_2030),
.B(n_1986),
.Y(n_2040)
);

INVxp67_ASAP7_75t_L g2041 ( 
.A(n_2030),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_2017),
.A2(n_1984),
.B1(n_1994),
.B2(n_2005),
.Y(n_2042)
);

AOI31xp33_ASAP7_75t_L g2043 ( 
.A1(n_2019),
.A2(n_2010),
.A3(n_1993),
.B(n_1995),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2032),
.Y(n_2044)
);

NOR2xp67_ASAP7_75t_SL g2045 ( 
.A(n_2014),
.B(n_1992),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_2024),
.B(n_1984),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2023),
.B(n_1992),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2032),
.Y(n_2048)
);

INVxp67_ASAP7_75t_SL g2049 ( 
.A(n_2020),
.Y(n_2049)
);

INVx1_ASAP7_75t_SL g2050 ( 
.A(n_2035),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_2028),
.B(n_1995),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2029),
.B(n_1996),
.Y(n_2052)
);

AOI221xp5_ASAP7_75t_L g2053 ( 
.A1(n_2043),
.A2(n_2020),
.B1(n_2036),
.B2(n_2021),
.C(n_2016),
.Y(n_2053)
);

AOI211x1_ASAP7_75t_L g2054 ( 
.A1(n_2045),
.A2(n_2026),
.B(n_1997),
.C(n_2018),
.Y(n_2054)
);

AOI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_2049),
.A2(n_2021),
.B(n_2022),
.Y(n_2055)
);

AOI211xp5_ASAP7_75t_SL g2056 ( 
.A1(n_2049),
.A2(n_2026),
.B(n_2018),
.C(n_2012),
.Y(n_2056)
);

AOI21xp33_ASAP7_75t_L g2057 ( 
.A1(n_2050),
.A2(n_2033),
.B(n_1996),
.Y(n_2057)
);

AOI21xp33_ASAP7_75t_SL g2058 ( 
.A1(n_2037),
.A2(n_1996),
.B(n_2012),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_2038),
.A2(n_2006),
.B(n_2008),
.Y(n_2059)
);

NAND3xp33_ASAP7_75t_L g2060 ( 
.A(n_2039),
.B(n_2008),
.C(n_2027),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_SL g2061 ( 
.A(n_2042),
.B(n_1985),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_2040),
.B(n_1985),
.Y(n_2062)
);

OAI211xp5_ASAP7_75t_L g2063 ( 
.A1(n_2047),
.A2(n_2051),
.B(n_2052),
.C(n_2041),
.Y(n_2063)
);

AOI211xp5_ASAP7_75t_L g2064 ( 
.A1(n_2040),
.A2(n_2006),
.B(n_2031),
.C(n_2008),
.Y(n_2064)
);

A2O1A1Ixp33_ASAP7_75t_L g2065 ( 
.A1(n_2046),
.A2(n_2005),
.B(n_1999),
.C(n_2007),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_L g2066 ( 
.A(n_2063),
.B(n_2041),
.Y(n_2066)
);

CKINVDCx20_ASAP7_75t_R g2067 ( 
.A(n_2061),
.Y(n_2067)
);

OAI21xp5_ASAP7_75t_SL g2068 ( 
.A1(n_2053),
.A2(n_2056),
.B(n_2059),
.Y(n_2068)
);

AOI211xp5_ASAP7_75t_L g2069 ( 
.A1(n_2057),
.A2(n_2044),
.B(n_2048),
.C(n_2007),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_2055),
.A2(n_2013),
.B(n_2009),
.Y(n_2070)
);

AND4x1_ASAP7_75t_L g2071 ( 
.A(n_2060),
.B(n_1957),
.C(n_1950),
.D(n_1959),
.Y(n_2071)
);

OAI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_2062),
.A2(n_2065),
.B(n_2058),
.Y(n_2072)
);

O2A1O1Ixp33_ASAP7_75t_L g2073 ( 
.A1(n_2064),
.A2(n_2013),
.B(n_1968),
.C(n_1963),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2071),
.Y(n_2074)
);

OAI21xp5_ASAP7_75t_L g2075 ( 
.A1(n_2068),
.A2(n_2054),
.B(n_2013),
.Y(n_2075)
);

INVx3_ASAP7_75t_L g2076 ( 
.A(n_2070),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2066),
.Y(n_2077)
);

NOR2x1_ASAP7_75t_L g2078 ( 
.A(n_2067),
.B(n_1963),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2072),
.B(n_1934),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2073),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_2069),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_2081),
.A2(n_2009),
.B1(n_1968),
.B2(n_1977),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2078),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2074),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_2081),
.A2(n_2009),
.B1(n_1889),
.B2(n_1888),
.Y(n_2085)
);

CKINVDCx20_ASAP7_75t_R g2086 ( 
.A(n_2079),
.Y(n_2086)
);

BUFx3_ASAP7_75t_L g2087 ( 
.A(n_2076),
.Y(n_2087)
);

NAND2x1p5_ASAP7_75t_L g2088 ( 
.A(n_2087),
.B(n_2076),
.Y(n_2088)
);

NAND3x1_ASAP7_75t_L g2089 ( 
.A(n_2083),
.B(n_2075),
.C(n_2077),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2086),
.Y(n_2090)
);

NOR3xp33_ASAP7_75t_L g2091 ( 
.A(n_2090),
.B(n_2076),
.C(n_2084),
.Y(n_2091)
);

OAI322xp33_ASAP7_75t_L g2092 ( 
.A1(n_2091),
.A2(n_2080),
.A3(n_2088),
.B1(n_2085),
.B2(n_2089),
.C1(n_2082),
.C2(n_1970),
.Y(n_2092)
);

OAI21xp5_ASAP7_75t_L g2093 ( 
.A1(n_2092),
.A2(n_2082),
.B(n_2009),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_2092),
.Y(n_2094)
);

INVx1_ASAP7_75t_SL g2095 ( 
.A(n_2094),
.Y(n_2095)
);

OAI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_2093),
.A2(n_2009),
.B(n_1970),
.Y(n_2096)
);

HB1xp67_ASAP7_75t_L g2097 ( 
.A(n_2096),
.Y(n_2097)
);

BUFx2_ASAP7_75t_L g2098 ( 
.A(n_2095),
.Y(n_2098)
);

HB1xp67_ASAP7_75t_L g2099 ( 
.A(n_2098),
.Y(n_2099)
);

AOI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_2099),
.A2(n_2097),
.B(n_2009),
.Y(n_2100)
);

AOI21xp5_ASAP7_75t_L g2101 ( 
.A1(n_2100),
.A2(n_2009),
.B(n_1977),
.Y(n_2101)
);

OAI21xp5_ASAP7_75t_L g2102 ( 
.A1(n_2101),
.A2(n_1978),
.B(n_1964),
.Y(n_2102)
);

AOI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_2102),
.A2(n_1978),
.B1(n_1964),
.B2(n_1942),
.Y(n_2103)
);

AOI211xp5_ASAP7_75t_L g2104 ( 
.A1(n_2103),
.A2(n_1942),
.B(n_1936),
.C(n_1935),
.Y(n_2104)
);


endmodule