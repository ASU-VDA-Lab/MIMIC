module fake_jpeg_7034_n_281 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_36),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_24),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_39),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_0),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_44),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_48),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_27),
.B(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_50),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_14),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_13),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_29),
.B(n_23),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_28),
.B1(n_19),
.B2(n_31),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_52),
.A2(n_88),
.B1(n_22),
.B2(n_21),
.Y(n_112)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_53),
.B(n_64),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVxp67_ASAP7_75t_SL g107 ( 
.A(n_57),
.Y(n_107)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_61),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_62),
.Y(n_115)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_66),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_43),
.A2(n_28),
.B1(n_19),
.B2(n_31),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_69),
.A2(n_80),
.B(n_21),
.C(n_13),
.Y(n_124)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_71),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_74),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_34),
.C(n_24),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_51),
.C(n_48),
.Y(n_109)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_81),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_26),
.B1(n_32),
.B2(n_22),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_22),
.B1(n_32),
.B2(n_26),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_85),
.Y(n_117)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_84),
.B1(n_12),
.B2(n_11),
.Y(n_127)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_113)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_39),
.A2(n_27),
.B1(n_33),
.B2(n_20),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_43),
.A2(n_33),
.B1(n_29),
.B2(n_23),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_54),
.B1(n_76),
.B2(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_37),
.B(n_34),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_98),
.Y(n_114)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_49),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_49),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_97),
.Y(n_104)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_30),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_43),
.B1(n_30),
.B2(n_22),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_101),
.A2(n_105),
.B1(n_116),
.B2(n_78),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_43),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_106),
.C(n_89),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_109),
.Y(n_158)
);

AOI22x1_ASAP7_75t_L g105 ( 
.A1(n_61),
.A2(n_49),
.B1(n_26),
.B2(n_32),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_92),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_108),
.A2(n_119),
.B1(n_1),
.B2(n_2),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_112),
.B(n_124),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_21),
.B1(n_32),
.B2(n_9),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_65),
.A2(n_12),
.A3(n_11),
.B1(n_10),
.B2(n_4),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_55),
.B(n_96),
.C(n_64),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_70),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_133),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_60),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_131),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_117),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_126),
.B(n_110),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_73),
.B(n_94),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_104),
.B(n_110),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_151),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_138),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_56),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_139),
.B(n_145),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_84),
.B1(n_73),
.B2(n_78),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_140),
.A2(n_160),
.B1(n_144),
.B2(n_153),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_154),
.B1(n_108),
.B2(n_100),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_147),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_57),
.B1(n_86),
.B2(n_56),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_115),
.B1(n_125),
.B2(n_120),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_68),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_149),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_118),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_150),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_68),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_1),
.Y(n_152)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_53),
.B1(n_95),
.B2(n_62),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_1),
.Y(n_157)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_104),
.B(n_1),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_132),
.B(n_158),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_165),
.B(n_154),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_185),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_100),
.B1(n_102),
.B2(n_115),
.Y(n_170)
);

HAxp5_ASAP7_75t_SL g172 ( 
.A(n_159),
.B(n_62),
.CON(n_172),
.SN(n_172)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_172),
.A2(n_133),
.B(n_136),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_120),
.B1(n_3),
.B2(n_4),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_135),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_95),
.C(n_125),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_191),
.C(n_152),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_148),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_155),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_189),
.B1(n_149),
.B2(n_128),
.Y(n_201)
);

A2O1A1O1Ixp25_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_137),
.B(n_132),
.C(n_139),
.D(n_145),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_134),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_131),
.B(n_7),
.C(n_3),
.Y(n_191)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_181),
.B(n_138),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_199),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_178),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_158),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_210),
.B(n_212),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_130),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_206),
.C(n_211),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_213),
.B1(n_176),
.B2(n_173),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_181),
.B(n_147),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_205),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_143),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

AOI221xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_157),
.B1(n_184),
.B2(n_174),
.C(n_7),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_158),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_183),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_142),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_146),
.B(n_142),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_166),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_165),
.B1(n_171),
.B2(n_180),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_214),
.A2(n_224),
.B1(n_201),
.B2(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_200),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_190),
.C(n_167),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_223),
.C(n_228),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_231),
.B1(n_202),
.B2(n_195),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_208),
.B(n_162),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_208),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_167),
.C(n_191),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_180),
.B1(n_186),
.B2(n_169),
.Y(n_224)
);

OAI322xp33_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_168),
.A3(n_179),
.B1(n_163),
.B2(n_166),
.C1(n_175),
.C2(n_172),
.Y(n_226)
);

NOR3xp33_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_199),
.C(n_196),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_170),
.C(n_160),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_192),
.A2(n_163),
.B1(n_140),
.B2(n_129),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_210),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_234),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_225),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_237),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_239),
.C(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_227),
.B(n_213),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_198),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_242),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_224),
.B1(n_221),
.B2(n_222),
.Y(n_240)
);

AOI322xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_218),
.A3(n_231),
.B1(n_233),
.B2(n_239),
.C1(n_242),
.C2(n_235),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_220),
.A2(n_221),
.B1(n_228),
.B2(n_217),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_215),
.C(n_223),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_203),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_245),
.A2(n_227),
.B(n_219),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_255),
.B(n_230),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_245),
.A2(n_220),
.B(n_222),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_184),
.B(n_174),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_254),
.C(n_241),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_216),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_207),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_229),
.C(n_204),
.Y(n_254)
);

OAI31xp33_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_236),
.A3(n_244),
.B(n_243),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_257),
.B(n_259),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_229),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_262),
.B(n_263),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_264),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_248),
.A2(n_197),
.B1(n_230),
.B2(n_143),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_261),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_6),
.B(n_2),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_2),
.C(n_5),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_259),
.B(n_250),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_260),
.Y(n_272)
);

INVxp33_ASAP7_75t_SL g270 ( 
.A(n_261),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

AOI31xp33_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_250),
.A3(n_253),
.B(n_5),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_258),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_273),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_264),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_268),
.C(n_270),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_275),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_278),
.A2(n_267),
.B(n_265),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_280),
.Y(n_281)
);


endmodule