module real_jpeg_5720_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_0),
.A2(n_48),
.B1(n_51),
.B2(n_54),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_0),
.A2(n_54),
.B1(n_202),
.B2(n_306),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_0),
.A2(n_54),
.B1(n_157),
.B2(n_158),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_0),
.A2(n_54),
.B1(n_325),
.B2(n_390),
.Y(n_389)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_1),
.Y(n_189)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_1),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_1),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g410 ( 
.A(n_1),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_2),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g346 ( 
.A(n_2),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_2),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_2),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_2),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_3),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_3),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_97),
.B1(n_126),
.B2(n_130),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_3),
.A2(n_58),
.B1(n_97),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_3),
.A2(n_97),
.B1(n_199),
.B2(n_374),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_4),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_4),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_4),
.A2(n_276),
.B1(n_354),
.B2(n_357),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_4),
.A2(n_276),
.B1(n_385),
.B2(n_388),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_L g440 ( 
.A1(n_4),
.A2(n_134),
.B1(n_276),
.B2(n_441),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_5),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_5),
.A2(n_60),
.B1(n_216),
.B2(n_224),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_5),
.A2(n_60),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_5),
.A2(n_60),
.B1(n_425),
.B2(n_426),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_6),
.A2(n_85),
.B1(n_87),
.B2(n_91),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_6),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_6),
.A2(n_51),
.B1(n_91),
.B2(n_133),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_6),
.A2(n_91),
.B1(n_275),
.B2(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_6),
.A2(n_91),
.B1(n_357),
.B2(n_400),
.Y(n_399)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_7),
.Y(n_323)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_8),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_9),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_9),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_9),
.A2(n_163),
.B1(n_198),
.B2(n_202),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_9),
.A2(n_163),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_9),
.A2(n_163),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_10),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_10),
.Y(n_172)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_12),
.Y(n_120)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_12),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_12),
.Y(n_192)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_14),
.Y(n_520)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_15),
.A2(n_178),
.B1(n_182),
.B2(n_183),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_15),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_15),
.A2(n_182),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_15),
.A2(n_182),
.B1(n_265),
.B2(n_351),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_15),
.A2(n_182),
.B1(n_393),
.B2(n_395),
.Y(n_392)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_17),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_17),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_17),
.B(n_172),
.C(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_17),
.B(n_72),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_17),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_17),
.B(n_166),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_17),
.B(n_260),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_18),
.A2(n_77),
.B1(n_157),
.B2(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_18),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_18),
.A2(n_208),
.B1(n_223),
.B2(n_228),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_18),
.A2(n_45),
.B1(n_208),
.B2(n_267),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_18),
.A2(n_31),
.B1(n_32),
.B2(n_208),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_516),
.B(n_518),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_146),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_144),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_141),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_23),
.B(n_141),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_131),
.C(n_138),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_24),
.A2(n_25),
.B1(n_512),
.B2(n_513),
.Y(n_511)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_61),
.C(n_98),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_26),
.B(n_504),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_47),
.B1(n_55),
.B2(n_57),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_27),
.A2(n_55),
.B1(n_57),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_27),
.A2(n_55),
.B1(n_132),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_27),
.A2(n_344),
.B(n_392),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_27),
.A2(n_38),
.B1(n_392),
.B2(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_27),
.A2(n_47),
.B1(n_55),
.B2(n_489),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_28),
.A2(n_341),
.B(n_343),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_28),
.B(n_345),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_38),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_33),
.Y(n_320)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_38),
.B(n_159),
.Y(n_303)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_40),
.Y(n_257)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_41),
.Y(n_425)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_43),
.Y(n_387)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_43),
.Y(n_428)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g342 ( 
.A(n_50),
.Y(n_342)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_55),
.A2(n_413),
.B(n_443),
.Y(n_453)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_56),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_56),
.B(n_440),
.Y(n_439)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_61),
.A2(n_98),
.B1(n_99),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_61),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_84),
.B1(n_92),
.B2(n_93),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_62),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_62),
.A2(n_92),
.B1(n_299),
.B2(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_62),
.A2(n_92),
.B1(n_384),
.B2(n_389),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_62),
.A2(n_84),
.B1(n_92),
.B2(n_493),
.Y(n_492)
);

OR2x2_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_72),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_63)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_64),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_71),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_71),
.Y(n_328)
);

BUFx5_ASAP7_75t_L g351 ( 
.A(n_71),
.Y(n_351)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_72),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

AOI22x1_ASAP7_75t_L g414 ( 
.A1(n_72),
.A2(n_139),
.B1(n_301),
.B2(n_415),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_72),
.A2(n_139),
.B1(n_423),
.B2(n_424),
.Y(n_422)
);

AO22x2_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_79),
.B2(n_81),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_75),
.Y(n_286)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g287 ( 
.A(n_77),
.B(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_77),
.Y(n_379)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_78),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_80),
.Y(n_356)
);

INVx6_ASAP7_75t_L g359 ( 
.A(n_80),
.Y(n_359)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_86),
.Y(n_266)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_90),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_92),
.B(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_92),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_94),
.Y(n_390)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_98),
.A2(n_99),
.B1(n_491),
.B2(n_492),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_98),
.B(n_488),
.C(n_491),
.Y(n_499)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_116),
.B(n_125),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_100),
.A2(n_156),
.B(n_160),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_100),
.A2(n_116),
.B1(n_207),
.B2(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_100),
.A2(n_160),
.B(n_250),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_100),
.A2(n_116),
.B1(n_353),
.B2(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_101),
.B(n_161),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_101),
.A2(n_166),
.B1(n_377),
.B2(n_378),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_101),
.A2(n_166),
.B1(n_378),
.B2(n_399),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_101),
.A2(n_166),
.B1(n_399),
.B2(n_431),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_116),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B1(n_109),
.B2(n_113),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx5_ASAP7_75t_SL g285 ( 
.A(n_113),
.Y(n_285)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_116),
.A2(n_207),
.B(n_209),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_116),
.A2(n_209),
.B(n_353),
.Y(n_352)
);

AOI22x1_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_119),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_120),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_120),
.Y(n_375)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_125),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_130),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_131),
.B(n_138),
.Y(n_513)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_134),
.B(n_159),
.Y(n_329)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_139),
.A2(n_256),
.B(n_263),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_139),
.B(n_301),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_139),
.A2(n_263),
.B(n_456),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_510),
.B(n_515),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_482),
.B(n_507),
.Y(n_147)
);

OAI311xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_362),
.A3(n_458),
.B1(n_476),
.C1(n_477),
.Y(n_148)
);

AOI21x1_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_312),
.B(n_361),
.Y(n_149)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_290),
.B(n_311),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_244),
.B(n_289),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_212),
.B(n_243),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_175),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_154),
.B(n_175),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_167),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_155),
.A2(n_167),
.B1(n_168),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_155),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_159),
.A2(n_186),
.B(n_193),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_SL g256 ( 
.A1(n_159),
.A2(n_257),
.B(n_258),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_SL g341 ( 
.A1(n_159),
.A2(n_329),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_162),
.Y(n_251)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_204),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_176),
.B(n_205),
.C(n_211),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_186),
.B(n_193),
.Y(n_176)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_179),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_185),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_186),
.A2(n_195),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_186),
.A2(n_368),
.B1(n_371),
.B2(n_373),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_186),
.A2(n_195),
.B(n_373),
.Y(n_401)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_197),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_187),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_187),
.A2(n_273),
.B1(n_305),
.B2(n_308),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_187),
.A2(n_334),
.B1(n_408),
.B2(n_409),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_189),
.Y(n_309)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx8_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_192),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_222),
.B(n_231),
.Y(n_221)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_210),
.B2(n_211),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_234),
.B(n_242),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_220),
.B(n_233),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_232),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_232),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_231),
.A2(n_272),
.B(n_279),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_240),
.Y(n_242)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_246),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_270),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_254),
.B2(n_255),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_254),
.C(n_270),
.Y(n_291)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_253),
.Y(n_381)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI32xp33_ASAP7_75t_L g282 ( 
.A1(n_259),
.A2(n_283),
.A3(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_282)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_269),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_282),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_282),
.Y(n_296)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_281),
.Y(n_372)
);

INVx4_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_291),
.B(n_292),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_297),
.B2(n_310),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_296),
.C(n_310),
.Y(n_313)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_302),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_303),
.C(n_304),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_313),
.B(n_314),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_338),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.Y(n_315)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_330),
.B2(n_331),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_318),
.B(n_330),
.Y(n_454)
);

OAI32xp33_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_320),
.A3(n_321),
.B1(n_324),
.B2(n_329),
.Y(n_318)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_325),
.Y(n_324)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_326),
.Y(n_325)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_335),
.B(n_337),
.C(n_338),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_348),
.B2(n_360),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_339),
.B(n_349),
.C(n_352),
.Y(n_467)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_347),
.Y(n_395)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_348),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_352),
.Y(n_348)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_350),
.Y(n_456)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NAND2xp33_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_444),
.Y(n_362)
);

A2O1A1Ixp33_ASAP7_75t_SL g477 ( 
.A1(n_363),
.A2(n_444),
.B(n_478),
.C(n_481),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_416),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_364),
.B(n_416),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_396),
.C(n_403),
.Y(n_364)
);

FAx1_ASAP7_75t_SL g457 ( 
.A(n_365),
.B(n_396),
.CI(n_403),
.CON(n_457),
.SN(n_457)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_382),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_366),
.B(n_383),
.C(n_391),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_376),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_367),
.B(n_376),
.Y(n_450)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_368),
.Y(n_408)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_377),
.Y(n_406)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_391),
.Y(n_382)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_386),
.Y(n_385)
);

INVx6_ASAP7_75t_SL g386 ( 
.A(n_387),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_389),
.Y(n_423)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_401),
.B2(n_402),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_398),
.B(n_401),
.Y(n_435)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_401),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_401),
.A2(n_402),
.B1(n_437),
.B2(n_438),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_401),
.A2(n_435),
.B(n_438),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_411),
.C(n_414),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_404),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_407),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_405),
.B(n_407),
.Y(n_466)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_411),
.A2(n_412),
.B1(n_414),
.B2(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_414),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_417),
.B(n_420),
.C(n_433),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_419),
.A2(n_420),
.B1(n_433),
.B2(n_434),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_429),
.B(n_432),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_430),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_424),
.Y(n_493)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

FAx1_ASAP7_75t_SL g484 ( 
.A(n_432),
.B(n_485),
.CI(n_486),
.CON(n_484),
.SN(n_484)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_432),
.B(n_485),
.C(n_486),
.Y(n_506)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_443),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_440),
.Y(n_489)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_457),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_445),
.B(n_457),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_450),
.C(n_451),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_446),
.A2(n_447),
.B1(n_450),
.B2(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_450),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_451),
.B(n_469),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_454),
.C(n_455),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_452),
.A2(n_453),
.B1(n_455),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_454),
.B(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_455),
.Y(n_464)
);

BUFx24_ASAP7_75t_SL g521 ( 
.A(n_457),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_459),
.B(n_471),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_460),
.A2(n_479),
.B(n_480),
.Y(n_478)
);

NOR2x1_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_468),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_468),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_465),
.C(n_467),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_462),
.B(n_474),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_465),
.A2(n_466),
.B1(n_467),
.B2(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_467),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_472),
.B(n_473),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_496),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_484),
.B(n_495),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_495),
.Y(n_508)
);

BUFx24_ASAP7_75t_SL g523 ( 
.A(n_484),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_487),
.A2(n_488),
.B1(n_490),
.B2(n_494),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_487),
.A2(n_488),
.B1(n_502),
.B2(n_503),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_487),
.B(n_498),
.C(n_502),
.Y(n_514)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_490),
.Y(n_494)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_496),
.A2(n_508),
.B(n_509),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_506),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_506),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_499),
.B1(n_500),
.B2(n_501),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_514),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_514),
.Y(n_515)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx6_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx13_ASAP7_75t_L g519 ( 
.A(n_517),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_520),
.Y(n_518)
);


endmodule