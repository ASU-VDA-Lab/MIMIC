module fake_jpeg_29136_n_324 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx8_ASAP7_75t_SL g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_13),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_41),
.B(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_10),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_59),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_26),
.B(n_9),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_21),
.B(n_9),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_60),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_16),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_65),
.B(n_32),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_47),
.Y(n_74)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_67),
.Y(n_110)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_70),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_27),
.B1(n_33),
.B2(n_35),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_71),
.A2(n_111),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_27),
.B1(n_35),
.B2(n_33),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_76),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_20),
.B1(n_35),
.B2(n_33),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_78),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_36),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_119),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_23),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_98),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_40),
.A2(n_39),
.B1(n_38),
.B2(n_31),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_95),
.B1(n_8),
.B2(n_6),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_43),
.A2(n_39),
.B1(n_38),
.B2(n_31),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_23),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_44),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g141 ( 
.A(n_99),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_46),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_47),
.B(n_20),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_58),
.B(n_34),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_32),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_70),
.A2(n_31),
.B1(n_37),
.B2(n_29),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_106),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_37),
.C(n_29),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_7),
.C(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_0),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_116),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_48),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_111)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_50),
.B(n_2),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_61),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_100),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_29),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_120),
.A2(n_126),
.B1(n_113),
.B2(n_97),
.Y(n_178)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_122),
.A2(n_124),
.B1(n_136),
.B2(n_139),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_8),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_125),
.B(n_128),
.Y(n_167)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_82),
.B(n_7),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_158),
.C(n_86),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_146),
.B(n_86),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_75),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_140),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_87),
.A2(n_107),
.B1(n_77),
.B2(n_85),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_87),
.B(n_84),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_99),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_88),
.A2(n_83),
.B1(n_92),
.B2(n_117),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_75),
.Y(n_140)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_91),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_150),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_90),
.A2(n_108),
.B1(n_93),
.B2(n_85),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_79),
.B(n_90),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_148),
.B(n_149),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_73),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_91),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_88),
.A2(n_114),
.B1(n_92),
.B2(n_83),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_152),
.A2(n_155),
.B1(n_141),
.B2(n_131),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_96),
.A2(n_108),
.B1(n_93),
.B2(n_80),
.Y(n_153)
);

AO22x1_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_154),
.B1(n_130),
.B2(n_155),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_96),
.A2(n_80),
.B1(n_118),
.B2(n_115),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_97),
.A2(n_81),
.B1(n_110),
.B2(n_115),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_99),
.B(n_86),
.C(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_160),
.B(n_163),
.Y(n_200)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_123),
.B(n_136),
.CI(n_129),
.CON(n_162),
.SN(n_162)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_162),
.B(n_124),
.Y(n_195)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_165),
.A2(n_153),
.B(n_154),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_170),
.B(n_173),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_190),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_137),
.C(n_148),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_179),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_156),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_174),
.B(n_187),
.Y(n_225)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_81),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_184),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_192),
.B1(n_152),
.B2(n_141),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_132),
.C(n_133),
.Y(n_179)
);

NAND2xp33_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_154),
.Y(n_206)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_135),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_122),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_167),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_132),
.B(n_133),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_128),
.B(n_145),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_191),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_126),
.A2(n_131),
.B1(n_147),
.B2(n_130),
.Y(n_192)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_193),
.Y(n_201)
);

XOR2x2_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_147),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_216),
.C(n_220),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_214),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_186),
.A2(n_146),
.B1(n_153),
.B2(n_154),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_207),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_153),
.B1(n_154),
.B2(n_134),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_215),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_180),
.A2(n_190),
.B1(n_165),
.B2(n_153),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_205),
.A2(n_210),
.B1(n_214),
.B2(n_217),
.Y(n_247)
);

AO22x2_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_204),
.B1(n_197),
.B2(n_196),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_180),
.A2(n_140),
.B1(n_143),
.B2(n_150),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_141),
.B(n_159),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_218),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_159),
.A2(n_162),
.B1(n_168),
.B2(n_185),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_188),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_171),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_177),
.A2(n_173),
.B1(n_176),
.B2(n_184),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_176),
.B1(n_182),
.B2(n_164),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_182),
.A2(n_161),
.B1(n_175),
.B2(n_181),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_198),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_164),
.A2(n_193),
.B1(n_166),
.B2(n_183),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_180),
.B1(n_192),
.B2(n_178),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_230),
.B(n_232),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_195),
.B1(n_210),
.B2(n_220),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_231),
.A2(n_242),
.B1(n_201),
.B2(n_208),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_239),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_215),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_237),
.Y(n_253)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_199),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_238),
.B(n_237),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_213),
.C(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_212),
.B1(n_202),
.B2(n_194),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_225),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_249),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_213),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_194),
.B(n_207),
.C(n_201),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_239),
.Y(n_265)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_208),
.B(n_219),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_250),
.A2(n_266),
.B(n_229),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_260),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_219),
.B(n_223),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_233),
.B(n_240),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_228),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_241),
.Y(n_281)
);

OAI21x1_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_268),
.B(n_238),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_234),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_227),
.B(n_226),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_236),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_235),
.B(n_227),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_269),
.B(n_271),
.Y(n_289)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_245),
.C(n_231),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_274),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_266),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_253),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_256),
.B(n_247),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_278),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_255),
.A2(n_251),
.B1(n_259),
.B2(n_230),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_229),
.B1(n_255),
.B2(n_252),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_281),
.A2(n_258),
.B1(n_259),
.B2(n_262),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_284),
.A2(n_285),
.B1(n_288),
.B2(n_290),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_247),
.B1(n_251),
.B2(n_263),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_281),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_293),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_268),
.B1(n_230),
.B2(n_250),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_274),
.A2(n_230),
.B1(n_258),
.B2(n_250),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_253),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_295),
.B(n_257),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_299),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_271),
.C(n_269),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_293),
.C(n_254),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_294),
.A2(n_260),
.B1(n_230),
.B2(n_282),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_300),
.A2(n_305),
.B1(n_285),
.B2(n_290),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_257),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_303),
.Y(n_313)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_280),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_306),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_282),
.B1(n_272),
.B2(n_278),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_279),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_309),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_301),
.A2(n_288),
.B(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_310),
.B(n_312),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_SL g312 ( 
.A(n_300),
.B(n_298),
.C(n_296),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_302),
.C(n_296),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_302),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_305),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

NOR3xp33_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_308),
.C(n_313),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_319),
.B(n_314),
.C(n_312),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_320),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_309),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_246),
.Y(n_324)
);


endmodule