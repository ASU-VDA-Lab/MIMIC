module real_jpeg_28867_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g48 ( 
.A(n_0),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_1),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_4),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_7),
.A2(n_10),
.B(n_47),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_8),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_8),
.A2(n_27),
.B1(n_46),
.B2(n_47),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_8),
.A2(n_27),
.B1(n_38),
.B2(n_39),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_30),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_10),
.A2(n_20),
.B1(n_21),
.B2(n_30),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_10),
.A2(n_20),
.B(n_23),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_10),
.A2(n_30),
.B1(n_46),
.B2(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_10),
.B(n_19),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_SL g117 ( 
.A1(n_10),
.A2(n_39),
.B(n_59),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_10),
.B(n_52),
.Y(n_142)
);

HAxp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_111),
.CON(n_11),
.SN(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_109),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_85),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_15),
.B(n_85),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_63),
.C(n_75),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_16),
.B(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_33),
.B1(n_61),
.B2(n_62),
.Y(n_16)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_17),
.B(n_34),
.C(n_50),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_24),
.B(n_28),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_19),
.A2(n_29),
.B1(n_31),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_20),
.A2(n_21),
.B1(n_53),
.B2(n_59),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_20),
.A2(n_30),
.B(n_60),
.C(n_117),
.Y(n_116)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_22),
.A2(n_26),
.B(n_30),
.C(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_30),
.A2(n_39),
.B(n_44),
.C(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_30),
.B(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_30),
.B(n_45),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_33),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_40),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_37),
.B(n_41),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_37),
.A2(n_41),
.B1(n_45),
.B2(n_101),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_46),
.B(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_71),
.Y(n_70)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_49),
.B(n_99),
.C(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_49),
.A2(n_50),
.B1(n_98),
.B2(n_99),
.Y(n_163)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_54),
.B(n_55),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_54),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_63),
.B(n_75),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_68),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_67),
.A2(n_68),
.B1(n_141),
.B2(n_144),
.Y(n_140)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_68),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_68),
.B(n_156),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_68),
.B(n_131),
.C(n_143),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_74),
.B(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_70),
.B(n_71),
.Y(n_120)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.C(n_83),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_76),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_76),
.A2(n_91),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_79),
.A2(n_83),
.B1(n_84),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_79),
.B(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_80),
.A2(n_106),
.B(n_108),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_93),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_104),
.B2(n_105),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_98),
.A2(n_99),
.B1(n_138),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_99),
.B(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_102),
.B(n_103),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_166),
.B(n_170),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_134),
.B(n_165),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_122),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_122),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_121),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_128),
.B2(n_129),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_131),
.C(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_125),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_126),
.B(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_130),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_133),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_160),
.B(n_164),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_145),
.B(n_159),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_140),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_138),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_141),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_149),
.B(n_158),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_155),
.B(n_157),
.Y(n_149)
);

INVx5_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_162),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_168),
.Y(n_170)
);


endmodule