module real_jpeg_31871_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_0),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_0),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_495),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_1),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_2),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_2),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_3),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_3),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_3),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_3),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_3),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_3),
.B(n_344),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_3),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_3),
.B(n_398),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_4),
.Y(n_342)
);

NAND2x1_ASAP7_75t_SL g39 ( 
.A(n_5),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_5),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_5),
.B(n_108),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_5),
.B(n_97),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_5),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_5),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_5),
.B(n_457),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_6),
.Y(n_82)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_6),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_6),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_7),
.B(n_55),
.Y(n_54)
);

NAND2xp67_ASAP7_75t_SL g74 ( 
.A(n_7),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_7),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_7),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_7),
.B(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_7),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_7),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_7),
.B(n_367),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_8),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_8),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_8),
.B(n_30),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_8),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_8),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_8),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_8),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g245 ( 
.A(n_8),
.B(n_128),
.Y(n_245)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_9),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_9),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_10),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_10),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_10),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_10),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_10),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_10),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_10),
.B(n_407),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_12),
.Y(n_381)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_13),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_13),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_14),
.B(n_30),
.Y(n_63)
);

NAND2x1_ASAP7_75t_L g73 ( 
.A(n_14),
.B(n_50),
.Y(n_73)
);

NAND2x1p5_ASAP7_75t_L g88 ( 
.A(n_14),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_14),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_14),
.B(n_159),
.Y(n_158)
);

BUFx24_ASAP7_75t_L g164 ( 
.A(n_14),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_15),
.B(n_30),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_15),
.B(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_15),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_15),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_15),
.B(n_463),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_16),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_17),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_17),
.B(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_17),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_17),
.B(n_333),
.Y(n_332)
);

AND2x2_ASAP7_75t_SL g378 ( 
.A(n_17),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_17),
.B(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_17),
.B(n_412),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_450),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OA21x2_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_325),
.B(n_442),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_265),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_23),
.A2(n_443),
.B(n_446),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_180),
.B1(n_224),
.B2(n_264),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_25),
.B(n_181),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_112),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_26),
.B(n_113),
.C(n_178),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_46),
.C(n_69),
.Y(n_26)
);

XOR2x1_ASAP7_75t_L g184 ( 
.A(n_27),
.B(n_47),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_35),
.C(n_39),
.Y(n_27)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_28),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

OA21x2_ASAP7_75t_L g270 ( 
.A1(n_29),
.A2(n_31),
.B(n_218),
.Y(n_270)
);

INVx4_ASAP7_75t_SL g350 ( 
.A(n_30),
.Y(n_350)
);

INVx8_ASAP7_75t_L g413 ( 
.A(n_30),
.Y(n_413)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_34),
.Y(n_177)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_34),
.Y(n_195)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_34),
.Y(n_240)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_34),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_35),
.B(n_39),
.Y(n_217)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_43),
.Y(n_404)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_45),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_45),
.Y(n_209)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_45),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_57),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_49),
.Y(n_56)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_51),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_53),
.B(n_56),
.C(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.C(n_64),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_58),
.B(n_62),
.C(n_64),
.Y(n_169)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_59),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_59),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_61),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_61),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_212)
);

AO22x1_ASAP7_75t_SL g371 ( 
.A1(n_62),
.A2(n_63),
.B1(n_135),
.B2(n_230),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_63),
.B(n_229),
.Y(n_287)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVxp67_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2x1_ASAP7_75t_L g183 ( 
.A(n_70),
.B(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_83),
.C(n_98),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_71),
.B(n_83),
.Y(n_314)
);

XOR2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_73),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_73),
.A2(n_154),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_74),
.B(n_152),
.C(n_153),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_76),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_80),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.C(n_93),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_84),
.B(n_272),
.Y(n_271)
);

BUFx4f_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_87),
.B(n_94),
.Y(n_272)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2x1_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_88),
.B(n_117),
.C(n_119),
.Y(n_256)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_92),
.Y(n_369)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_98),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.C(n_107),
.Y(n_98)
);

XNOR2x1_ASAP7_75t_SL g188 ( 
.A(n_99),
.B(n_104),
.Y(n_188)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_103),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_104),
.A2(n_472),
.B1(n_473),
.B2(n_478),
.Y(n_471)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_104),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_107),
.B(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_107),
.B(n_188),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_110),
.Y(n_354)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_111),
.Y(n_396)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_111),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_146),
.B1(n_178),
.B2(n_179),
.Y(n_112)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_114),
.B(n_122),
.C(n_133),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_120),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_158),
.C(n_163),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_119),
.B(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_120),
.B(n_356),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_133),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.C(n_130),
.Y(n_122)
);

XOR2x2_ASAP7_75t_SL g148 ( 
.A(n_123),
.B(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2x1_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_130),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_134),
.A2(n_229),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_135),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_139),
.B(n_229),
.C(n_231),
.Y(n_228)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_142),
.Y(n_384)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_143),
.Y(n_231)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_145),
.Y(n_465)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_167),
.Y(n_146)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_147),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_155),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_148),
.Y(n_223)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_153),
.Y(n_482)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_161),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_156),
.A2(n_157),
.B1(n_462),
.B2(n_466),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_162),
.A2(n_163),
.B1(n_191),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_164),
.B(n_239),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g475 ( 
.A(n_164),
.B(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_170),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_171),
.B(n_173),
.C(n_175),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g467 ( 
.A(n_175),
.B(n_251),
.C(n_255),
.Y(n_467)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_176),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.C(n_219),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_183),
.B(n_220),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_185),
.B(n_324),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_210),
.C(n_215),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_186),
.B(n_317),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.C(n_196),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_189),
.A2(n_190),
.B1(n_196),
.B2(n_197),
.Y(n_309)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_191),
.Y(n_305)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.C(n_206),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_198),
.A2(n_206),
.B1(n_207),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_198),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_202),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_203),
.B(n_291),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_207),
.B1(n_243),
.B2(n_246),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_206),
.A2(n_207),
.B1(n_474),
.B2(n_475),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_206),
.B(n_229),
.C(n_245),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_210),
.A2(n_211),
.B1(n_216),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_216),
.Y(n_318)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_224),
.B(n_264),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_224),
.B(n_264),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_260),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_247),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_226),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_242),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_232),
.B1(n_233),
.B2(n_241),
.Y(n_227)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_232),
.B(n_241),
.C(n_242),
.Y(n_468)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2x2_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_235),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_235),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_238),
.Y(n_483)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

INVxp33_ASAP7_75t_SL g490 ( 
.A(n_247),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_259),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_258),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_249),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_249)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_258),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_259),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_260),
.B(n_490),
.C(n_491),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_260)
);

NOR2x1_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_319),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_310),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_267),
.B(n_310),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_288),
.C(n_306),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_268),
.B(n_440),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_273),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_270),
.B(n_271),
.C(n_273),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_281),
.C(n_287),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_274),
.A2(n_275),
.B1(n_281),
.B2(n_282),
.Y(n_431)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_287),
.B(n_431),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_289),
.B(n_307),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_293),
.C(n_303),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_290),
.B(n_433),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_293),
.A2(n_303),
.B1(n_304),
.B2(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_293),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.C(n_301),
.Y(n_293)
);

XNOR2x1_ASAP7_75t_SL g362 ( 
.A(n_294),
.B(n_301),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_SL g361 ( 
.A(n_297),
.B(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_300),
.Y(n_336)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_316),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_315),
.Y(n_311)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_321),
.C(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_316),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_319),
.A2(n_444),
.B(n_445),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_320),
.B(n_323),
.Y(n_445)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_437),
.B(n_441),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_424),
.B(n_436),
.Y(n_326)
);

OAI21x1_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_373),
.B(n_423),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_358),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_329),
.B(n_358),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_347),
.C(n_355),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_331),
.B(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_337),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_338),
.C(n_343),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_343),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_347),
.A2(n_348),
.B1(n_355),
.B2(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_352),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_349),
.B(n_352),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_355),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_363),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_360),
.B(n_361),
.C(n_363),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_372),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_366),
.B1(n_370),
.B2(n_371),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_365),
.B(n_371),
.C(n_372),
.Y(n_428)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_388),
.B(n_422),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_385),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_375),
.B(n_385),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.C(n_382),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_376),
.A2(n_377),
.B1(n_418),
.B2(n_419),
.Y(n_417)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_378),
.A2(n_382),
.B1(n_383),
.B2(n_420),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_378),
.Y(n_420)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_415),
.B(n_421),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_405),
.B(n_414),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_402),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_402),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_397),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_392),
.B(n_397),
.Y(n_416)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_SL g398 ( 
.A(n_399),
.Y(n_398)
);

INVx8_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_411),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_416),
.B(n_417),
.Y(n_421)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_435),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_435),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_432),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_428),
.B1(n_429),
.B2(n_430),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_429),
.C(n_432),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_430),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_438),
.B(n_439),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_448),
.B(n_449),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_493),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_489),
.Y(n_451)
);

NOR2x1_ASAP7_75t_L g494 ( 
.A(n_452),
.B(n_489),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_469),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_468),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_467),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_461),
.Y(n_455)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_462),
.Y(n_466)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_485),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_479),
.Y(n_470)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_475),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_484),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.C(n_483),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_487),
.C(n_488),
.Y(n_485)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_498),
.Y(n_495)
);

INVx5_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);


endmodule