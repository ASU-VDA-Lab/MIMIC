module fake_jpeg_30845_n_441 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_441);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx2_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_45),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_51),
.A2(n_23),
.B1(n_19),
.B2(n_38),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_57),
.Y(n_93)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_56),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_63),
.Y(n_97)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_11),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_11),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_71),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_33),
.B(n_11),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_80),
.Y(n_116)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_85),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_34),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_88),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_32),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_98),
.B(n_128),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_37),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_120),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_45),
.A2(n_37),
.B1(n_23),
.B2(n_26),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_119),
.A2(n_127),
.B1(n_77),
.B2(n_83),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_50),
.B(n_38),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_134),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_35),
.B1(n_34),
.B2(n_26),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_66),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_52),
.B1(n_86),
.B2(n_88),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_35),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_49),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_47),
.B(n_9),
.Y(n_134)
);

BUFx8_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_140),
.Y(n_185)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_53),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_144),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_64),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_93),
.B(n_48),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_145),
.Y(n_194)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_47),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_149),
.B(n_152),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_99),
.A2(n_68),
.B1(n_67),
.B2(n_58),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_150),
.A2(n_74),
.B1(n_72),
.B2(n_96),
.Y(n_192)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_77),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_153),
.A2(n_158),
.B1(n_168),
.B2(n_108),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_119),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_154),
.B(n_164),
.Y(n_184)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

CKINVDCx12_ASAP7_75t_R g157 ( 
.A(n_114),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_161),
.B1(n_163),
.B2(n_165),
.Y(n_179)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_169),
.Y(n_181)
);

CKINVDCx12_ASAP7_75t_R g167 ( 
.A(n_104),
.Y(n_167)
);

NOR2x1_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_104),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_62),
.B1(n_46),
.B2(n_54),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_122),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_108),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_127),
.B(n_123),
.C(n_51),
.Y(n_173)
);

A2O1A1O1Ixp25_ASAP7_75t_L g208 ( 
.A1(n_173),
.A2(n_196),
.B(n_59),
.C(n_90),
.D(n_69),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_135),
.Y(n_214)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_191),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_192),
.A2(n_150),
.B1(n_92),
.B2(n_129),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_147),
.A2(n_95),
.B(n_82),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_169),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_166),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_109),
.C(n_113),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_159),
.C(n_160),
.Y(n_207)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_171),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_207),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_187),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_210),
.Y(n_229)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_219),
.B1(n_186),
.B2(n_94),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_208),
.A2(n_180),
.B(n_190),
.Y(n_251)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_217),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_15),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_221),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_135),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_215),
.Y(n_231)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_165),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_162),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_220),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_173),
.A2(n_79),
.B1(n_73),
.B2(n_96),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_156),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_223),
.B(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_151),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_225),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_142),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_113),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_180),
.Y(n_249)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_191),
.A3(n_192),
.B1(n_175),
.B2(n_178),
.Y(n_228)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_179),
.B1(n_129),
.B2(n_89),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_232),
.A2(n_237),
.B1(n_240),
.B2(n_206),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_242),
.B1(n_244),
.B2(n_204),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_249),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_185),
.B1(n_91),
.B2(n_92),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_205),
.A2(n_91),
.B1(n_94),
.B2(n_61),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_216),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_186),
.B1(n_193),
.B2(n_137),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_193),
.B1(n_199),
.B2(n_172),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_217),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_SL g253 ( 
.A1(n_247),
.A2(n_251),
.B(n_228),
.C(n_246),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_188),
.B(n_176),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_211),
.B(n_226),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_211),
.Y(n_252)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_253),
.A2(n_255),
.B(n_257),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_227),
.B(n_213),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_254),
.B(n_256),
.Y(n_304)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_210),
.B(n_212),
.C(n_211),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_227),
.B(n_225),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_229),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_258),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_215),
.B(n_224),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_259),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_261),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_207),
.Y(n_262)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_271),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_223),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_268),
.Y(n_287)
);

XNOR2x2_ASAP7_75t_SL g266 ( 
.A(n_247),
.B(n_202),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_281),
.Y(n_283)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_221),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_201),
.Y(n_269)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_275),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_177),
.B(n_176),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_209),
.Y(n_272)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_231),
.Y(n_274)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_274),
.Y(n_307)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_204),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_277),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_247),
.A2(n_177),
.B(n_190),
.Y(n_277)
);

OA21x2_ASAP7_75t_L g279 ( 
.A1(n_247),
.A2(n_183),
.B(n_199),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_183),
.C(n_172),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_244),
.C(n_242),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_233),
.A2(n_189),
.B1(n_132),
.B2(n_182),
.Y(n_281)
);

NOR4xp25_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_239),
.C(n_248),
.D(n_249),
.Y(n_282)
);

NAND3xp33_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_266),
.C(n_272),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_248),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_285),
.B(n_286),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_236),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_228),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_279),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_299),
.C(n_308),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_258),
.B(n_231),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_302),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_259),
.B(n_244),
.C(n_232),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_265),
.B(n_230),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_242),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_305),
.B(n_270),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_233),
.C(n_230),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_256),
.B(n_240),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_237),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_284),
.B(n_304),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_323),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_325),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_291),
.A2(n_264),
.B1(n_281),
.B2(n_271),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_313),
.A2(n_295),
.B1(n_292),
.B2(n_301),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_277),
.B(n_252),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_315),
.A2(n_261),
.B(n_309),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_278),
.C(n_260),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_326),
.C(n_331),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_324),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_291),
.A2(n_264),
.B1(n_252),
.B2(n_267),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_318),
.A2(n_333),
.B1(n_293),
.B2(n_288),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_SL g320 ( 
.A(n_283),
.B(n_266),
.C(n_253),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_320),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_284),
.A2(n_257),
.B1(n_275),
.B2(n_268),
.Y(n_321)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_288),
.Y(n_322)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_322),
.Y(n_350)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_286),
.C(n_285),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_296),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_330),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_294),
.B(n_255),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_328),
.B(n_329),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_307),
.A2(n_255),
.B(n_269),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_276),
.C(n_261),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_287),
.B(n_238),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_332),
.B(n_306),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_295),
.A2(n_253),
.B1(n_279),
.B2(n_269),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_283),
.B(n_279),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_290),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_337),
.A2(n_354),
.B1(n_358),
.B2(n_161),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_308),
.C(n_299),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_347),
.C(n_326),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_287),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_348),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_309),
.C(n_305),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_335),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_316),
.B(n_306),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_351),
.B(n_355),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_353),
.A2(n_327),
.B1(n_317),
.B2(n_324),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_318),
.A2(n_292),
.B1(n_301),
.B2(n_303),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_331),
.B(n_290),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_263),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_356),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_253),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_357),
.B(n_313),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_333),
.A2(n_253),
.B1(n_235),
.B2(n_274),
.Y(n_358)
);

OAI21xp33_ASAP7_75t_L g359 ( 
.A1(n_342),
.A2(n_315),
.B(n_334),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_359),
.B(n_376),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_339),
.B(n_312),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_378),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_363),
.B(n_366),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_364),
.A2(n_372),
.B1(n_358),
.B2(n_374),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_365),
.B(n_337),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_341),
.B(n_235),
.C(n_238),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_367),
.B(n_369),
.C(n_370),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_SL g368 ( 
.A(n_352),
.B(n_347),
.C(n_349),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_368),
.A2(n_346),
.B(n_336),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_274),
.C(n_195),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_338),
.B(n_195),
.C(n_182),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_263),
.C(n_138),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_374),
.C(n_336),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_340),
.A2(n_118),
.B1(n_65),
.B2(n_101),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_146),
.C(n_141),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_136),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_345),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_350),
.B(n_18),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_373),
.Y(n_379)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_379),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_380),
.A2(n_383),
.B(n_370),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_360),
.A2(n_365),
.B(n_369),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_361),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_385),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_354),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_387),
.B(n_390),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_389),
.B(n_391),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_371),
.B(n_346),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_392),
.B(n_393),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_363),
.B(n_161),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_394),
.B(n_15),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_376),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_403),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_392),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_14),
.Y(n_415)
);

NOR2xp67_ASAP7_75t_SL g401 ( 
.A(n_381),
.B(n_359),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_401),
.B(n_14),
.Y(n_416)
);

BUFx24_ASAP7_75t_SL g403 ( 
.A(n_391),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_375),
.C(n_360),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_404),
.B(n_406),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_389),
.B(n_136),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_102),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_118),
.C(n_101),
.Y(n_406)
);

OA21x2_ASAP7_75t_SL g407 ( 
.A1(n_396),
.A2(n_381),
.B(n_386),
.Y(n_407)
);

AOI31xp33_ASAP7_75t_L g424 ( 
.A1(n_407),
.A2(n_8),
.A3(n_16),
.B(n_13),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_397),
.A2(n_386),
.B1(n_393),
.B2(n_117),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_411),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_131),
.C(n_90),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_413),
.C(n_12),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_155),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_414),
.A2(n_416),
.B(n_417),
.Y(n_422)
);

AOI322xp5_ASAP7_75t_L g423 ( 
.A1(n_415),
.A2(n_12),
.A3(n_17),
.B1(n_16),
.B2(n_13),
.C1(n_9),
.C2(n_8),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_395),
.B(n_132),
.C(n_117),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_410),
.A2(n_405),
.B(n_400),
.Y(n_418)
);

MAJx2_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_421),
.C(n_424),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_425),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_415),
.A2(n_102),
.B(n_12),
.Y(n_421)
);

OA21x2_ASAP7_75t_L g428 ( 
.A1(n_423),
.A2(n_424),
.B(n_0),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_84),
.C(n_76),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_412),
.A2(n_81),
.B1(n_56),
.B2(n_13),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_426),
.B(n_414),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_1),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_419),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_429),
.A2(n_430),
.B1(n_431),
.B2(n_1),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_0),
.C(n_1),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_432),
.B(n_7),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_433),
.B(n_434),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_435),
.B(n_427),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_436),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_437),
.B(n_6),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_439),
.A2(n_7),
.B1(n_4),
.B2(n_6),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_7),
.Y(n_441)
);


endmodule