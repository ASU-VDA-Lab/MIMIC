module fake_jpeg_13846_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_26),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_12),
.B(n_3),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_17),
.C(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_0),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_46),
.B1(n_55),
.B2(n_52),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_52),
.B1(n_56),
.B2(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_79),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_53),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_93),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_29),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_85),
.C(n_8),
.Y(n_106)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_46),
.A3(n_45),
.B1(n_58),
.B2(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_100),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_89),
.B(n_96),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_52),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_9),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_41),
.B1(n_40),
.B2(n_2),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_97),
.B1(n_98),
.B2(n_7),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_0),
.B(n_1),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_3),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_80),
.B1(n_6),
.B2(n_7),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_9),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_72),
.B(n_5),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_107),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_112),
.C(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_108),
.A2(n_115),
.B(n_119),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_84),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_39),
.C(n_28),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_10),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_14),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_15),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_16),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_123),
.B(n_130),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_125),
.Y(n_131)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_113),
.B(n_22),
.CI(n_23),
.CON(n_125),
.SN(n_125)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_104),
.C(n_116),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_123),
.B1(n_128),
.B2(n_129),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_115),
.C(n_106),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_135),
.B(n_120),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_114),
.C(n_102),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_137),
.B(n_138),
.Y(n_139)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_122),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_132),
.B(n_121),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_141),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_127),
.B(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);


endmodule