module fake_jpeg_11293_n_348 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_48),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_8),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_8),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_24),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_70)
);

NAND2x1_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_19),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_86),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_74),
.B(n_96),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_55),
.Y(n_78)
);

OAI21x1_ASAP7_75t_SL g130 ( 
.A1(n_78),
.A2(n_18),
.B(n_35),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_40),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_87),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_17),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_40),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_33),
.B(n_41),
.C(n_19),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_78),
.B(n_76),
.C(n_72),
.Y(n_123)
);

INVx11_ASAP7_75t_SL g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_93),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_38),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_41),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_104),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_57),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_58),
.A2(n_31),
.B1(n_19),
.B2(n_42),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_98),
.A2(n_115),
.B1(n_39),
.B2(n_35),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_43),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_110),
.B1(n_32),
.B2(n_42),
.Y(n_126)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_51),
.B(n_27),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_38),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_52),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_2),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_88),
.B1(n_84),
.B2(n_99),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_32),
.B1(n_37),
.B2(n_26),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_25),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_114),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_60),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_49),
.A2(n_19),
.B1(n_39),
.B2(n_42),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_37),
.B1(n_32),
.B2(n_42),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_118),
.A2(n_126),
.B1(n_144),
.B2(n_99),
.Y(n_175)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_25),
.B1(n_19),
.B2(n_37),
.Y(n_120)
);

XNOR2x1_ASAP7_75t_SL g161 ( 
.A(n_120),
.B(n_151),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_123),
.A2(n_131),
.B(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_86),
.B(n_27),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_124),
.B(n_135),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_127),
.Y(n_185)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_78),
.B1(n_113),
.B2(n_112),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_129),
.A2(n_138),
.B1(n_157),
.B2(n_97),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_130),
.A2(n_82),
.B(n_117),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_76),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_71),
.A2(n_35),
.B(n_28),
.C(n_18),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_150),
.B(n_2),
.C(n_4),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_81),
.B(n_22),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_137),
.A2(n_91),
.B1(n_100),
.B2(n_77),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_28),
.B1(n_26),
.B2(n_22),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_109),
.B(n_10),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_153),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_75),
.B(n_28),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_146),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_83),
.A2(n_18),
.B1(n_7),
.B2(n_11),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_75),
.B(n_0),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_73),
.B(n_0),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_155),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_93),
.A2(n_13),
.B(n_12),
.C(n_7),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_79),
.B(n_1),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_103),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_90),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_97),
.B1(n_100),
.B2(n_91),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_73),
.B(n_1),
.Y(n_155)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_90),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_116),
.B1(n_92),
.B2(n_84),
.Y(n_158)
);

AO21x2_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_184),
.B(n_176),
.Y(n_209)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_170),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_161),
.A2(n_155),
.B1(n_149),
.B2(n_146),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_150),
.Y(n_197)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_125),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_169),
.B(n_187),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_7),
.C(n_12),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_175),
.A2(n_177),
.B1(n_185),
.B2(n_173),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_177),
.B1(n_144),
.B2(n_132),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_116),
.A3(n_101),
.B1(n_92),
.B2(n_16),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_182),
.Y(n_199)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_184),
.Y(n_224)
);

AOI32xp33_ASAP7_75t_L g186 ( 
.A1(n_122),
.A2(n_101),
.A3(n_82),
.B1(n_16),
.B2(n_13),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_133),
.B(n_140),
.C(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_151),
.A2(n_117),
.B1(n_16),
.B2(n_4),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_130),
.B(n_148),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_125),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_190),
.B(n_193),
.Y(n_198)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_141),
.A2(n_123),
.B1(n_140),
.B2(n_121),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_192),
.A2(n_185),
.B1(n_158),
.B2(n_188),
.Y(n_227)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_197),
.A2(n_200),
.B(n_203),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_183),
.A2(n_142),
.B1(n_122),
.B2(n_120),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_204),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_179),
.B(n_124),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_205),
.B(n_225),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_143),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_207),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_183),
.A2(n_140),
.B1(n_126),
.B2(n_157),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_213),
.B1(n_224),
.B2(n_218),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_134),
.B(n_131),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_222),
.B(n_191),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_118),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_212),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_153),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

INVx6_ASAP7_75t_SL g250 ( 
.A(n_214),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_194),
.B(n_139),
.CI(n_138),
.CON(n_215),
.SN(n_215)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_216),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_162),
.B(n_121),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_214),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_165),
.B(n_121),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_223),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_161),
.B(n_132),
.C(n_158),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_171),
.C(n_167),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_158),
.A2(n_175),
.B(n_180),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_173),
.Y(n_225)
);

INVx2_ASAP7_75t_R g226 ( 
.A(n_182),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_159),
.B(n_193),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_222),
.A2(n_172),
.B1(n_174),
.B2(n_166),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_241),
.B1(n_244),
.B2(n_246),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_172),
.C(n_174),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_233),
.C(n_231),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_243),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_235),
.A2(n_233),
.B1(n_254),
.B2(n_231),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_245),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_206),
.B(n_201),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_199),
.A2(n_209),
.B1(n_213),
.B2(n_211),
.Y(n_241)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_195),
.B(n_216),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_215),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_209),
.A2(n_224),
.B1(n_220),
.B2(n_203),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_208),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_249),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_196),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_210),
.B(n_221),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_253),
.Y(n_274)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_197),
.B(n_219),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_236),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_204),
.B(n_200),
.C(n_223),
.D(n_207),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_257),
.A2(n_272),
.B(n_229),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_218),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_229),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_209),
.B1(n_226),
.B2(n_221),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_209),
.B1(n_226),
.B2(n_217),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_214),
.B1(n_217),
.B2(n_247),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_251),
.A2(n_214),
.B1(n_217),
.B2(n_247),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_252),
.B1(n_239),
.B2(n_234),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_267),
.B(n_236),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_268),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_244),
.B1(n_228),
.B2(n_246),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_273),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_235),
.A2(n_232),
.B1(n_238),
.B2(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_250),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_277),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_248),
.Y(n_277)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_276),
.Y(n_279)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_271),
.C(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_292),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_230),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_287),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_235),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_288),
.B(n_289),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_240),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_293),
.Y(n_298)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_260),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_263),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_266),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_295),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_306),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_271),
.B(n_272),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_287),
.Y(n_317)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_259),
.B1(n_261),
.B2(n_264),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_305),
.A2(n_288),
.B1(n_278),
.B2(n_279),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_256),
.C(n_273),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.C(n_310),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_269),
.C(n_265),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_281),
.A2(n_265),
.B1(n_257),
.B2(n_262),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_308),
.A2(n_283),
.B1(n_250),
.B2(n_253),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_275),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_283),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_274),
.C(n_262),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_311),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_296),
.A2(n_284),
.B(n_289),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_314),
.B(n_321),
.Y(n_328)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_315),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_316),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_305),
.A2(n_242),
.B(n_307),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_310),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_297),
.C(n_298),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_313),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_318),
.Y(n_337)
);

AO221x1_ASAP7_75t_L g329 ( 
.A1(n_312),
.A2(n_301),
.B1(n_303),
.B2(n_308),
.C(n_309),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_329),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_325),
.Y(n_331)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_331),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_322),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_336),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_327),
.A2(n_311),
.B1(n_325),
.B2(n_330),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_335),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_313),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_337),
.A2(n_324),
.B(n_317),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_341),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_340),
.B(n_332),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_342),
.A2(n_338),
.B(n_343),
.Y(n_344)
);

OAI21xp33_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_339),
.B(n_331),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_327),
.C(n_323),
.Y(n_346)
);

OAI21xp33_ASAP7_75t_SL g347 ( 
.A1(n_346),
.A2(n_320),
.B(n_319),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_298),
.Y(n_348)
);


endmodule