module fake_jpeg_17491_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_41),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_18),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_19),
.B1(n_16),
.B2(n_32),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_53),
.B1(n_23),
.B2(n_20),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_30),
.B1(n_32),
.B2(n_16),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_29),
.B1(n_28),
.B2(n_21),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_24),
.B1(n_28),
.B2(n_20),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_30),
.B1(n_32),
.B2(n_16),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_75),
.B1(n_29),
.B2(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_27),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_45),
.C(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_63),
.Y(n_87)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_22),
.C(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_66),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_30),
.B1(n_34),
.B2(n_25),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_31),
.B1(n_33),
.B2(n_22),
.Y(n_109)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_36),
.A2(n_30),
.B1(n_32),
.B2(n_16),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_77),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_73),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_28),
.B1(n_24),
.B2(n_18),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_78),
.A2(n_109),
.B1(n_72),
.B2(n_60),
.Y(n_137)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_91),
.B1(n_95),
.B2(n_100),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_85),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_97),
.B1(n_59),
.B2(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_50),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_21),
.B1(n_20),
.B2(n_23),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_101),
.B1(n_102),
.B2(n_110),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_65),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_51),
.A2(n_18),
.B1(n_33),
.B2(n_23),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_82),
.B1(n_81),
.B2(n_89),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_53),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_26),
.B1(n_18),
.B2(n_15),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_26),
.B1(n_9),
.B2(n_14),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_53),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_108),
.Y(n_111)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_53),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_52),
.B(n_53),
.C(n_66),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_112),
.A2(n_22),
.B(n_31),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_58),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_117),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_58),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_137),
.B1(n_96),
.B2(n_97),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_95),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_61),
.B1(n_74),
.B2(n_59),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_126),
.A2(n_130),
.B1(n_136),
.B2(n_67),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_90),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_57),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_138),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_61),
.B1(n_74),
.B2(n_59),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_86),
.B1(n_87),
.B2(n_91),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_87),
.A2(n_63),
.B1(n_68),
.B2(n_72),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_82),
.B(n_22),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_79),
.B(n_81),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_139),
.B(n_79),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_98),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_150),
.B(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_145),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_144),
.B(n_149),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_134),
.B(n_76),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_151),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_139),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_118),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_156),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_109),
.C(n_67),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_157),
.C(n_136),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_107),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_78),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_99),
.B1(n_96),
.B2(n_88),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_168),
.Y(n_207)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_112),
.A2(n_67),
.B(n_90),
.C(n_99),
.D(n_33),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_132),
.C(n_127),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_112),
.A2(n_99),
.B(n_105),
.C(n_96),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_103),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_163),
.B(n_169),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_165)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_22),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_119),
.Y(n_181)
);

AOI32xp33_ASAP7_75t_L g167 ( 
.A1(n_118),
.A2(n_67),
.A3(n_103),
.B1(n_31),
.B2(n_33),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_172),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_121),
.B(n_11),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_118),
.A2(n_0),
.B(n_1),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_136),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_173)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_176),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_177),
.B(n_180),
.Y(n_212)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_170),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_201),
.Y(n_214)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_117),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_190),
.C(n_191),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_138),
.C(n_121),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_127),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_196),
.C(n_155),
.Y(n_228)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_195),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_127),
.C(n_119),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_199),
.Y(n_208)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_150),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_203),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_204),
.A2(n_200),
.B1(n_199),
.B2(n_153),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_205),
.A2(n_172),
.B(n_141),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_228),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_224),
.B1(n_225),
.B2(n_229),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_204),
.A2(n_201),
.B1(n_193),
.B2(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_150),
.C(n_143),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_194),
.C(n_188),
.Y(n_237)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_186),
.A2(n_132),
.B1(n_149),
.B2(n_145),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_154),
.B1(n_167),
.B2(n_158),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_157),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_196),
.C(n_175),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_158),
.B1(n_159),
.B2(n_164),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_231),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_141),
.B1(n_161),
.B2(n_155),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_208),
.B1(n_219),
.B2(n_234),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_192),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_233),
.B(n_131),
.Y(n_259)
);

XOR2x2_ASAP7_75t_L g234 ( 
.A(n_174),
.B(n_166),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_234),
.A2(n_189),
.B(n_202),
.Y(n_248)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_178),
.Y(n_244)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_195),
.C(n_219),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_197),
.Y(n_239)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_251),
.C(n_228),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_175),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_226),
.Y(n_264)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_244),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_215),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_247),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_182),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_249),
.B(n_214),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_174),
.C(n_182),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_257),
.Y(n_278)
);

NOR2x1_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_181),
.Y(n_253)
);

OAI22x1_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_179),
.B1(n_198),
.B2(n_197),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_161),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_255),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g257 ( 
.A1(n_209),
.A2(n_173),
.B(n_184),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_206),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_258),
.B(n_227),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_259),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_248),
.A2(n_214),
.B(n_208),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_260),
.A2(n_253),
.B(n_249),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_262),
.A2(n_256),
.B1(n_184),
.B2(n_245),
.Y(n_293)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_267),
.C(n_268),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_250),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_222),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_270),
.C(n_271),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_225),
.C(n_232),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_215),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_220),
.C(n_223),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_277),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_275),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_165),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_231),
.C(n_221),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_281),
.A2(n_265),
.B(n_279),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_236),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_288),
.C(n_289),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_243),
.B1(n_254),
.B2(n_247),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_274),
.B1(n_124),
.B2(n_126),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_266),
.B(n_123),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_286),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_218),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_276),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_255),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_243),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_246),
.Y(n_291)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_273),
.A2(n_256),
.B1(n_241),
.B2(n_238),
.Y(n_294)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_272),
.C(n_267),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_303),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_300),
.A2(n_10),
.B(n_1),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_269),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_292),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_125),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_295),
.B1(n_280),
.B2(n_283),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_169),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_309),
.Y(n_317)
);

OAI322xp33_ASAP7_75t_L g307 ( 
.A1(n_282),
.A2(n_264),
.A3(n_268),
.B1(n_137),
.B2(n_113),
.C1(n_126),
.C2(n_120),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_307),
.A2(n_300),
.B(n_298),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_120),
.C(n_113),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_310),
.B(n_315),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_294),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_311),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_297),
.C(n_299),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_289),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_301),
.A2(n_130),
.B1(n_292),
.B2(n_285),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_SL g320 ( 
.A1(n_316),
.A2(n_318),
.B(n_298),
.C(n_301),
.Y(n_320)
);

AOI322xp5_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_305),
.A3(n_297),
.B1(n_302),
.B2(n_10),
.C1(n_5),
.C2(n_6),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_320),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_323),
.Y(n_329)
);

AOI31xp67_ASAP7_75t_L g328 ( 
.A1(n_324),
.A2(n_327),
.A3(n_3),
.B(n_4),
.Y(n_328)
);

AOI322xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_305),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_0),
.C2(n_6),
.Y(n_325)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_320),
.B(n_5),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_3),
.C(n_4),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_326),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_8),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_332),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_322),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_334),
.C(n_329),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_331),
.C(n_316),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_338)
);


endmodule