module fake_jpeg_17346_n_219 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVxp33_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_28),
.B(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_7),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_7),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_27),
.B1(n_21),
.B2(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_0),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_14),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_48),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_24),
.B1(n_17),
.B2(n_21),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_28),
.B(n_21),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_50),
.B1(n_41),
.B2(n_39),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_20),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_24),
.B1(n_26),
.B2(n_18),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_18),
.B1(n_16),
.B2(n_24),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_16),
.B1(n_24),
.B2(n_15),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_29),
.A2(n_22),
.B1(n_27),
.B2(n_19),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_38),
.B1(n_27),
.B2(n_32),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_60),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_0),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_72),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_66),
.B1(n_45),
.B2(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_46),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_65),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_36),
.B1(n_32),
.B2(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_0),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_46),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_90),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_56),
.A3(n_71),
.B1(n_70),
.B2(n_60),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_85),
.B1(n_56),
.B2(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_100),
.B1(n_74),
.B2(n_76),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_97),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_50),
.B(n_56),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_99),
.B(n_108),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_88),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_54),
.B(n_67),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_70),
.B1(n_39),
.B2(n_69),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_33),
.C(n_63),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_105),
.C(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_107),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_39),
.B1(n_47),
.B2(n_43),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_34),
.C(n_55),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_83),
.C(n_88),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_81),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_98),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_79),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_112),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_119),
.B(n_120),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_84),
.B1(n_78),
.B2(n_85),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_123),
.B1(n_47),
.B2(n_68),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_117),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_76),
.A3(n_75),
.B1(n_73),
.B2(n_85),
.C1(n_52),
.C2(n_81),
.Y(n_114)
);

NOR4xp25_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_40),
.C(n_34),
.D(n_19),
.Y(n_142)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_106),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_77),
.B(n_87),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_77),
.B(n_27),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_102),
.B1(n_103),
.B2(n_94),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_107),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_110),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_55),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_135),
.C(n_144),
.Y(n_149)
);

AOI22x1_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_90),
.B1(n_86),
.B2(n_68),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_141),
.B1(n_137),
.B2(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_51),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_136),
.B(n_138),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_39),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_121),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_91),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

XNOR2x2_ASAP7_75t_SL g156 ( 
.A(n_142),
.B(n_115),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_47),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_125),
.C(n_117),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_19),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_150),
.C(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_133),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_110),
.C(n_113),
.Y(n_154)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_133),
.B1(n_140),
.B2(n_130),
.C(n_131),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_111),
.C(n_118),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_159),
.C(n_132),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_120),
.C(n_114),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_158),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_163),
.B1(n_169),
.B2(n_9),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_153),
.B1(n_152),
.B2(n_159),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_164),
.B(n_170),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_157),
.B(n_131),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_168),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_127),
.B1(n_90),
.B2(n_10),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_149),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_86),
.C(n_59),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_174),
.C(n_145),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_86),
.C(n_40),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_178),
.C(n_185),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_156),
.C(n_86),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_8),
.B(n_13),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_179),
.A2(n_181),
.B(n_13),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_8),
.B(n_13),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_9),
.Y(n_182)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_171),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_40),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_22),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_7),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_186),
.B(n_10),
.Y(n_193)
);

OAI21x1_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_166),
.B(n_174),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_190),
.Y(n_198)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_184),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_22),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_167),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_90),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_177),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_192),
.B(n_193),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_196),
.B(n_12),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_195),
.A2(n_180),
.B(n_185),
.C(n_178),
.D(n_11),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_200),
.C(n_201),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_195),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_204),
.B(n_190),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_205),
.B(n_206),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_202),
.A2(n_191),
.B(n_11),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_0),
.C(n_1),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_3),
.Y(n_213)
);

AOI21x1_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_1),
.B(n_2),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_210),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_208),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_1),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_213),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_SL g217 ( 
.A1(n_215),
.A2(n_214),
.B(n_4),
.C(n_5),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_216),
.B(n_4),
.C(n_6),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_3),
.C(n_4),
.Y(n_219)
);


endmodule