module fake_jpeg_3611_n_213 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_213);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_12),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_17),
.B(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_0),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_0),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_68),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_77),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_2),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_61),
.C(n_48),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_65),
.B1(n_58),
.B2(n_69),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_75),
.B1(n_65),
.B2(n_79),
.Y(n_104)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_69),
.B1(n_58),
.B2(n_55),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_78),
.B1(n_56),
.B2(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_94),
.B(n_51),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_67),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_81),
.B(n_74),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g119 ( 
.A(n_103),
.Y(n_119)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_75),
.B1(n_91),
.B2(n_79),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_48),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_71),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_54),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_113),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_56),
.B1(n_54),
.B2(n_63),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_65),
.Y(n_126)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_63),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_91),
.B1(n_88),
.B2(n_89),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_133),
.B1(n_66),
.B2(n_59),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_59),
.Y(n_147)
);

NAND2x1_ASAP7_75t_SL g118 ( 
.A(n_107),
.B(n_79),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_98),
.B(n_106),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_68),
.C(n_53),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_132),
.C(n_79),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_71),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_3),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_125),
.B(n_131),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_103),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_53),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_53),
.B1(n_60),
.B2(n_66),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_98),
.B(n_97),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_143),
.B(n_5),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_121),
.B(n_97),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_139),
.C(n_145),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_53),
.C(n_49),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_150),
.C(n_6),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_123),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_59),
.B1(n_49),
.B2(n_66),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_3),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_144),
.B(n_149),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_130),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_147),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_49),
.B(n_5),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_13),
.B(n_14),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_23),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_119),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_151),
.B(n_156),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_24),
.B1(n_43),
.B2(n_42),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_115),
.B(n_120),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_163),
.B(n_31),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_172),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_45),
.B(n_41),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_154),
.B(n_4),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_164),
.B(n_169),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_155),
.C(n_143),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_136),
.B(n_8),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_175),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_11),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_14),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_139),
.C(n_140),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_181),
.C(n_29),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_142),
.B(n_141),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_183),
.A2(n_171),
.B(n_159),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_176),
.A2(n_171),
.B1(n_170),
.B2(n_162),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_189),
.B(n_177),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_185),
.B(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_21),
.B(n_38),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_15),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_182),
.B(n_180),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_193),
.B(n_196),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_167),
.A3(n_165),
.B1(n_172),
.B2(n_168),
.C1(n_174),
.C2(n_163),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_195),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_35),
.C(n_39),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_187),
.B(n_28),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_197),
.A2(n_190),
.B1(n_37),
.B2(n_40),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_202),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_190),
.B(n_188),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_203),
.B(n_36),
.Y(n_205)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_205),
.A2(n_200),
.B1(n_201),
.B2(n_18),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_204),
.A2(n_15),
.B(n_17),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_207),
.B(n_18),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_209),
.B(n_206),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_19),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_19),
.Y(n_213)
);


endmodule