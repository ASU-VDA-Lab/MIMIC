module fake_netlist_6_302_n_68 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_68);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_68;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_24;
wire n_37;
wire n_33;
wire n_54;
wire n_67;
wire n_27;
wire n_38;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_55;
wire n_35;
wire n_28;
wire n_58;
wire n_23;
wire n_50;
wire n_49;
wire n_30;
wire n_64;
wire n_43;
wire n_47;
wire n_48;
wire n_29;
wire n_62;
wire n_31;
wire n_65;
wire n_25;
wire n_40;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx4_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

AND2x4_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_4),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_14),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_26),
.B(n_2),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_3),
.B1(n_20),
.B2(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_22),
.B(n_3),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_24),
.B(n_32),
.Y(n_48)
);

OAI21x1_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_36),
.B(n_28),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_32),
.B(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

OAI21x1_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_41),
.B(n_45),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

AOI222xp33_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_45),
.B1(n_44),
.B2(n_41),
.C1(n_39),
.C2(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_59),
.B(n_58),
.Y(n_62)
);

OAI221xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_61),
.B1(n_22),
.B2(n_42),
.C(n_37),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_SL g64 ( 
.A(n_63),
.B(n_53),
.C(n_30),
.Y(n_64)
);

AOI222xp33_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_23),
.B1(n_30),
.B2(n_31),
.C1(n_42),
.C2(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);


endmodule