module fake_jpeg_24377_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_7),
.B(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_40),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_7),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_34),
.Y(n_74)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

OR2x2_ASAP7_75t_SL g47 ( 
.A(n_28),
.B(n_0),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_28),
.C(n_34),
.Y(n_76)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_52),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_16),
.B1(n_32),
.B2(n_19),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_57),
.B1(n_75),
.B2(n_37),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_16),
.B1(n_19),
.B2(n_32),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_54),
.B1(n_68),
.B2(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_32),
.B1(n_28),
.B2(n_22),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_33),
.B1(n_25),
.B2(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_17),
.Y(n_62)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_24),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_67),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_28),
.B1(n_33),
.B2(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_24),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_69),
.Y(n_110)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_74),
.B(n_9),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_37),
.A2(n_25),
.B1(n_33),
.B2(n_28),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_15),
.Y(n_84)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_SL g118 ( 
.A1(n_78),
.A2(n_84),
.B(n_101),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_79),
.A2(n_42),
.B1(n_66),
.B2(n_21),
.Y(n_126)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_95),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_37),
.B1(n_18),
.B2(n_47),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_89),
.B1(n_90),
.B2(n_75),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_85),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_40),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_18),
.B1(n_26),
.B2(n_21),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_26),
.B1(n_21),
.B2(n_35),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_94),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_29),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_44),
.B1(n_45),
.B2(n_30),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_66),
.B1(n_77),
.B2(n_65),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_29),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_105),
.Y(n_135)
);

CKINVDCx9p33_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_44),
.B1(n_45),
.B2(n_42),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_104),
.B(n_111),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_35),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_35),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_72),
.B(n_9),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_0),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_35),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_133),
.B1(n_144),
.B2(n_104),
.Y(n_158)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_42),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_140),
.C(n_111),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_54),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_133),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_126),
.B1(n_100),
.B2(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_123),
.B(n_136),
.Y(n_155)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_134),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_80),
.A2(n_61),
.B1(n_49),
.B2(n_70),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_127),
.A2(n_131),
.B1(n_114),
.B2(n_109),
.Y(n_172)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_30),
.B1(n_23),
.B2(n_73),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_132),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_78),
.A2(n_30),
.B1(n_23),
.B2(n_2),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_93),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_12),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_141),
.Y(n_154)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_83),
.B(n_12),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_146),
.A2(n_3),
.B(n_4),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_134),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_147),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_85),
.B(n_112),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_148),
.A2(n_150),
.B(n_171),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_84),
.B1(n_82),
.B2(n_105),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_159),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_156),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_158),
.B1(n_166),
.B2(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_84),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_163),
.Y(n_180)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_102),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_165),
.Y(n_192)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_177),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_128),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_168),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_125),
.A2(n_130),
.B1(n_120),
.B2(n_135),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_169),
.A2(n_179),
.B1(n_130),
.B2(n_135),
.Y(n_187)
);

AO22x2_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_91),
.B1(n_95),
.B2(n_103),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_142),
.B1(n_133),
.B2(n_124),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_128),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_173),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_86),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_174),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_106),
.Y(n_175)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_106),
.C(n_82),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_143),
.B(n_110),
.Y(n_183)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_117),
.A2(n_110),
.B1(n_113),
.B2(n_87),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_183),
.B(n_195),
.Y(n_224)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_207),
.B1(n_170),
.B2(n_205),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_206),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_177),
.A2(n_125),
.B1(n_131),
.B2(n_145),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_188),
.A2(n_189),
.B1(n_168),
.B2(n_166),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_148),
.A2(n_145),
.B1(n_113),
.B2(n_87),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_196),
.B(n_198),
.Y(n_238)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_146),
.A2(n_143),
.B(n_1),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_202),
.A2(n_209),
.B(n_153),
.Y(n_217)
);

A2O1A1O1Ixp25_ASAP7_75t_L g203 ( 
.A1(n_169),
.A2(n_11),
.B(n_10),
.C(n_8),
.D(n_4),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_179),
.C(n_160),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_0),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

AOI21x1_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_0),
.B(n_1),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_210),
.B(n_173),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_155),
.Y(n_206)
);

AOI22x1_ASAP7_75t_SL g207 ( 
.A1(n_170),
.A2(n_98),
.B1(n_10),
.B2(n_8),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_150),
.A2(n_1),
.B(n_3),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_178),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_187),
.B(n_158),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_213),
.B(n_214),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_159),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_221),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_217),
.A2(n_227),
.B(n_204),
.Y(n_262)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_212),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_147),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_231),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_151),
.C(n_165),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_228),
.C(n_229),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_170),
.Y(n_226)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_172),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_164),
.C(n_171),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_212),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_186),
.B(n_167),
.C(n_4),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_236),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_193),
.B1(n_229),
.B2(n_226),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_3),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_237),
.C(n_239),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_3),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_240),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_186),
.B(n_4),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_5),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_5),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_241),
.A2(n_257),
.B1(n_260),
.B2(n_252),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_238),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_244),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_235),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_214),
.B(n_223),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_252),
.C(n_256),
.Y(n_269)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_215),
.B(n_197),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_216),
.A2(n_185),
.B1(n_182),
.B2(n_233),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_254),
.A2(n_216),
.B1(n_184),
.B2(n_227),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_213),
.B(n_202),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_228),
.A2(n_209),
.B1(n_192),
.B2(n_184),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_192),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_262),
.B(n_255),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_217),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_216),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_265),
.A2(n_276),
.B1(n_258),
.B2(n_251),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_275),
.B(n_280),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_237),
.C(n_220),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_281),
.C(n_283),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_185),
.B1(n_222),
.B2(n_207),
.Y(n_272)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_242),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_273),
.Y(n_295)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_194),
.B(n_210),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_246),
.A2(n_195),
.B1(n_184),
.B2(n_220),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_282),
.B1(n_274),
.B2(n_266),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_234),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_253),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_249),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_199),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_262),
.A2(n_194),
.B(n_181),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_181),
.C(n_180),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_200),
.B1(n_199),
.B2(n_206),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_211),
.C(n_203),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_278),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_248),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_287),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_256),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_245),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_288),
.B(n_289),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_298),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_294),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_282),
.A2(n_255),
.B1(n_258),
.B2(n_261),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_297),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_266),
.B(n_251),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_285),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_281),
.C(n_271),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_302),
.C(n_283),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_269),
.C(n_280),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_295),
.B(n_264),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_303),
.B(n_308),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_293),
.A2(n_284),
.B(n_292),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_310),
.B(n_311),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_208),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_269),
.B(n_275),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_267),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_250),
.Y(n_312)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_312),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_307),
.A2(n_290),
.B(n_296),
.Y(n_313)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_313),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_320),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_265),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_301),
.C(n_302),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_253),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_304),
.Y(n_321)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_321),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_183),
.Y(n_324)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_324),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_318),
.C(n_319),
.Y(n_329)
);

AOI322xp5_ASAP7_75t_L g333 ( 
.A1(n_329),
.A2(n_6),
.A3(n_309),
.B1(n_323),
.B2(n_322),
.C1(n_328),
.C2(n_320),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_315),
.Y(n_330)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g332 ( 
.A1(n_330),
.A2(n_325),
.B(n_323),
.C(n_327),
.D(n_326),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_333),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_331),
.Y(n_336)
);


endmodule