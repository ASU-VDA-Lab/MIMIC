module fake_jpeg_6664_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx9p33_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_17),
.Y(n_22)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_0),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_20),
.B(n_13),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_24),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_8),
.B1(n_14),
.B2(n_15),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_25),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_29),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_19),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_14),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_19),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_15),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_18),
.C(n_17),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_31),
.B1(n_29),
.B2(n_23),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_40),
.B1(n_43),
.B2(n_12),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_23),
.B1(n_8),
.B2(n_11),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_12),
.B1(n_10),
.B2(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_12),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_48),
.B1(n_39),
.B2(n_41),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_1),
.C(n_2),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_49),
.B1(n_51),
.B2(n_43),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_42),
.B1(n_4),
.B2(n_5),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_2),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_54),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_55),
.B(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_58),
.B(n_6),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_7),
.Y(n_60)
);


endmodule