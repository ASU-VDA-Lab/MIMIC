module fake_jpeg_11214_n_24 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_0),
.B(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_1),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx12_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

AND2x4_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_7),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_17),
.C(n_18),
.Y(n_21)
);

OAI32xp33_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_0),
.A3(n_1),
.B1(n_4),
.B2(n_8),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_13),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_10),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_20),
.B(n_12),
.C(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_15),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_18),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_23),
.A2(n_21),
.B1(n_16),
.B2(n_11),
.Y(n_24)
);


endmodule