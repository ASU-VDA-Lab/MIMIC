module fake_netlist_6_728_n_770 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_770);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_770;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_575;
wire n_368;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_153;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_508;
wire n_361;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_23),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_9),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_135),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_56),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_13),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_27),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_31),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_109),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_100),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_28),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_71),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_99),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_124),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_23),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_62),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_10),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_41),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_83),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_87),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_11),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_36),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_50),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_103),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_86),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_10),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_67),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_20),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_73),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_15),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_13),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_47),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_21),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_3),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_108),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_3),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_25),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_66),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_91),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_74),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_106),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_75),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_5),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_33),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_192),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_152),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_0),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_147),
.B(n_0),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_147),
.B(n_1),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_1),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_2),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_147),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_147),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_2),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_4),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_148),
.Y(n_219)
);

AND2x6_ASAP7_75t_L g220 ( 
.A(n_148),
.B(n_26),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_147),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_151),
.Y(n_224)
);

BUFx8_ASAP7_75t_SL g225 ( 
.A(n_169),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_147),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_149),
.B(n_4),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_146),
.B(n_5),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_164),
.B(n_6),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_164),
.B(n_6),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_150),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_171),
.B(n_7),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_155),
.B(n_7),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_172),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_188),
.B1(n_167),
.B2(n_157),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_210),
.A2(n_174),
.B1(n_192),
.B2(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_160),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_210),
.A2(n_179),
.B1(n_184),
.B2(n_191),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_216),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_153),
.Y(n_246)
);

AND2x2_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_8),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_229),
.A2(n_197),
.B1(n_193),
.B2(n_189),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_186),
.B1(n_183),
.B2(n_181),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_178),
.B1(n_177),
.B2(n_176),
.Y(n_250)
);

AO22x2_ASAP7_75t_L g251 ( 
.A1(n_205),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_R g252 ( 
.A1(n_235),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_252)
);

AO22x2_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_217),
.B1(n_209),
.B2(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_206),
.A2(n_175),
.B1(n_170),
.B2(n_166),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_12),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

NAND2xp33_ASAP7_75t_SL g258 ( 
.A(n_209),
.B(n_156),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_208),
.A2(n_165),
.B1(n_163),
.B2(n_162),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_237),
.A2(n_161),
.B1(n_158),
.B2(n_17),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_204),
.B(n_230),
.Y(n_262)
);

OR2x6_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_14),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_29),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_217),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_265)
);

AO22x2_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_213),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_220),
.B(n_19),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g269 ( 
.A1(n_238),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_30),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_236),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_201),
.A2(n_24),
.B1(n_32),
.B2(n_34),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_213),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_236),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_236),
.B(n_39),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_40),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_239),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_200),
.B(n_45),
.Y(n_280)
);

AND2x4_ASAP7_75t_L g281 ( 
.A(n_227),
.B(n_46),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_219),
.Y(n_282)
);

AO22x2_ASAP7_75t_L g283 ( 
.A1(n_223),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_213),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_223),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_L g286 ( 
.A1(n_223),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_227),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_200),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_219),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_243),
.B(n_223),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_241),
.B(n_225),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_241),
.B(n_59),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_200),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_242),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_249),
.B(n_60),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_246),
.B(n_219),
.Y(n_301)
);

AND2x6_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_215),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_259),
.B(n_200),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_259),
.B(n_200),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_244),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_249),
.B(n_226),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_245),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_254),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_244),
.B(n_226),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_240),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_R g313 ( 
.A(n_263),
.B(n_61),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_256),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_284),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_273),
.B(n_63),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_255),
.B(n_219),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_258),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_263),
.B(n_226),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_253),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_247),
.B(n_219),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_253),
.B(n_219),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_270),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_266),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_266),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_268),
.A2(n_222),
.B(n_215),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_283),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_221),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_251),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_265),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_251),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_260),
.Y(n_341)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_285),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_279),
.B(n_64),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_279),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_275),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_252),
.B(n_221),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_272),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_267),
.Y(n_348)
);

AND2x6_ASAP7_75t_L g349 ( 
.A(n_264),
.B(n_215),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_257),
.B(n_222),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_324),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_327),
.A2(n_220),
.B(n_222),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_287),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_319),
.B(n_221),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_289),
.B(n_221),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_290),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_221),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_302),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_309),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_348),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_322),
.B(n_200),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_293),
.B(n_221),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_301),
.B(n_220),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_314),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_295),
.B(n_322),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_321),
.B(n_202),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_350),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_292),
.B(n_202),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_301),
.B(n_220),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_327),
.A2(n_220),
.B(n_212),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_316),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_315),
.B(n_65),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_292),
.B(n_202),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_202),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_350),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_323),
.A2(n_318),
.B(n_344),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_338),
.Y(n_382)
);

AND2x2_ASAP7_75t_SL g383 ( 
.A(n_342),
.B(n_220),
.Y(n_383)
);

INVx3_ASAP7_75t_SL g384 ( 
.A(n_308),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_288),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_347),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_325),
.B(n_220),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_330),
.B(n_220),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_331),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_318),
.B(n_202),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_294),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_320),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_332),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_297),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_345),
.A2(n_212),
.B(n_214),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_334),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_300),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_337),
.B(n_68),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_339),
.B(n_69),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_302),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_302),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_312),
.B(n_70),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_313),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_338),
.B(n_218),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_332),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_291),
.B(n_218),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_335),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_342),
.B(n_218),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_328),
.B(n_346),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_302),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_302),
.B(n_218),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_298),
.B(n_72),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_303),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_359),
.B(n_328),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_359),
.B(n_304),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_363),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_370),
.B(n_340),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_413),
.B(n_346),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_370),
.B(n_326),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_363),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_336),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_381),
.B(n_306),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_406),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_363),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_401),
.B(n_336),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_341),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_363),
.Y(n_432)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_392),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_76),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_400),
.B(n_317),
.Y(n_437)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_360),
.Y(n_438)
);

INVx8_ASAP7_75t_L g439 ( 
.A(n_408),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_363),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_382),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_349),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_382),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_372),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_349),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_353),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_371),
.B(n_343),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_371),
.B(n_349),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_373),
.B(n_349),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_382),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_411),
.B(n_218),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_372),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_373),
.B(n_296),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_417),
.B(n_354),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_382),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g458 ( 
.A(n_416),
.B(n_218),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_414),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_372),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_378),
.B(n_389),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_408),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_391),
.Y(n_463)
);

BUFx12f_ASAP7_75t_L g464 ( 
.A(n_354),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_401),
.B(n_402),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_378),
.B(n_379),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_402),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_394),
.B(n_77),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_391),
.Y(n_469)
);

OR2x6_ASAP7_75t_L g470 ( 
.A(n_401),
.B(n_214),
.Y(n_470)
);

BUFx4f_ASAP7_75t_L g471 ( 
.A(n_408),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_389),
.B(n_379),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_465),
.B(n_421),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_441),
.Y(n_474)
);

INVx6_ASAP7_75t_L g475 ( 
.A(n_464),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_428),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_423),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_464),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_434),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_433),
.B(n_402),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_469),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_422),
.B(n_384),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_422),
.B(n_384),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_463),
.Y(n_484)
);

NAND2x1p5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_408),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_469),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_463),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_459),
.Y(n_488)
);

BUFx2_ASAP7_75t_SL g489 ( 
.A(n_423),
.Y(n_489)
);

INVx5_ASAP7_75t_SL g490 ( 
.A(n_430),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_423),
.Y(n_491)
);

BUFx12f_ASAP7_75t_L g492 ( 
.A(n_427),
.Y(n_492)
);

INVx6_ASAP7_75t_SL g493 ( 
.A(n_430),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_462),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_426),
.B(n_389),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_437),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_462),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_427),
.Y(n_498)
);

BUFx10_ASAP7_75t_L g499 ( 
.A(n_465),
.Y(n_499)
);

CKINVDCx6p67_ASAP7_75t_R g500 ( 
.A(n_430),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_421),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_436),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_462),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_455),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_455),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_449),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_421),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_426),
.B(n_402),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_425),
.B(n_384),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_430),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_436),
.Y(n_511)
);

NAND2x1p5_ASAP7_75t_L g512 ( 
.A(n_471),
.B(n_408),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_428),
.Y(n_513)
);

BUFx12f_ASAP7_75t_L g514 ( 
.A(n_468),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_445),
.Y(n_515)
);

BUFx12f_ASAP7_75t_L g516 ( 
.A(n_468),
.Y(n_516)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_428),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_449),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_462),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_428),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_498),
.Y(n_521)
);

BUFx4f_ASAP7_75t_SL g522 ( 
.A(n_492),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_484),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_482),
.B(n_425),
.Y(n_524)
);

INVx6_ASAP7_75t_L g525 ( 
.A(n_475),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_508),
.A2(n_418),
.B1(n_416),
.B2(n_431),
.Y(n_526)
);

CKINVDCx11_ASAP7_75t_R g527 ( 
.A(n_492),
.Y(n_527)
);

NAND2x1p5_ASAP7_75t_L g528 ( 
.A(n_517),
.B(n_471),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_475),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_484),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_480),
.A2(n_467),
.B1(n_458),
.B2(n_465),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_480),
.A2(n_467),
.B1(n_458),
.B2(n_465),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_509),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_500),
.A2(n_458),
.B1(n_456),
.B2(n_470),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_500),
.A2(n_470),
.B1(n_472),
.B2(n_461),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_481),
.Y(n_536)
);

NAND2x1p5_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_441),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_486),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_495),
.A2(n_416),
.B1(n_419),
.B2(n_466),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_496),
.A2(n_435),
.B1(n_405),
.B2(n_416),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_483),
.A2(n_466),
.B1(n_435),
.B2(n_377),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_498),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_509),
.A2(n_435),
.B1(n_361),
.B2(n_362),
.Y(n_543)
);

HB1xp67_ASAP7_75t_SL g544 ( 
.A(n_505),
.Y(n_544)
);

BUFx4_ASAP7_75t_SL g545 ( 
.A(n_506),
.Y(n_545)
);

INVx6_ASAP7_75t_L g546 ( 
.A(n_475),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_487),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_488),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_490),
.A2(n_470),
.B1(n_438),
.B2(n_433),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_514),
.A2(n_435),
.B1(n_447),
.B2(n_439),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_514),
.A2(n_439),
.B1(n_383),
.B2(n_462),
.Y(n_551)
);

BUFx4f_ASAP7_75t_L g552 ( 
.A(n_516),
.Y(n_552)
);

CKINVDCx11_ASAP7_75t_R g553 ( 
.A(n_479),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_491),
.B(n_510),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_510),
.A2(n_361),
.B1(n_362),
.B2(n_365),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_505),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_SL g557 ( 
.A1(n_516),
.A2(n_439),
.B1(n_383),
.B2(n_441),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_499),
.Y(n_558)
);

CKINVDCx11_ASAP7_75t_R g559 ( 
.A(n_504),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_517),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_490),
.A2(n_470),
.B1(n_438),
.B2(n_433),
.Y(n_561)
);

AOI222xp33_ASAP7_75t_L g562 ( 
.A1(n_524),
.A2(n_506),
.B1(n_477),
.B2(n_559),
.C1(n_504),
.C2(n_526),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_523),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_560),
.Y(n_564)
);

BUFx12f_ASAP7_75t_L g565 ( 
.A(n_527),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_SL g566 ( 
.A1(n_534),
.A2(n_518),
.B1(n_490),
.B2(n_489),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_540),
.A2(n_369),
.B1(n_365),
.B2(n_493),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_536),
.Y(n_568)
);

OAI222xp33_ASAP7_75t_L g569 ( 
.A1(n_543),
.A2(n_478),
.B1(n_502),
.B2(n_515),
.C1(n_511),
.C2(n_512),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_525),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_SL g571 ( 
.A1(n_522),
.A2(n_383),
.B1(n_443),
.B2(n_428),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_538),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_547),
.Y(n_573)
);

INVx5_ASAP7_75t_SL g574 ( 
.A(n_545),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_529),
.B(n_473),
.Y(n_575)
);

AOI222xp33_ASAP7_75t_L g576 ( 
.A1(n_526),
.A2(n_351),
.B1(n_473),
.B2(n_507),
.C1(n_501),
.C2(n_385),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_541),
.A2(n_473),
.B1(n_493),
.B2(n_507),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_523),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_554),
.B(n_501),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_541),
.A2(n_493),
.B1(n_386),
.B2(n_369),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_543),
.A2(n_386),
.B1(n_385),
.B2(n_376),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_556),
.B(n_398),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_530),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_533),
.B(n_398),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_539),
.A2(n_386),
.B1(n_376),
.B2(n_380),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_539),
.A2(n_376),
.B1(n_380),
.B2(n_451),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_558),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_530),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_533),
.A2(n_451),
.B1(n_391),
.B2(n_367),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_555),
.A2(n_367),
.B1(n_390),
.B2(n_454),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_521),
.A2(n_450),
.B1(n_499),
.B2(n_387),
.Y(n_591)
);

BUFx12f_ASAP7_75t_L g592 ( 
.A(n_553),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_521),
.A2(n_555),
.B1(n_550),
.B2(n_551),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_SL g594 ( 
.A1(n_522),
.A2(n_444),
.B1(n_443),
.B2(n_439),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_548),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_552),
.A2(n_450),
.B1(n_499),
.B2(n_387),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_548),
.B(n_542),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_557),
.A2(n_485),
.B1(n_512),
.B2(n_503),
.Y(n_598)
);

BUFx12f_ASAP7_75t_L g599 ( 
.A(n_525),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_525),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_558),
.Y(n_601)
);

OAI21xp33_ASAP7_75t_L g602 ( 
.A1(n_535),
.A2(n_356),
.B(n_355),
.Y(n_602)
);

BUFx8_ASAP7_75t_SL g603 ( 
.A(n_552),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_SL g604 ( 
.A1(n_531),
.A2(n_444),
.B1(n_443),
.B2(n_432),
.Y(n_604)
);

AOI222xp33_ASAP7_75t_L g605 ( 
.A1(n_532),
.A2(n_387),
.B1(n_352),
.B2(n_375),
.C1(n_397),
.C2(n_395),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_546),
.A2(n_445),
.B1(n_454),
.B2(n_460),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_544),
.A2(n_366),
.B1(n_408),
.B2(n_387),
.Y(n_607)
);

BUFx12f_ASAP7_75t_L g608 ( 
.A(n_546),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_546),
.A2(n_460),
.B1(n_395),
.B2(n_397),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_562),
.A2(n_432),
.B1(n_424),
.B2(n_364),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_566),
.A2(n_424),
.B1(n_358),
.B2(n_364),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_597),
.B(n_488),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_L g613 ( 
.A(n_576),
.B(n_567),
.C(n_593),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_566),
.A2(n_364),
.B1(n_357),
.B2(n_358),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_568),
.B(n_497),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_567),
.A2(n_358),
.B1(n_357),
.B2(n_420),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_578),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_579),
.B(n_519),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_SL g619 ( 
.A1(n_574),
.A2(n_561),
.B1(n_549),
.B2(n_485),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_571),
.A2(n_528),
.B1(n_438),
.B2(n_433),
.Y(n_620)
);

OAI221xp5_ASAP7_75t_L g621 ( 
.A1(n_580),
.A2(n_396),
.B1(n_412),
.B2(n_528),
.C(n_357),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_573),
.B(n_440),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_577),
.A2(n_457),
.B1(n_420),
.B2(n_393),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_572),
.B(n_440),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_591),
.A2(n_457),
.B1(n_393),
.B2(n_399),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_SL g626 ( 
.A1(n_574),
.A2(n_443),
.B1(n_444),
.B2(n_560),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_563),
.B(n_448),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_604),
.A2(n_393),
.B1(n_403),
.B2(n_399),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_571),
.A2(n_433),
.B1(n_438),
.B2(n_393),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_595),
.B(n_448),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_604),
.A2(n_404),
.B1(n_403),
.B2(n_399),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_583),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_575),
.A2(n_404),
.B1(n_403),
.B2(n_443),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_575),
.A2(n_586),
.B1(n_596),
.B2(n_574),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_598),
.A2(n_404),
.B1(n_444),
.B2(n_442),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_589),
.A2(n_444),
.B1(n_446),
.B2(n_429),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_588),
.B(n_476),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_584),
.B(n_429),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_589),
.A2(n_452),
.B1(n_429),
.B2(n_414),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_569),
.A2(n_388),
.B(n_537),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_585),
.A2(n_452),
.B1(n_414),
.B2(n_368),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_582),
.A2(n_452),
.B1(n_374),
.B2(n_388),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_601),
.B(n_476),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_581),
.A2(n_590),
.B1(n_609),
.B2(n_594),
.Y(n_644)
);

AOI222xp33_ASAP7_75t_L g645 ( 
.A1(n_565),
.A2(n_388),
.B1(n_407),
.B2(n_453),
.C1(n_459),
.C2(n_415),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_592),
.A2(n_388),
.B1(n_474),
.B2(n_494),
.Y(n_646)
);

NOR3xp33_ASAP7_75t_L g647 ( 
.A(n_613),
.B(n_619),
.C(n_644),
.Y(n_647)
);

AOI221xp5_ASAP7_75t_L g648 ( 
.A1(n_613),
.A2(n_607),
.B1(n_600),
.B2(n_570),
.C(n_602),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_618),
.B(n_612),
.Y(n_649)
);

OAI221xp5_ASAP7_75t_L g650 ( 
.A1(n_646),
.A2(n_594),
.B1(n_587),
.B2(n_609),
.C(n_590),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_615),
.B(n_587),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_640),
.A2(n_605),
.B(n_603),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_615),
.B(n_564),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_617),
.B(n_564),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_617),
.B(n_564),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_632),
.B(n_564),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_632),
.B(n_599),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_645),
.B(n_606),
.C(n_409),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_634),
.A2(n_606),
.B1(n_608),
.B2(n_537),
.Y(n_659)
);

OAI211xp5_ASAP7_75t_L g660 ( 
.A1(n_640),
.A2(n_494),
.B(n_203),
.C(n_202),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_SL g661 ( 
.A(n_643),
.B(n_494),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_638),
.B(n_474),
.Y(n_662)
);

AOI221xp5_ASAP7_75t_L g663 ( 
.A1(n_644),
.A2(n_203),
.B1(n_207),
.B2(n_214),
.C(n_211),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_645),
.B(n_513),
.C(n_476),
.Y(n_664)
);

NAND4xp25_ASAP7_75t_L g665 ( 
.A(n_642),
.B(n_459),
.C(n_474),
.D(n_360),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_637),
.B(n_476),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_637),
.B(n_513),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_630),
.B(n_643),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_630),
.B(n_513),
.Y(n_669)
);

NAND4xp25_ASAP7_75t_L g670 ( 
.A(n_635),
.B(n_610),
.C(n_611),
.D(n_624),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_620),
.B(n_629),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_622),
.B(n_513),
.Y(n_672)
);

AOI221xp5_ASAP7_75t_L g673 ( 
.A1(n_614),
.A2(n_214),
.B1(n_211),
.B2(n_207),
.C(n_203),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_627),
.B(n_78),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_636),
.B(n_79),
.Y(n_675)
);

OAI221xp5_ASAP7_75t_SL g676 ( 
.A1(n_628),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.C(n_85),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_668),
.Y(n_677)
);

AOI211xp5_ASAP7_75t_L g678 ( 
.A1(n_647),
.A2(n_652),
.B(n_676),
.C(n_664),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_649),
.B(n_626),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_657),
.Y(n_680)
);

OAI211xp5_ASAP7_75t_SL g681 ( 
.A1(n_647),
.A2(n_633),
.B(n_631),
.C(n_623),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_648),
.B(n_661),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_653),
.B(n_639),
.Y(n_683)
);

NOR3xp33_ASAP7_75t_L g684 ( 
.A(n_660),
.B(n_621),
.C(n_616),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_651),
.B(n_625),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_655),
.B(n_88),
.Y(n_686)
);

NAND3xp33_ASAP7_75t_L g687 ( 
.A(n_663),
.B(n_641),
.C(n_214),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_656),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_654),
.B(n_662),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_666),
.B(n_89),
.Y(n_690)
);

NAND3xp33_ASAP7_75t_L g691 ( 
.A(n_671),
.B(n_214),
.C(n_207),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_669),
.B(n_90),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_688),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_688),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_677),
.B(n_667),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_678),
.B(n_671),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_680),
.Y(n_697)
);

INVxp67_ASAP7_75t_SL g698 ( 
.A(n_689),
.Y(n_698)
);

XNOR2xp5_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_659),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_677),
.B(n_672),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_680),
.B(n_670),
.Y(n_701)
);

NAND2x1p5_ASAP7_75t_L g702 ( 
.A(n_682),
.B(n_517),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_693),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_697),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_694),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_697),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_698),
.Y(n_707)
);

BUFx2_ASAP7_75t_SL g708 ( 
.A(n_704),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_704),
.Y(n_709)
);

OAI22x1_ASAP7_75t_L g710 ( 
.A1(n_707),
.A2(n_696),
.B1(n_699),
.B2(n_701),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_706),
.A2(n_696),
.B1(n_701),
.B2(n_702),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_SL g712 ( 
.A1(n_706),
.A2(n_702),
.B1(n_679),
.B2(n_691),
.Y(n_712)
);

XNOR2x1_ASAP7_75t_L g713 ( 
.A(n_705),
.B(n_692),
.Y(n_713)
);

OAI322xp33_ASAP7_75t_L g714 ( 
.A1(n_711),
.A2(n_703),
.A3(n_700),
.B1(n_687),
.B2(n_695),
.C1(n_675),
.C2(n_650),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_709),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_708),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_710),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_713),
.Y(n_718)
);

AOI221xp5_ASAP7_75t_L g719 ( 
.A1(n_717),
.A2(n_712),
.B1(n_703),
.B2(n_684),
.C(n_681),
.Y(n_719)
);

NAND4xp75_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_686),
.C(n_690),
.D(n_674),
.Y(n_720)
);

OA22x2_ASAP7_75t_SL g721 ( 
.A1(n_718),
.A2(n_665),
.B1(n_685),
.B2(n_683),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_719),
.Y(n_722)
);

AND4x1_ASAP7_75t_L g723 ( 
.A(n_721),
.B(n_715),
.C(n_714),
.D(n_658),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_SL g724 ( 
.A1(n_720),
.A2(n_685),
.B(n_683),
.C(n_94),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_719),
.Y(n_725)
);

AOI221xp5_ASAP7_75t_L g726 ( 
.A1(n_722),
.A2(n_673),
.B1(n_211),
.B2(n_207),
.C(n_203),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_725),
.A2(n_203),
.B1(n_207),
.B2(n_211),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_723),
.A2(n_203),
.B1(n_207),
.B2(n_211),
.Y(n_728)
);

NOR4xp25_ASAP7_75t_L g729 ( 
.A(n_724),
.B(n_92),
.C(n_93),
.D(n_95),
.Y(n_729)
);

AOI221xp5_ASAP7_75t_L g730 ( 
.A1(n_722),
.A2(n_211),
.B1(n_98),
.B2(n_101),
.C(n_102),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_722),
.A2(n_520),
.B1(n_517),
.B2(n_438),
.Y(n_731)
);

NOR2x1_ASAP7_75t_L g732 ( 
.A(n_728),
.B(n_729),
.Y(n_732)
);

INVxp67_ASAP7_75t_SL g733 ( 
.A(n_727),
.Y(n_733)
);

AND3x2_ASAP7_75t_L g734 ( 
.A(n_730),
.B(n_97),
.C(n_104),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_731),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_726),
.A2(n_520),
.B1(n_438),
.B2(n_433),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_729),
.A2(n_520),
.B1(n_212),
.B2(n_113),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_727),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_737),
.A2(n_520),
.B1(n_212),
.B2(n_114),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_732),
.A2(n_520),
.B1(n_212),
.B2(n_115),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_735),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_733),
.Y(n_742)
);

AND4x1_ASAP7_75t_L g743 ( 
.A(n_738),
.B(n_105),
.C(n_112),
.D(n_116),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_736),
.Y(n_744)
);

NOR2x1_ASAP7_75t_L g745 ( 
.A(n_734),
.B(n_118),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_735),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_737),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_742),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_741),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_746),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_744),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_743),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_740),
.Y(n_753)
);

INVxp67_ASAP7_75t_SL g754 ( 
.A(n_745),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_747),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_739),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_SL g757 ( 
.A1(n_754),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_748),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_752),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_754),
.Y(n_760)
);

OA22x2_ASAP7_75t_L g761 ( 
.A1(n_749),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_758),
.B(n_750),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_760),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_763),
.A2(n_751),
.B1(n_753),
.B2(n_755),
.Y(n_764)
);

AO22x2_ASAP7_75t_L g765 ( 
.A1(n_762),
.A2(n_756),
.B1(n_761),
.B2(n_757),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_765),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_766),
.A2(n_764),
.B1(n_759),
.B2(n_138),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_767),
.Y(n_768)
);

AOI221xp5_ASAP7_75t_L g769 ( 
.A1(n_768),
.A2(n_136),
.B1(n_137),
.B2(n_139),
.C(n_140),
.Y(n_769)
);

AOI211xp5_ASAP7_75t_L g770 ( 
.A1(n_769),
.A2(n_141),
.B(n_142),
.C(n_143),
.Y(n_770)
);


endmodule