module fake_jpeg_15698_n_244 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_244);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_6),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_19),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_26),
.B1(n_29),
.B2(n_27),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_46),
.B1(n_48),
.B2(n_53),
.Y(n_69)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_26),
.B1(n_14),
.B2(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_55),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_26),
.B1(n_19),
.B2(n_20),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_14),
.B1(n_25),
.B2(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_23),
.Y(n_55)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_57),
.A2(n_20),
.B1(n_19),
.B2(n_23),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_60),
.B1(n_65),
.B2(n_82),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_20),
.B1(n_22),
.B2(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_22),
.B1(n_17),
.B2(n_3),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_29),
.B(n_27),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_40),
.B(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_41),
.B(n_10),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_76),
.Y(n_92)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_46),
.B(n_10),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_28),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_29),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_42),
.A2(n_37),
.B(n_31),
.C(n_30),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_97),
.Y(n_116)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_100),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_27),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_72),
.A2(n_40),
.B1(n_50),
.B2(n_37),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_98),
.B1(n_105),
.B2(n_67),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_50),
.B1(n_30),
.B2(n_31),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_104),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_63),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_1),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_82),
.B1(n_71),
.B2(n_1),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_56),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_37),
.B1(n_31),
.B2(n_56),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_119),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_112),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_107),
.B(n_28),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_83),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_86),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_2),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_128),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_28),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_101),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_15),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_86),
.Y(n_127)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_75),
.B1(n_74),
.B2(n_4),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_121),
.B1(n_106),
.B2(n_125),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_27),
.B(n_51),
.C(n_17),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_87),
.B(n_98),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_151),
.B1(n_2),
.B2(n_85),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_96),
.C(n_87),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_122),
.C(n_129),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_91),
.B1(n_95),
.B2(n_92),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_140),
.B1(n_146),
.B2(n_109),
.Y(n_161)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_101),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_84),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_113),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_130),
.A2(n_88),
.B1(n_103),
.B2(n_100),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_108),
.A2(n_94),
.B1(n_89),
.B2(n_105),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_127),
.Y(n_164)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_130),
.B(n_110),
.C(n_117),
.D(n_118),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_138),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_157),
.C(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_123),
.C(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_163),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_112),
.C(n_127),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_124),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_165),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_134),
.B1(n_151),
.B2(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_164),
.A2(n_172),
.B1(n_142),
.B2(n_150),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_84),
.C(n_89),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_167),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_102),
.C(n_79),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_147),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_170),
.C(n_143),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_148),
.B(n_109),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_141),
.B(n_106),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_134),
.B1(n_150),
.B2(n_131),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_144),
.B(n_140),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_85),
.B1(n_128),
.B2(n_51),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_177),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_SL g177 ( 
.A(n_166),
.B(n_132),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_182),
.B(n_183),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_8),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_168),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_146),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_157),
.C(n_165),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g187 ( 
.A(n_153),
.B(n_132),
.CI(n_145),
.CON(n_187),
.SN(n_187)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_187),
.B(n_17),
.Y(n_195)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_155),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_191),
.Y(n_202)
);

AO22x1_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_154),
.B1(n_135),
.B2(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_200),
.C(n_201),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_198),
.Y(n_212)
);

BUFx12_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_149),
.B1(n_85),
.B2(n_5),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_199),
.B(n_185),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_15),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_193),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_196),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_179),
.C(n_176),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_209),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_179),
.C(n_176),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_178),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_199),
.Y(n_222)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_191),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_186),
.B(n_197),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_212),
.B(n_188),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_216),
.B(n_218),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_204),
.B(n_180),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_211),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_SL g228 ( 
.A1(n_220),
.A2(n_221),
.B(n_209),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_192),
.B1(n_189),
.B2(n_174),
.Y(n_221)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_224),
.B(n_207),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_210),
.B(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_226),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_215),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_228),
.B(n_206),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_231),
.A2(n_8),
.B(n_3),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_213),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_7),
.B1(n_3),
.B2(n_5),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_13),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_237),
.B(n_229),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_64),
.C(n_15),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_13),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_238),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_240),
.C(n_7),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_242),
.A2(n_2),
.B1(n_9),
.B2(n_241),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_9),
.Y(n_244)
);


endmodule