module real_aes_8379_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g513 ( .A1(n_0), .A2(n_177), .B(n_514), .C(n_517), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_1), .B(n_509), .Y(n_518) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g175 ( .A(n_3), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_4), .B(n_178), .Y(n_582) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_5), .A2(n_131), .B1(n_134), .B2(n_135), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_5), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_6), .A2(n_477), .B(n_553), .Y(n_552) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_7), .A2(n_185), .B(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_8), .A2(n_38), .B1(n_165), .B2(n_213), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_9), .B(n_185), .Y(n_193) );
AND2x6_ASAP7_75t_L g180 ( .A(n_10), .B(n_181), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_11), .A2(n_180), .B(n_482), .C(n_526), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_12), .A2(n_42), .B1(n_132), .B2(n_133), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_12), .Y(n_132) );
INVx1_ASAP7_75t_L g110 ( .A(n_13), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_13), .B(n_39), .Y(n_127) );
INVx1_ASAP7_75t_L g159 ( .A(n_14), .Y(n_159) );
INVx1_ASAP7_75t_L g156 ( .A(n_15), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_16), .B(n_161), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_17), .B(n_178), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_18), .B(n_152), .Y(n_259) );
AO32x2_ASAP7_75t_L g229 ( .A1(n_19), .A2(n_151), .A3(n_185), .B1(n_204), .B2(n_230), .Y(n_229) );
AOI222xp33_ASAP7_75t_SL g129 ( .A1(n_20), .A2(n_130), .B1(n_136), .B2(n_755), .C1(n_756), .C2(n_758), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_21), .B(n_165), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_22), .B(n_152), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_23), .A2(n_57), .B1(n_165), .B2(n_213), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_24), .Y(n_128) );
AOI22xp33_ASAP7_75t_SL g215 ( .A1(n_25), .A2(n_84), .B1(n_161), .B2(n_165), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_26), .B(n_165), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_27), .A2(n_204), .B(n_482), .C(n_500), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_28), .A2(n_204), .B(n_482), .C(n_535), .Y(n_534) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_29), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_30), .B(n_206), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_31), .A2(n_477), .B(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_32), .B(n_206), .Y(n_247) );
INVx2_ASAP7_75t_L g163 ( .A(n_33), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_34), .A2(n_480), .B(n_484), .C(n_490), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_35), .B(n_165), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_36), .B(n_206), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_37), .B(n_224), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_39), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_40), .B(n_498), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_41), .Y(n_530) );
INVx1_ASAP7_75t_L g133 ( .A(n_42), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_43), .B(n_178), .Y(n_547) );
OAI22xp5_ASAP7_75t_SL g768 ( .A1(n_44), .A2(n_769), .B1(n_771), .B2(n_772), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_44), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_45), .B(n_477), .Y(n_533) );
OAI22xp5_ASAP7_75t_SL g138 ( .A1(n_46), .A2(n_139), .B1(n_140), .B2(n_461), .Y(n_138) );
INVx1_ASAP7_75t_L g461 ( .A(n_46), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g769 ( .A1(n_46), .A2(n_48), .B1(n_461), .B2(n_770), .Y(n_769) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_47), .A2(n_480), .B(n_490), .C(n_545), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_48), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_49), .B(n_165), .Y(n_188) );
INVx1_ASAP7_75t_L g515 ( .A(n_50), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_51), .A2(n_93), .B1(n_213), .B2(n_214), .Y(n_212) );
INVx1_ASAP7_75t_L g546 ( .A(n_52), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_53), .B(n_165), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_54), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_55), .B(n_477), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_56), .B(n_173), .Y(n_192) );
AOI22xp33_ASAP7_75t_SL g257 ( .A1(n_58), .A2(n_62), .B1(n_161), .B2(n_165), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_59), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_60), .B(n_165), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_61), .B(n_165), .Y(n_221) );
INVx1_ASAP7_75t_L g181 ( .A(n_63), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_64), .B(n_477), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_65), .B(n_509), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_66), .A2(n_167), .B(n_173), .C(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_67), .B(n_165), .Y(n_176) );
INVx1_ASAP7_75t_L g155 ( .A(n_68), .Y(n_155) );
OAI22xp33_ASAP7_75t_SL g765 ( .A1(n_69), .A2(n_766), .B1(n_773), .B2(n_774), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_69), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_70), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_71), .B(n_178), .Y(n_488) );
AO32x2_ASAP7_75t_L g210 ( .A1(n_72), .A2(n_185), .A3(n_204), .B1(n_211), .B2(n_216), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_73), .B(n_179), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_74), .A2(n_105), .B1(n_116), .B2(n_776), .Y(n_104) );
INVx1_ASAP7_75t_L g200 ( .A(n_75), .Y(n_200) );
INVx1_ASAP7_75t_L g242 ( .A(n_76), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_77), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_78), .B(n_487), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g579 ( .A1(n_79), .A2(n_482), .B(n_490), .C(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_80), .B(n_161), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g554 ( .A(n_81), .Y(n_554) );
INVx1_ASAP7_75t_L g115 ( .A(n_82), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_83), .B(n_486), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_85), .B(n_213), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_86), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_87), .B(n_161), .Y(n_246) );
INVx2_ASAP7_75t_L g153 ( .A(n_88), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_89), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_90), .B(n_203), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_91), .B(n_161), .Y(n_189) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_92), .B(n_112), .C(n_113), .Y(n_111) );
OR2x2_ASAP7_75t_L g124 ( .A(n_92), .B(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g464 ( .A(n_92), .B(n_126), .Y(n_464) );
INVx2_ASAP7_75t_L g468 ( .A(n_92), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_94), .A2(n_103), .B1(n_161), .B2(n_162), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_95), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g485 ( .A(n_96), .Y(n_485) );
INVxp67_ASAP7_75t_L g557 ( .A(n_97), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_98), .B(n_161), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_99), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g523 ( .A(n_100), .Y(n_523) );
INVx1_ASAP7_75t_L g581 ( .A(n_101), .Y(n_581) );
AND2x2_ASAP7_75t_L g548 ( .A(n_102), .B(n_206), .Y(n_548) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx5_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_108), .Y(n_777) );
OR2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND2x2_ASAP7_75t_L g126 ( .A(n_112), .B(n_127), .Y(n_126) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_129), .B1(n_761), .B2(n_764), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_122), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g763 ( .A(n_121), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_122), .A2(n_765), .B(n_775), .Y(n_764) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_128), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_124), .Y(n_775) );
NOR2x2_ASAP7_75t_L g760 ( .A(n_125), .B(n_468), .Y(n_760) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g467 ( .A(n_126), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g755 ( .A(n_130), .Y(n_755) );
CKINVDCx14_ASAP7_75t_R g134 ( .A(n_131), .Y(n_134) );
OAI22x1_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_462), .B1(n_465), .B2(n_469), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_138), .A2(n_462), .B1(n_467), .B2(n_757), .Y(n_756) );
OAI22xp5_ASAP7_75t_SL g766 ( .A1(n_139), .A2(n_140), .B1(n_767), .B2(n_768), .Y(n_766) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_141), .B(n_427), .Y(n_140) );
NOR3xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_331), .C(n_415), .Y(n_141) );
NAND4xp25_ASAP7_75t_L g142 ( .A(n_143), .B(n_274), .C(n_296), .D(n_312), .Y(n_142) );
AOI221xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_207), .B1(n_233), .B2(n_252), .C(n_260), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_183), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_146), .B(n_252), .Y(n_286) );
NAND4xp25_ASAP7_75t_L g326 ( .A(n_146), .B(n_314), .C(n_327), .D(n_329), .Y(n_326) );
INVxp67_ASAP7_75t_L g443 ( .A(n_146), .Y(n_443) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OR2x2_ASAP7_75t_L g325 ( .A(n_147), .B(n_263), .Y(n_325) );
AND2x2_ASAP7_75t_L g349 ( .A(n_147), .B(n_183), .Y(n_349) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g316 ( .A(n_148), .B(n_251), .Y(n_316) );
AND2x2_ASAP7_75t_L g356 ( .A(n_148), .B(n_337), .Y(n_356) );
AND2x2_ASAP7_75t_L g373 ( .A(n_148), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_148), .B(n_184), .Y(n_397) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g250 ( .A(n_149), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g268 ( .A(n_149), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g280 ( .A(n_149), .B(n_184), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_149), .B(n_194), .Y(n_302) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_157), .B(n_182), .Y(n_149) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_150), .A2(n_195), .B(n_205), .Y(n_194) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_151), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_153), .B(n_154), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
OAI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_171), .B(n_180), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_164), .C(n_167), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_160), .A2(n_527), .B(n_528), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_160), .A2(n_536), .B(n_537), .Y(n_535) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g166 ( .A(n_163), .Y(n_166) );
INVx1_ASAP7_75t_L g174 ( .A(n_163), .Y(n_174) );
INVx3_ASAP7_75t_L g241 ( .A(n_165), .Y(n_241) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_165), .Y(n_583) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_166), .Y(n_214) );
AND2x6_ASAP7_75t_L g482 ( .A(n_166), .B(n_483), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g580 ( .A1(n_167), .A2(n_581), .B(n_582), .C(n_583), .Y(n_580) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_168), .A2(n_245), .B(n_246), .Y(n_244) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g487 ( .A(n_169), .Y(n_487) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx3_ASAP7_75t_L g179 ( .A(n_170), .Y(n_179) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_170), .Y(n_203) );
INVx1_ASAP7_75t_L g224 ( .A(n_170), .Y(n_224) );
AND2x2_ASAP7_75t_L g478 ( .A(n_170), .B(n_174), .Y(n_478) );
INVx1_ASAP7_75t_L g483 ( .A(n_170), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_176), .C(n_177), .Y(n_171) );
O2A1O1Ixp5_ASAP7_75t_L g199 ( .A1(n_172), .A2(n_200), .B(n_201), .C(n_202), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_172), .A2(n_501), .B(n_502), .Y(n_500) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_177), .A2(n_191), .B(n_192), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_177), .A2(n_203), .B1(n_231), .B2(n_232), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_177), .A2(n_203), .B1(n_256), .B2(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_178), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_178), .A2(n_197), .B(n_198), .Y(n_196) );
O2A1O1Ixp5_ASAP7_75t_SL g240 ( .A1(n_178), .A2(n_241), .B(n_242), .C(n_243), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_178), .B(n_557), .Y(n_556) );
INVx5_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g211 ( .A1(n_179), .A2(n_203), .B1(n_212), .B2(n_215), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_180), .A2(n_187), .B(n_190), .Y(n_186) );
BUFx3_ASAP7_75t_L g204 ( .A(n_180), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_180), .A2(n_220), .B(n_225), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_180), .A2(n_240), .B(n_244), .Y(n_239) );
AND2x4_ASAP7_75t_L g477 ( .A(n_180), .B(n_478), .Y(n_477) );
INVx4_ASAP7_75t_SL g491 ( .A(n_180), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g524 ( .A(n_180), .B(n_478), .Y(n_524) );
AND2x2_ASAP7_75t_L g283 ( .A(n_183), .B(n_284), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_183), .A2(n_333), .B1(n_336), .B2(n_338), .C(n_342), .Y(n_332) );
AND2x2_ASAP7_75t_L g391 ( .A(n_183), .B(n_356), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_183), .B(n_373), .Y(n_425) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_194), .Y(n_183) );
INVx3_ASAP7_75t_L g251 ( .A(n_184), .Y(n_251) );
AND2x2_ASAP7_75t_L g300 ( .A(n_184), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g354 ( .A(n_184), .B(n_269), .Y(n_354) );
AND2x2_ASAP7_75t_L g412 ( .A(n_184), .B(n_413), .Y(n_412) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_193), .Y(n_184) );
INVx4_ASAP7_75t_L g254 ( .A(n_185), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_185), .A2(n_533), .B(n_534), .Y(n_532) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_185), .Y(n_551) );
AND2x2_ASAP7_75t_L g252 ( .A(n_194), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g269 ( .A(n_194), .Y(n_269) );
INVx1_ASAP7_75t_L g324 ( .A(n_194), .Y(n_324) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_194), .Y(n_330) );
AND2x2_ASAP7_75t_L g375 ( .A(n_194), .B(n_251), .Y(n_375) );
OR2x2_ASAP7_75t_L g414 ( .A(n_194), .B(n_253), .Y(n_414) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_199), .B(n_204), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_202), .A2(n_226), .B(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx4_ASAP7_75t_L g516 ( .A(n_203), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g273 ( .A(n_204), .B(n_254), .C(n_255), .Y(n_273) );
INVx2_ASAP7_75t_L g216 ( .A(n_206), .Y(n_216) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_206), .A2(n_219), .B(n_228), .Y(n_218) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_206), .A2(n_239), .B(n_247), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_206), .A2(n_476), .B(n_479), .Y(n_475) );
INVx1_ASAP7_75t_L g506 ( .A(n_206), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_206), .A2(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_207), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_217), .Y(n_207) );
AND2x2_ASAP7_75t_L g410 ( .A(n_208), .B(n_407), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_208), .B(n_392), .Y(n_442) );
BUFx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g341 ( .A(n_209), .B(n_265), .Y(n_341) );
AND2x2_ASAP7_75t_L g390 ( .A(n_209), .B(n_236), .Y(n_390) );
INVx1_ASAP7_75t_L g436 ( .A(n_209), .Y(n_436) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
AND2x2_ASAP7_75t_L g291 ( .A(n_210), .B(n_265), .Y(n_291) );
INVx1_ASAP7_75t_L g308 ( .A(n_210), .Y(n_308) );
AND2x2_ASAP7_75t_L g314 ( .A(n_210), .B(n_229), .Y(n_314) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_214), .Y(n_489) );
INVx2_ASAP7_75t_L g517 ( .A(n_214), .Y(n_517) );
INVx1_ASAP7_75t_L g503 ( .A(n_216), .Y(n_503) );
AND2x2_ASAP7_75t_L g382 ( .A(n_217), .B(n_290), .Y(n_382) );
INVx2_ASAP7_75t_L g447 ( .A(n_217), .Y(n_447) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_229), .Y(n_217) );
AND2x2_ASAP7_75t_L g264 ( .A(n_218), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g277 ( .A(n_218), .B(n_237), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_218), .B(n_236), .Y(n_305) );
INVx1_ASAP7_75t_L g311 ( .A(n_218), .Y(n_311) );
INVx1_ASAP7_75t_L g328 ( .A(n_218), .Y(n_328) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_218), .Y(n_340) );
INVx2_ASAP7_75t_L g408 ( .A(n_218), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g265 ( .A(n_229), .Y(n_265) );
BUFx2_ASAP7_75t_L g362 ( .A(n_229), .Y(n_362) );
AND2x2_ASAP7_75t_L g407 ( .A(n_229), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_248), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_235), .B(n_344), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_235), .A2(n_406), .B(n_420), .Y(n_430) );
AND2x2_ASAP7_75t_L g455 ( .A(n_235), .B(n_341), .Y(n_455) );
BUFx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g377 ( .A(n_237), .Y(n_377) );
AND2x2_ASAP7_75t_L g406 ( .A(n_237), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_238), .Y(n_290) );
INVx2_ASAP7_75t_L g309 ( .A(n_238), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_238), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g263 ( .A(n_249), .Y(n_263) );
OR2x2_ASAP7_75t_L g276 ( .A(n_249), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g344 ( .A(n_249), .B(n_340), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_249), .B(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g445 ( .A(n_249), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_249), .B(n_382), .Y(n_457) );
AND2x2_ASAP7_75t_L g336 ( .A(n_250), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g359 ( .A(n_250), .B(n_252), .Y(n_359) );
INVx2_ASAP7_75t_L g271 ( .A(n_251), .Y(n_271) );
AND2x2_ASAP7_75t_L g299 ( .A(n_251), .B(n_272), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_251), .B(n_324), .Y(n_380) );
AND2x2_ASAP7_75t_L g294 ( .A(n_252), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g441 ( .A(n_252), .Y(n_441) );
AND2x2_ASAP7_75t_L g453 ( .A(n_252), .B(n_316), .Y(n_453) );
AND2x2_ASAP7_75t_L g279 ( .A(n_253), .B(n_269), .Y(n_279) );
INVx1_ASAP7_75t_L g374 ( .A(n_253), .Y(n_374) );
AO21x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B(n_258), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_254), .B(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g509 ( .A(n_254), .Y(n_509) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_254), .A2(n_522), .B(n_529), .Y(n_521) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_254), .A2(n_578), .B(n_585), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_254), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g272 ( .A(n_259), .B(n_273), .Y(n_272) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_266), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_263), .B(n_310), .Y(n_319) );
OR2x2_ASAP7_75t_L g451 ( .A(n_263), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g368 ( .A(n_264), .B(n_309), .Y(n_368) );
AND2x2_ASAP7_75t_L g376 ( .A(n_264), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g435 ( .A(n_264), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g459 ( .A(n_264), .B(n_306), .Y(n_459) );
NOR2xp67_ASAP7_75t_L g417 ( .A(n_265), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g446 ( .A(n_265), .B(n_309), .Y(n_446) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2x1p5_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
AND2x2_ASAP7_75t_L g298 ( .A(n_268), .B(n_299), .Y(n_298) );
INVxp67_ASAP7_75t_L g460 ( .A(n_268), .Y(n_460) );
NOR2x1_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g295 ( .A(n_271), .Y(n_295) );
AND2x2_ASAP7_75t_L g346 ( .A(n_271), .B(n_279), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_271), .B(n_414), .Y(n_440) );
INVx2_ASAP7_75t_L g285 ( .A(n_272), .Y(n_285) );
INVx3_ASAP7_75t_L g337 ( .A(n_272), .Y(n_337) );
OR2x2_ASAP7_75t_L g365 ( .A(n_272), .B(n_366), .Y(n_365) );
AOI311xp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_278), .A3(n_280), .B(n_281), .C(n_292), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g312 ( .A1(n_275), .A2(n_313), .B(n_315), .C(n_317), .Y(n_312) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_SL g297 ( .A(n_277), .Y(n_297) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g315 ( .A(n_279), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_279), .B(n_295), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_279), .B(n_280), .Y(n_448) );
AND2x2_ASAP7_75t_L g370 ( .A(n_280), .B(n_284), .Y(n_370) );
AOI21xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_286), .B(n_287), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g428 ( .A(n_284), .B(n_316), .Y(n_428) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_285), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g322 ( .A(n_285), .Y(n_322) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
AND2x2_ASAP7_75t_L g313 ( .A(n_289), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g358 ( .A(n_291), .Y(n_358) );
AND2x4_ASAP7_75t_L g420 ( .A(n_291), .B(n_389), .Y(n_420) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI222xp33_ASAP7_75t_L g371 ( .A1(n_294), .A2(n_360), .B1(n_372), .B2(n_376), .C1(n_378), .C2(n_382), .Y(n_371) );
A2O1A1Ixp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B(n_300), .C(n_303), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_297), .B(n_341), .Y(n_364) );
INVx1_ASAP7_75t_L g386 ( .A(n_299), .Y(n_386) );
INVx1_ASAP7_75t_L g320 ( .A(n_301), .Y(n_320) );
OR2x2_ASAP7_75t_L g385 ( .A(n_302), .B(n_386), .Y(n_385) );
OAI21xp33_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_306), .B(n_310), .Y(n_303) );
NAND3xp33_ASAP7_75t_L g321 ( .A(n_304), .B(n_322), .C(n_323), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_304), .A2(n_341), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_308), .Y(n_361) );
AND2x2_ASAP7_75t_SL g327 ( .A(n_309), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g418 ( .A(n_309), .Y(n_418) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_309), .Y(n_434) );
INVx2_ASAP7_75t_L g392 ( .A(n_310), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_314), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g366 ( .A(n_316), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_320), .B1(n_321), .B2(n_325), .C(n_326), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_320), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g454 ( .A(n_320), .Y(n_454) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g335 ( .A(n_327), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_327), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g393 ( .A(n_327), .B(n_341), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_327), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g426 ( .A(n_327), .B(n_361), .Y(n_426) );
BUFx3_ASAP7_75t_L g389 ( .A(n_328), .Y(n_389) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND5xp2_ASAP7_75t_L g331 ( .A(n_332), .B(n_350), .C(n_371), .D(n_383), .E(n_398), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AOI32xp33_ASAP7_75t_L g423 ( .A1(n_335), .A2(n_362), .A3(n_378), .B1(n_424), .B2(n_426), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_337), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_SL g347 ( .A(n_341), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_345), .B1(n_347), .B2(n_348), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_357), .B1(n_359), .B2(n_360), .C(n_363), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g422 ( .A(n_354), .B(n_373), .Y(n_422) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_359), .A2(n_420), .B1(n_438), .B2(n_443), .C(n_444), .Y(n_437) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx2_ASAP7_75t_L g403 ( .A(n_362), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_367), .B2(n_369), .Y(n_363) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_L g381 ( .A(n_373), .Y(n_381) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
AOI222xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_387), .B1(n_391), .B2(n_392), .C1(n_393), .C2(n_394), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g438 ( .A1(n_392), .A2(n_439), .B1(n_441), .B2(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_409), .B(n_411), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g452 ( .A(n_407), .Y(n_452) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
A2O1A1Ixp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_419), .B(n_421), .C(n_423), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI211xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B(n_431), .C(n_456), .Y(n_427) );
CKINVDCx16_ASAP7_75t_R g432 ( .A(n_428), .Y(n_432) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI211xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B(n_437), .C(n_449), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_447), .B(n_448), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_453), .B1(n_454), .B2(n_455), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AOI21xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B(n_460), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g757 ( .A(n_469), .Y(n_757) );
OR3x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_669), .C(n_712), .Y(n_469) );
NAND5xp2_ASAP7_75t_L g470 ( .A(n_471), .B(n_596), .C(n_626), .D(n_643), .E(n_658), .Y(n_470) );
AOI221xp5_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_519), .B1(n_559), .B2(n_565), .C(n_569), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_494), .Y(n_472) );
OR2x2_ASAP7_75t_L g574 ( .A(n_473), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g613 ( .A(n_473), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g631 ( .A(n_473), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_473), .B(n_567), .Y(n_648) );
OR2x2_ASAP7_75t_L g660 ( .A(n_473), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_473), .B(n_619), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_473), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_473), .B(n_597), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_473), .B(n_605), .Y(n_711) );
AND2x2_ASAP7_75t_L g743 ( .A(n_473), .B(n_507), .Y(n_743) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_473), .Y(n_751) );
INVx5_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_474), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g571 ( .A(n_474), .B(n_549), .Y(n_571) );
BUFx2_ASAP7_75t_L g593 ( .A(n_474), .Y(n_593) );
AND2x2_ASAP7_75t_L g622 ( .A(n_474), .B(n_495), .Y(n_622) );
AND2x2_ASAP7_75t_L g677 ( .A(n_474), .B(n_575), .Y(n_677) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_492), .Y(n_474) );
BUFx2_ASAP7_75t_L g498 ( .A(n_477), .Y(n_498) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g511 ( .A1(n_481), .A2(n_491), .B(n_512), .C(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g553 ( .A1(n_481), .A2(n_491), .B(n_554), .C(n_555), .Y(n_553) );
INVx5_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_488), .C(n_489), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_486), .A2(n_489), .B(n_546), .C(n_547), .Y(n_545) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_494), .B(n_631), .Y(n_640) );
OAI32xp33_ASAP7_75t_L g654 ( .A1(n_494), .A2(n_590), .A3(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_494), .B(n_656), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_494), .B(n_574), .Y(n_697) );
INVx1_ASAP7_75t_SL g726 ( .A(n_494), .Y(n_726) );
NAND4xp25_ASAP7_75t_L g735 ( .A(n_494), .B(n_521), .C(n_677), .D(n_736), .Y(n_735) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_507), .Y(n_494) );
INVx5_ASAP7_75t_L g568 ( .A(n_495), .Y(n_568) );
AND2x2_ASAP7_75t_L g597 ( .A(n_495), .B(n_508), .Y(n_597) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_495), .Y(n_676) );
AND2x2_ASAP7_75t_L g746 ( .A(n_495), .B(n_693), .Y(n_746) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_504), .Y(n_495) );
AOI21xp5_ASAP7_75t_SL g496 ( .A1(n_497), .A2(n_499), .B(n_503), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x4_ASAP7_75t_L g619 ( .A(n_507), .B(n_568), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_507), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g653 ( .A(n_507), .B(n_575), .Y(n_653) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g567 ( .A(n_508), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g605 ( .A(n_508), .B(n_577), .Y(n_605) );
AND2x2_ASAP7_75t_L g614 ( .A(n_508), .B(n_576), .Y(n_614) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_518), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
AOI222xp33_ASAP7_75t_L g682 ( .A1(n_519), .A2(n_683), .B1(n_685), .B2(n_687), .C1(n_690), .C2(n_691), .Y(n_682) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_538), .Y(n_519) );
AND2x2_ASAP7_75t_L g615 ( .A(n_520), .B(n_616), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g732 ( .A(n_520), .B(n_593), .C(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_531), .Y(n_520) );
INVx5_ASAP7_75t_SL g564 ( .A(n_521), .Y(n_564) );
OAI322xp33_ASAP7_75t_L g569 ( .A1(n_521), .A2(n_570), .A3(n_572), .B1(n_573), .B2(n_587), .C1(n_590), .C2(n_592), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_521), .B(n_562), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_521), .B(n_550), .Y(n_741) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_525), .Y(n_522) );
INVx2_ASAP7_75t_L g562 ( .A(n_531), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_531), .B(n_540), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_538), .B(n_600), .Y(n_655) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g634 ( .A(n_539), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_549), .Y(n_539) );
OR2x2_ASAP7_75t_L g563 ( .A(n_540), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_540), .B(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g602 ( .A(n_540), .B(n_550), .Y(n_602) );
AND2x2_ASAP7_75t_L g625 ( .A(n_540), .B(n_562), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_540), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g641 ( .A(n_540), .B(n_600), .Y(n_641) );
AND2x2_ASAP7_75t_L g649 ( .A(n_540), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_540), .B(n_609), .Y(n_699) );
INVx5_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g589 ( .A(n_541), .B(n_564), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_541), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g616 ( .A(n_541), .B(n_550), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_541), .B(n_663), .Y(n_704) );
OR2x2_ASAP7_75t_L g720 ( .A(n_541), .B(n_664), .Y(n_720) );
AND2x2_ASAP7_75t_SL g727 ( .A(n_541), .B(n_681), .Y(n_727) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_541), .Y(n_734) );
OR2x6_ASAP7_75t_L g541 ( .A(n_542), .B(n_548), .Y(n_541) );
AND2x2_ASAP7_75t_L g588 ( .A(n_549), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g638 ( .A(n_549), .B(n_562), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_549), .B(n_564), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_549), .B(n_600), .Y(n_722) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_550), .B(n_564), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_550), .B(n_562), .Y(n_610) );
OR2x2_ASAP7_75t_L g664 ( .A(n_550), .B(n_562), .Y(n_664) );
AND2x2_ASAP7_75t_L g681 ( .A(n_550), .B(n_561), .Y(n_681) );
INVxp67_ASAP7_75t_L g703 ( .A(n_550), .Y(n_703) );
AND2x2_ASAP7_75t_L g730 ( .A(n_550), .B(n_600), .Y(n_730) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_550), .Y(n_737) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_552), .B(n_558), .Y(n_550) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_561), .B(n_611), .Y(n_684) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g600 ( .A(n_562), .B(n_564), .Y(n_600) );
OR2x2_ASAP7_75t_L g667 ( .A(n_562), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g611 ( .A(n_563), .Y(n_611) );
OR2x2_ASAP7_75t_L g672 ( .A(n_563), .B(n_664), .Y(n_672) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g572 ( .A(n_567), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_567), .B(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g573 ( .A(n_568), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_568), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_568), .B(n_575), .Y(n_607) );
INVx2_ASAP7_75t_L g652 ( .A(n_568), .Y(n_652) );
AND2x2_ASAP7_75t_L g665 ( .A(n_568), .B(n_605), .Y(n_665) );
AND2x2_ASAP7_75t_L g690 ( .A(n_568), .B(n_614), .Y(n_690) );
INVx1_ASAP7_75t_L g642 ( .A(n_573), .Y(n_642) );
INVx2_ASAP7_75t_SL g629 ( .A(n_574), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_575), .Y(n_632) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_576), .Y(n_595) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
BUFx2_ASAP7_75t_L g693 ( .A(n_577), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_584), .Y(n_578) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g662 ( .A(n_589), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g668 ( .A(n_589), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_589), .A2(n_671), .B1(n_673), .B2(n_678), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_589), .B(n_681), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_590), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g624 ( .A(n_591), .Y(n_624) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OR2x2_ASAP7_75t_L g606 ( .A(n_593), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_593), .B(n_597), .Y(n_657) );
AND2x2_ASAP7_75t_L g680 ( .A(n_593), .B(n_681), .Y(n_680) );
BUFx2_ASAP7_75t_L g656 ( .A(n_595), .Y(n_656) );
AOI211xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_603), .C(n_617), .Y(n_596) );
INVx1_ASAP7_75t_L g620 ( .A(n_597), .Y(n_620) );
OAI221xp5_ASAP7_75t_SL g728 ( .A1(n_597), .A2(n_729), .B1(n_731), .B2(n_732), .C(n_735), .Y(n_728) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g747 ( .A(n_600), .Y(n_747) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g696 ( .A(n_602), .B(n_635), .Y(n_696) );
A2O1A1Ixp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_606), .B(n_608), .C(n_612), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
OAI32xp33_ASAP7_75t_L g721 ( .A1(n_610), .A2(n_611), .A3(n_674), .B1(n_711), .B2(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
AND2x2_ASAP7_75t_L g753 ( .A(n_613), .B(n_652), .Y(n_753) );
AND2x2_ASAP7_75t_L g700 ( .A(n_614), .B(n_652), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_614), .B(n_622), .Y(n_718) );
AOI31xp33_ASAP7_75t_SL g617 ( .A1(n_618), .A2(n_620), .A3(n_621), .B(n_623), .Y(n_617) );
INVxp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_619), .B(n_631), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_619), .B(n_629), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g738 ( .A1(n_619), .A2(n_649), .B1(n_739), .B2(n_742), .C(n_744), .Y(n_738) );
CKINVDCx16_ASAP7_75t_R g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
AND2x2_ASAP7_75t_L g644 ( .A(n_624), .B(n_645), .Y(n_644) );
AOI222xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_633), .B1(n_636), .B2(n_639), .C1(n_641), .C2(n_642), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g709 ( .A(n_628), .Y(n_709) );
INVx1_ASAP7_75t_L g731 ( .A(n_631), .Y(n_731) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_634), .A2(n_745), .B1(n_747), .B2(n_748), .Y(n_744) );
INVx1_ASAP7_75t_L g650 ( .A(n_635), .Y(n_650) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_647), .B1(n_649), .B2(n_651), .C(n_654), .Y(n_643) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g688 ( .A(n_646), .B(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g740 ( .A(n_646), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g715 ( .A(n_651), .Y(n_715) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g679 ( .A(n_652), .Y(n_679) );
INVx1_ASAP7_75t_L g661 ( .A(n_653), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_656), .B(n_743), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .B1(n_665), .B2(n_666), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g752 ( .A(n_665), .Y(n_752) );
INVxp33_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_667), .B(n_711), .Y(n_710) );
OAI32xp33_ASAP7_75t_L g701 ( .A1(n_668), .A2(n_702), .A3(n_703), .B1(n_704), .B2(n_705), .Y(n_701) );
NAND4xp25_ASAP7_75t_L g669 ( .A(n_670), .B(n_682), .C(n_694), .D(n_706), .Y(n_669) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
NAND2xp33_ASAP7_75t_SL g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_677), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
CKINVDCx16_ASAP7_75t_R g687 ( .A(n_688), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_691), .A2(n_707), .B1(n_724), .B2(n_727), .C(n_728), .Y(n_723) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g742 ( .A(n_693), .B(n_743), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_697), .B1(n_698), .B2(n_700), .C(n_701), .Y(n_694) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_703), .B(n_734), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B(n_710), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND4xp25_ASAP7_75t_L g712 ( .A(n_713), .B(n_723), .C(n_738), .D(n_749), .Y(n_712) );
O2A1O1Ixp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_717), .B(n_719), .C(n_721), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g754 ( .A(n_741), .Y(n_754) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_753), .B(n_754), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
BUFx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g774 ( .A(n_766), .Y(n_774) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_769), .Y(n_772) );
INVx1_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
endmodule