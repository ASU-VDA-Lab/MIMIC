module fake_jpeg_11362_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_10),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_62),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_1),
.B(n_2),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_44),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_3),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_44),
.B1(n_43),
.B2(n_45),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_74),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_57),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_45),
.B1(n_52),
.B2(n_51),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_50),
.B1(n_49),
.B2(n_47),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_58),
.B1(n_42),
.B2(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_3),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_88),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_99),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_93),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_92),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_98),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_72),
.A2(n_55),
.B1(n_41),
.B2(n_6),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_12),
.B(n_15),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_41),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_4),
.Y(n_98)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_108),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_41),
.B1(n_6),
.B2(n_7),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_5),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_5),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_8),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_114),
.C(n_116),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_8),
.B(n_9),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_116),
.C(n_109),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_10),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_37),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_117),
.B(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_130),
.B1(n_118),
.B2(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_125),
.B(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_125),
.B1(n_122),
.B2(n_123),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_134),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_132),
.C(n_133),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.C(n_104),
.Y(n_141)
);

OAI31xp33_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_127),
.A3(n_137),
.B(n_101),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_127),
.A3(n_102),
.B1(n_104),
.B2(n_107),
.C1(n_26),
.C2(n_27),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_23),
.B(n_30),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_32),
.Y(n_146)
);


endmodule