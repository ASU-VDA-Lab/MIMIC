module fake_jpeg_7292_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_31;
wire n_25;
wire n_17;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx6_ASAP7_75t_SL g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx4f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_19),
.A2(n_22),
.B1(n_13),
.B2(n_14),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_18),
.B(n_1),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_15),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_20),
.B(n_22),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_33),
.C(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_34),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_10),
.B(n_23),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_10),
.B(n_12),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_10),
.Y(n_37)
);

AND2x6_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_39),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_30),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_10),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_14),
.B1(n_11),
.B2(n_16),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_17),
.B1(n_16),
.B2(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_47),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_53),
.Y(n_60)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_37),
.C(n_36),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_44),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_53),
.C(n_55),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_41),
.B1(n_48),
.B2(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_24),
.B1(n_12),
.B2(n_6),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_51),
.B1(n_57),
.B2(n_12),
.Y(n_64)
);

NOR3xp33_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_51),
.C(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_63),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_59),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_60),
.B(n_24),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_59),
.B1(n_57),
.B2(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_3),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_70),
.B(n_67),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_71),
.A2(n_72),
.B(n_5),
.Y(n_73)
);

OA21x2_ASAP7_75t_SL g72 ( 
.A1(n_70),
.A2(n_68),
.B(n_7),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_5),
.Y(n_74)
);


endmodule