module fake_netlist_6_4551_n_804 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_804);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_804;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_760;
wire n_741;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_683;
wire n_420;
wire n_620;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_787;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_44),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_18),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_2),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_89),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_50),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_42),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_7),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_14),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_122),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_99),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_90),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_51),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_65),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_105),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_57),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_113),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_94),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_76),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_46),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_108),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_21),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_141),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_20),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_78),
.Y(n_192)
);

NOR2xp67_ASAP7_75t_L g193 ( 
.A(n_80),
.B(n_109),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_137),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_29),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_14),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_77),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_70),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_126),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_0),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_33),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_48),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_5),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_45),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_112),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_L g210 ( 
.A(n_49),
.B(n_102),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_95),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_132),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_135),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_24),
.Y(n_215)
);

CKINVDCx11_ASAP7_75t_R g216 ( 
.A(n_169),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_159),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_159),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_22),
.Y(n_223)
);

AND2x4_ASAP7_75t_SL g224 ( 
.A(n_194),
.B(n_23),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_25),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_173),
.B(n_0),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

OA21x2_ASAP7_75t_L g232 ( 
.A1(n_196),
.A2(n_1),
.B(n_2),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_26),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_173),
.B(n_187),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_161),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_1),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_167),
.B(n_27),
.Y(n_245)
);

BUFx8_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_190),
.B(n_3),
.Y(n_249)
);

BUFx8_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_162),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_170),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_184),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_205),
.B(n_3),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_189),
.Y(n_259)
);

NOR2x1p5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_206),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_220),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_194),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_217),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_164),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_169),
.B1(n_207),
.B2(n_200),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_217),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_223),
.B(n_227),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_220),
.B(n_160),
.Y(n_278)
);

CKINVDCx6p67_ASAP7_75t_R g279 ( 
.A(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_216),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_226),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_253),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_230),
.B(n_191),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

OR2x6_ASAP7_75t_L g286 ( 
.A(n_242),
.B(n_193),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_223),
.B(n_199),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_SL g288 ( 
.A(n_249),
.B(n_197),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_218),
.B(n_165),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_258),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_223),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_251),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_252),
.A2(n_227),
.B1(n_233),
.B2(n_245),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_217),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_245),
.B(n_197),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_218),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_245),
.B(n_227),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_236),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_222),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_233),
.B(n_200),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_222),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_222),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_222),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_222),
.Y(n_307)
);

AND3x2_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_204),
.C(n_208),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_278),
.Y(n_309)
);

BUFx5_ASAP7_75t_L g310 ( 
.A(n_290),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_262),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_233),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

NAND2xp33_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_257),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_267),
.B(n_224),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_168),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_224),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_218),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_269),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_290),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_228),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_246),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_171),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_246),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_228),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_260),
.A2(n_232),
.B1(n_234),
.B2(n_238),
.Y(n_327)
);

BUFx6f_ASAP7_75t_SL g328 ( 
.A(n_286),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_291),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_228),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_299),
.B(n_237),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_246),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_263),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_273),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_293),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_292),
.B(n_250),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_287),
.B(n_250),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_271),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_240),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_279),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_270),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_288),
.A2(n_215),
.B1(n_174),
.B2(n_175),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_273),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_274),
.B(n_275),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_288),
.B(n_172),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_274),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_L g349 ( 
.A(n_282),
.B(n_219),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_L g350 ( 
.A(n_268),
.B(n_229),
.C(n_243),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_275),
.B(n_250),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_284),
.B(n_231),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_284),
.B(n_231),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_286),
.A2(n_232),
.B1(n_234),
.B2(n_259),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_285),
.B(n_231),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_286),
.B(n_276),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_L g357 ( 
.A(n_285),
.B(n_176),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_266),
.B(n_219),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_308),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_266),
.B(n_219),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_266),
.B(n_219),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_276),
.B(n_210),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_304),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_282),
.B(n_219),
.Y(n_364)
);

O2A1O1Ixp33_ASAP7_75t_L g365 ( 
.A1(n_281),
.A2(n_232),
.B(n_234),
.C(n_203),
.Y(n_365)
);

BUFx6f_ASAP7_75t_SL g366 ( 
.A(n_279),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_304),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_294),
.B(n_221),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_294),
.B(n_221),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_281),
.B(n_177),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_294),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_307),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_293),
.B(n_255),
.Y(n_373)
);

NAND3xp33_ASAP7_75t_L g374 ( 
.A(n_297),
.B(n_214),
.C(n_183),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_315),
.Y(n_375)
);

AOI21x1_ASAP7_75t_L g376 ( 
.A1(n_352),
.A2(n_307),
.B(n_306),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_312),
.A2(n_221),
.B(n_277),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_318),
.B(n_179),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_326),
.A2(n_186),
.B1(n_192),
.B2(n_195),
.Y(n_379)
);

A2O1A1Ixp33_ASAP7_75t_L g380 ( 
.A1(n_365),
.A2(n_297),
.B(n_261),
.C(n_264),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_327),
.B(n_354),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_313),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_322),
.B(n_327),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_319),
.B(n_216),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_340),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_316),
.B(n_280),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_365),
.A2(n_261),
.B(n_264),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_311),
.Y(n_388)
);

BUFx12f_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_319),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_314),
.A2(n_221),
.B(n_277),
.Y(n_391)
);

NOR2x2_ASAP7_75t_L g392 ( 
.A(n_328),
.B(n_4),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_209),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_320),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_353),
.A2(n_221),
.B(n_277),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_355),
.A2(n_277),
.B(n_271),
.Y(n_396)
);

AOI21x1_ASAP7_75t_L g397 ( 
.A1(n_346),
.A2(n_306),
.B(n_305),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_336),
.B(n_302),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_341),
.A2(n_212),
.B1(n_302),
.B2(n_296),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_309),
.Y(n_400)
);

A2O1A1Ixp33_ASAP7_75t_L g401 ( 
.A1(n_354),
.A2(n_305),
.B(n_296),
.C(n_302),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_356),
.B(n_4),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_336),
.A2(n_255),
.B(n_248),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_344),
.A2(n_255),
.B1(n_241),
.B2(n_247),
.Y(n_404)
);

CKINVDCx10_ASAP7_75t_R g405 ( 
.A(n_366),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_356),
.B(n_255),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_349),
.B(n_255),
.Y(n_407)
);

O2A1O1Ixp33_ASAP7_75t_L g408 ( 
.A1(n_350),
.A2(n_225),
.B(n_241),
.C(n_247),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_364),
.B(n_225),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_332),
.B(n_225),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_331),
.A2(n_248),
.B(n_247),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_321),
.Y(n_412)
);

AND2x4_ASAP7_75t_SL g413 ( 
.A(n_359),
.B(n_271),
.Y(n_413)
);

AOI33xp33_ASAP7_75t_L g414 ( 
.A1(n_362),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.B3(n_9),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_362),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_331),
.B(n_350),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_335),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_323),
.A2(n_277),
.B(n_271),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_310),
.B(n_329),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_325),
.B(n_271),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_347),
.B(n_28),
.Y(n_421)
);

AOI21x1_ASAP7_75t_L g422 ( 
.A1(n_358),
.A2(n_248),
.B(n_247),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_330),
.B(n_225),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_351),
.A2(n_248),
.B(n_247),
.Y(n_424)
);

AO21x1_ASAP7_75t_L g425 ( 
.A1(n_317),
.A2(n_6),
.B(n_8),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_333),
.A2(n_248),
.B(n_241),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_338),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_334),
.B(n_225),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_337),
.A2(n_241),
.B(n_82),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_343),
.B(n_241),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_357),
.A2(n_81),
.B(n_155),
.Y(n_431)
);

A2O1A1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_324),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_370),
.B(n_10),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_360),
.A2(n_83),
.B(n_154),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_L g435 ( 
.A1(n_363),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_371),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_367),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_361),
.A2(n_79),
.B(n_153),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_345),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_374),
.B(n_12),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_372),
.B(n_30),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_348),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_328),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_416),
.A2(n_310),
.B1(n_339),
.B2(n_373),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_381),
.B(n_310),
.Y(n_446)
);

O2A1O1Ixp5_ASAP7_75t_L g447 ( 
.A1(n_397),
.A2(n_339),
.B(n_373),
.C(n_368),
.Y(n_447)
);

OAI21xp33_ASAP7_75t_L g448 ( 
.A1(n_393),
.A2(n_366),
.B(n_369),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_381),
.B(n_310),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_385),
.A2(n_433),
.B(n_402),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_390),
.B(n_31),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_384),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_383),
.B(n_310),
.Y(n_453)
);

AO221x2_ASAP7_75t_L g454 ( 
.A1(n_443),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_454)
);

AOI21x1_ASAP7_75t_L g455 ( 
.A1(n_376),
.A2(n_310),
.B(n_87),
.Y(n_455)
);

OR2x6_ASAP7_75t_L g456 ( 
.A(n_389),
.B(n_388),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_417),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_390),
.B(n_17),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_421),
.A2(n_88),
.B1(n_32),
.B2(n_34),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_412),
.B(n_19),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_400),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

OA21x2_ASAP7_75t_L g463 ( 
.A1(n_387),
.A2(n_91),
.B(n_35),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_415),
.Y(n_464)
);

OR2x6_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_19),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_421),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_420),
.A2(n_39),
.B(n_40),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_418),
.A2(n_419),
.B(n_396),
.Y(n_468)
);

A2O1A1Ixp33_ASAP7_75t_L g469 ( 
.A1(n_375),
.A2(n_41),
.B(n_43),
.C(n_47),
.Y(n_469)
);

BUFx12f_ASAP7_75t_L g470 ( 
.A(n_427),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_386),
.B(n_52),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_419),
.A2(n_156),
.B(n_54),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_398),
.B(n_53),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_377),
.A2(n_55),
.B(n_56),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_413),
.B(n_58),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_394),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_440),
.Y(n_477)
);

OAI21x1_ASAP7_75t_L g478 ( 
.A1(n_422),
.A2(n_152),
.B(n_60),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_394),
.Y(n_479)
);

BUFx12f_ASAP7_75t_L g480 ( 
.A(n_436),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_442),
.B(n_59),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_378),
.B(n_61),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_401),
.A2(n_62),
.B(n_63),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_439),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_379),
.Y(n_485)
);

AO21x2_ASAP7_75t_L g486 ( 
.A1(n_387),
.A2(n_149),
.B(n_66),
.Y(n_486)
);

AO31x2_ASAP7_75t_L g487 ( 
.A1(n_380),
.A2(n_425),
.A3(n_432),
.B(n_435),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_391),
.A2(n_148),
.B(n_67),
.Y(n_488)
);

A2O1A1Ixp33_ASAP7_75t_L g489 ( 
.A1(n_399),
.A2(n_64),
.B(n_68),
.C(n_69),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_439),
.B(n_71),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_441),
.A2(n_72),
.B(n_73),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_406),
.A2(n_411),
.B(n_410),
.Y(n_492)
);

AOI221xp5_ASAP7_75t_L g493 ( 
.A1(n_408),
.A2(n_74),
.B1(n_75),
.B2(n_84),
.C(n_85),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_403),
.B(n_86),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_423),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_428),
.A2(n_92),
.B(n_93),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

A2O1A1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_411),
.A2(n_96),
.B(n_97),
.C(n_100),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_429),
.B(n_101),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_403),
.B(n_430),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_426),
.B(n_104),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_474),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_462),
.Y(n_503)
);

AOI22x1_ASAP7_75t_L g504 ( 
.A1(n_492),
.A2(n_431),
.B1(n_434),
.B2(n_438),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_468),
.A2(n_424),
.B(n_395),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_461),
.Y(n_506)
);

NAND3xp33_ASAP7_75t_L g507 ( 
.A(n_450),
.B(n_404),
.C(n_409),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_445),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_407),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_455),
.A2(n_404),
.B(n_110),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_447),
.A2(n_107),
.B(n_114),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_445),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_488),
.A2(n_115),
.B(n_116),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_457),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_478),
.A2(n_117),
.B(n_118),
.Y(n_515)
);

AO21x2_ASAP7_75t_L g516 ( 
.A1(n_473),
.A2(n_120),
.B(n_121),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_483),
.A2(n_123),
.B(n_125),
.Y(n_517)
);

BUFx6f_ASAP7_75t_SL g518 ( 
.A(n_456),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_472),
.A2(n_496),
.B(n_449),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_446),
.A2(n_128),
.B(n_131),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_470),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_457),
.Y(n_522)
);

BUFx4f_ASAP7_75t_SL g523 ( 
.A(n_480),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_479),
.Y(n_524)
);

AO21x2_ASAP7_75t_L g525 ( 
.A1(n_500),
.A2(n_134),
.B(n_138),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_464),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_453),
.A2(n_139),
.B(n_140),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_490),
.A2(n_142),
.B(n_143),
.Y(n_528)
);

CKINVDCx8_ASAP7_75t_R g529 ( 
.A(n_456),
.Y(n_529)
);

BUFx2_ASAP7_75t_SL g530 ( 
.A(n_464),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_452),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_495),
.A2(n_144),
.B(n_145),
.Y(n_532)
);

AO21x2_ASAP7_75t_L g533 ( 
.A1(n_444),
.A2(n_146),
.B(n_147),
.Y(n_533)
);

OA21x2_ASAP7_75t_L g534 ( 
.A1(n_495),
.A2(n_392),
.B(n_405),
.Y(n_534)
);

AO21x2_ASAP7_75t_L g535 ( 
.A1(n_458),
.A2(n_494),
.B(n_451),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_485),
.A2(n_482),
.B(n_451),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_498),
.A2(n_477),
.B(n_460),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_476),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_497),
.B(n_484),
.Y(n_539)
);

AO21x2_ASAP7_75t_L g540 ( 
.A1(n_486),
.A2(n_489),
.B(n_481),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_501),
.A2(n_463),
.B(n_467),
.Y(n_541)
);

NAND2x1p5_ASAP7_75t_L g542 ( 
.A(n_475),
.B(n_464),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_499),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_499),
.Y(n_544)
);

AO21x2_ASAP7_75t_L g545 ( 
.A1(n_486),
.A2(n_448),
.B(n_469),
.Y(n_545)
);

BUFx4f_ASAP7_75t_SL g546 ( 
.A(n_471),
.Y(n_546)
);

OAI21x1_ASAP7_75t_SL g547 ( 
.A1(n_466),
.A2(n_459),
.B(n_463),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_497),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_497),
.Y(n_549)
);

BUFx4_ASAP7_75t_SL g550 ( 
.A(n_465),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_505),
.A2(n_491),
.B(n_493),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_508),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_L g553 ( 
.A1(n_546),
.A2(n_465),
.B1(n_454),
.B2(n_487),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_512),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_544),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_537),
.B(n_487),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_514),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_522),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_524),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_526),
.B(n_487),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_506),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_503),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_524),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_550),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_538),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_543),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_539),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_506),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_531),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_544),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_548),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_544),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_549),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_543),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_548),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_543),
.Y(n_576)
);

CKINVDCx8_ASAP7_75t_R g577 ( 
.A(n_530),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_521),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_543),
.Y(n_579)
);

OAI21x1_ASAP7_75t_L g580 ( 
.A1(n_505),
.A2(n_454),
.B(n_519),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_548),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_536),
.B(n_507),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_548),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_509),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_509),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_529),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_542),
.Y(n_587)
);

AO21x2_ASAP7_75t_L g588 ( 
.A1(n_547),
.A2(n_519),
.B(n_540),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_543),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_546),
.B(n_542),
.Y(n_590)
);

AO21x1_ASAP7_75t_SL g591 ( 
.A1(n_533),
.A2(n_545),
.B(n_532),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_517),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_526),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_533),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_511),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_567),
.B(n_526),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_567),
.B(n_534),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_569),
.Y(n_598)
);

NAND2x1_ASAP7_75t_L g599 ( 
.A(n_555),
.B(n_502),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_556),
.B(n_545),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_556),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_561),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_563),
.B(n_533),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_552),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_582),
.B(n_534),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_559),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_568),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_554),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_566),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_559),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_582),
.B(n_540),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_580),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_580),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_560),
.B(n_527),
.Y(n_614)
);

INVxp67_ASAP7_75t_R g615 ( 
.A(n_571),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_560),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_560),
.B(n_527),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_568),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_577),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_566),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_557),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_558),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_562),
.B(n_525),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_587),
.B(n_513),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_562),
.B(n_525),
.Y(n_625)
);

AND2x4_ASAP7_75t_SL g626 ( 
.A(n_566),
.B(n_502),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_590),
.B(n_534),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_570),
.B(n_516),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_570),
.B(n_516),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_SL g630 ( 
.A1(n_586),
.A2(n_518),
.B1(n_523),
.B2(n_504),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_565),
.Y(n_631)
);

NOR2x1_ASAP7_75t_R g632 ( 
.A(n_564),
.B(n_523),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_584),
.B(n_513),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_572),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_572),
.B(n_520),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_594),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_566),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_565),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_594),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_553),
.A2(n_518),
.B1(n_535),
.B2(n_517),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_586),
.B(n_529),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_555),
.B(n_520),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_555),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_585),
.A2(n_518),
.B1(n_535),
.B2(n_502),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_574),
.B(n_532),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_588),
.B(n_535),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_621),
.Y(n_647)
);

NAND3xp33_ASAP7_75t_L g648 ( 
.A(n_605),
.B(n_578),
.C(n_573),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_627),
.B(n_583),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_621),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_597),
.B(n_598),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_601),
.B(n_588),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_638),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_601),
.B(n_575),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_618),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_616),
.B(n_611),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_634),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_631),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_618),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_602),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_638),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_596),
.B(n_581),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_636),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_636),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_616),
.B(n_593),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_641),
.A2(n_564),
.B1(n_574),
.B2(n_589),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_630),
.A2(n_588),
.B1(n_591),
.B2(n_589),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_609),
.B(n_576),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_611),
.B(n_603),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_639),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_639),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_606),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_604),
.B(n_576),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_606),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_608),
.B(n_592),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_603),
.B(n_591),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_619),
.A2(n_579),
.B1(n_566),
.B2(n_592),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_640),
.A2(n_551),
.B1(n_579),
.B2(n_592),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_622),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_609),
.B(n_579),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_623),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_610),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_607),
.B(n_577),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_607),
.B(n_610),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_634),
.B(n_528),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_643),
.B(n_579),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_623),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_664),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_663),
.B(n_613),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_655),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_651),
.B(n_600),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_669),
.B(n_600),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_670),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_669),
.B(n_656),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_649),
.B(n_625),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_681),
.B(n_646),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_663),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_656),
.B(n_617),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_687),
.B(n_613),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_681),
.B(n_617),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_660),
.B(n_625),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_652),
.B(n_646),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_671),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_647),
.Y(n_704)
);

OA21x2_ASAP7_75t_L g705 ( 
.A1(n_678),
.A2(n_612),
.B(n_595),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_650),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_658),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_662),
.B(n_643),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_665),
.B(n_644),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_679),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_676),
.B(n_614),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_676),
.B(n_614),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_653),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_648),
.B(n_666),
.C(n_678),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_652),
.B(n_612),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_683),
.A2(n_615),
.B1(n_609),
.B2(n_620),
.Y(n_716)
);

NAND2x1p5_ASAP7_75t_L g717 ( 
.A(n_655),
.B(n_599),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_683),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_702),
.B(n_675),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_697),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_690),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_707),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_702),
.B(n_657),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_691),
.B(n_659),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_710),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_704),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_692),
.B(n_659),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_692),
.B(n_653),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_690),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_694),
.B(n_685),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_706),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_688),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_713),
.Y(n_733)
);

OAI211xp5_ASAP7_75t_L g734 ( 
.A1(n_714),
.A2(n_667),
.B(n_677),
.C(n_684),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_694),
.B(n_661),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_696),
.B(n_654),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_698),
.B(n_667),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_693),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_696),
.B(n_673),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_703),
.Y(n_740)
);

NAND2x1_ASAP7_75t_SL g741 ( 
.A(n_733),
.B(n_715),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_726),
.Y(n_742)
);

OAI21xp33_ASAP7_75t_L g743 ( 
.A1(n_734),
.A2(n_709),
.B(n_718),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_730),
.B(n_711),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_731),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_734),
.A2(n_716),
.B1(n_701),
.B2(n_698),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_732),
.Y(n_747)
);

AOI32xp33_ASAP7_75t_L g748 ( 
.A1(n_737),
.A2(n_712),
.A3(n_711),
.B1(n_700),
.B2(n_715),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_SL g749 ( 
.A1(n_721),
.A2(n_729),
.B(n_722),
.C(n_725),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_724),
.B(n_695),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_738),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_736),
.Y(n_752)
);

OAI211xp5_ASAP7_75t_SL g753 ( 
.A1(n_743),
.A2(n_729),
.B(n_721),
.C(n_740),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_L g754 ( 
.A(n_746),
.B(n_708),
.C(n_723),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_749),
.B(n_739),
.C(n_719),
.Y(n_755)
);

AOI322xp5_ASAP7_75t_L g756 ( 
.A1(n_752),
.A2(n_735),
.A3(n_712),
.B1(n_700),
.B2(n_728),
.C1(n_699),
.C2(n_720),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_SL g757 ( 
.A1(n_748),
.A2(n_727),
.B(n_728),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_742),
.A2(n_720),
.B(n_717),
.Y(n_758)
);

OAI21xp33_ASAP7_75t_L g759 ( 
.A1(n_755),
.A2(n_752),
.B(n_750),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_754),
.A2(n_751),
.B1(n_747),
.B2(n_745),
.Y(n_760)
);

OAI22xp33_ASAP7_75t_SL g761 ( 
.A1(n_758),
.A2(n_717),
.B1(n_741),
.B2(n_615),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_753),
.Y(n_762)
);

AOI221xp5_ASAP7_75t_L g763 ( 
.A1(n_757),
.A2(n_744),
.B1(n_699),
.B2(n_697),
.C(n_713),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_756),
.A2(n_699),
.B1(n_705),
.B2(n_689),
.Y(n_764)
);

AND4x1_ASAP7_75t_L g765 ( 
.A(n_759),
.B(n_632),
.C(n_686),
.D(n_629),
.Y(n_765)
);

NAND3xp33_ASAP7_75t_L g766 ( 
.A(n_760),
.B(n_668),
.C(n_682),
.Y(n_766)
);

NOR2x1_ASAP7_75t_L g767 ( 
.A(n_762),
.B(n_620),
.Y(n_767)
);

NOR4xp25_ASAP7_75t_L g768 ( 
.A(n_764),
.B(n_713),
.C(n_628),
.D(n_629),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_763),
.B(n_689),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_767),
.Y(n_770)
);

NAND3xp33_ASAP7_75t_L g771 ( 
.A(n_768),
.B(n_668),
.C(n_680),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_770),
.B(n_766),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_771),
.A2(n_761),
.B1(n_769),
.B2(n_765),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_770),
.B(n_668),
.C(n_680),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_773),
.A2(n_680),
.B1(n_689),
.B2(n_705),
.Y(n_775)
);

NAND2x1_ASAP7_75t_L g776 ( 
.A(n_774),
.B(n_705),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_772),
.B(n_674),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_773),
.A2(n_637),
.B1(n_633),
.B2(n_624),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_772),
.B(n_620),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_778),
.B(n_637),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_779),
.A2(n_633),
.B(n_624),
.Y(n_781)
);

NAND3xp33_ASAP7_75t_L g782 ( 
.A(n_775),
.B(n_579),
.C(n_624),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_777),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_776),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_779),
.B(n_672),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_R g786 ( 
.A1(n_783),
.A2(n_674),
.B(n_672),
.C(n_595),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_785),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_784),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_780),
.A2(n_528),
.B(n_551),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_782),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_SL g791 ( 
.A(n_787),
.B(n_781),
.C(n_599),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_788),
.Y(n_792)
);

AOI21xp33_ASAP7_75t_L g793 ( 
.A1(n_788),
.A2(n_633),
.B(n_645),
.Y(n_793)
);

OAI21x1_ASAP7_75t_SL g794 ( 
.A1(n_790),
.A2(n_626),
.B(n_515),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_789),
.A2(n_786),
.B1(n_628),
.B2(n_642),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_792),
.A2(n_515),
.B(n_511),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_791),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_795),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_798),
.A2(n_793),
.B1(n_794),
.B2(n_642),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_797),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_800),
.A2(n_796),
.B(n_541),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_801),
.B(n_799),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_802),
.A2(n_510),
.B(n_541),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_803),
.A2(n_635),
.B1(n_645),
.B2(n_626),
.Y(n_804)
);


endmodule