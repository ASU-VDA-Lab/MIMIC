module fake_jpeg_12687_n_63 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_3),
.A2(n_1),
.B1(n_14),
.B2(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_32),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

OA21x2_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_26),
.B(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_0),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_22),
.B1(n_24),
.B2(n_27),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_40),
.B1(n_41),
.B2(n_30),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_27),
.B1(n_25),
.B2(n_23),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_8),
.B1(n_18),
.B2(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_48),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_29),
.B(n_1),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_19),
.C(n_13),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_49),
.C(n_42),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_50),
.B1(n_49),
.B2(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_2),
.B(n_3),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_2),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_53),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_9),
.C(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_5),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_11),
.Y(n_55)
);

OAI221xp5_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_51),
.B1(n_56),
.B2(n_7),
.C(n_5),
.Y(n_58)
);

NOR2xp67_ASAP7_75t_R g60 ( 
.A(n_57),
.B(n_58),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_60),
.B(n_59),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_55),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_6),
.Y(n_63)
);


endmodule