module fake_jpeg_6253_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_43),
.Y(n_69)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_19),
.B1(n_31),
.B2(n_33),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_29),
.B1(n_34),
.B2(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx2_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_30),
.C(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_65),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_51),
.B1(n_59),
.B2(n_61),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_19),
.B1(n_29),
.B2(n_33),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_25),
.B(n_28),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_30),
.C(n_28),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_55),
.B(n_60),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_17),
.B1(n_24),
.B2(n_35),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_58),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_29),
.B1(n_23),
.B2(n_18),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_23),
.B1(n_27),
.B2(n_17),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_35),
.Y(n_65)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_72),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_55),
.B1(n_49),
.B2(n_69),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_94),
.B1(n_53),
.B2(n_71),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_74),
.A2(n_80),
.B1(n_86),
.B2(n_58),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_47),
.B1(n_44),
.B2(n_42),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_75),
.A2(n_95),
.B1(n_102),
.B2(n_32),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_69),
.A2(n_17),
.B1(n_24),
.B2(n_25),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_81),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_24),
.B1(n_44),
.B2(n_47),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_98),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_53),
.Y(n_103)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_90),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_21),
.A3(n_25),
.B1(n_22),
.B2(n_20),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_76),
.C(n_73),
.Y(n_110)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_92),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

OA22x2_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_25),
.B1(n_30),
.B2(n_28),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_66),
.B(n_71),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_32),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_30),
.B1(n_28),
.B2(n_32),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_71),
.B1(n_68),
.B2(n_53),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_26),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_32),
.B1(n_26),
.B2(n_30),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_105),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_107),
.B1(n_108),
.B2(n_115),
.Y(n_138)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_114),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_112),
.A2(n_0),
.B(n_1),
.Y(n_155)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_52),
.B1(n_68),
.B2(n_72),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_72),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_126),
.B1(n_88),
.B2(n_78),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_52),
.B1(n_64),
.B2(n_58),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_123),
.B1(n_93),
.B2(n_81),
.Y(n_151)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_122),
.B(n_125),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_52),
.B1(n_64),
.B2(n_58),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_64),
.B1(n_58),
.B2(n_3),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_64),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_77),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_85),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_129),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_130),
.B(n_97),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_116),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_132),
.A2(n_155),
.B(n_161),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_147),
.B1(n_151),
.B2(n_153),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_89),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_156),
.C(n_12),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_137),
.B(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_146),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_97),
.B1(n_79),
.B2(n_78),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_101),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_111),
.B(n_90),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_101),
.B1(n_82),
.B2(n_95),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_77),
.B1(n_92),
.B2(n_96),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_127),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_158),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_81),
.B1(n_1),
.B2(n_3),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_0),
.C(n_1),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_160),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_119),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_108),
.B(n_3),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_4),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_118),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_181),
.C(n_143),
.Y(n_210)
);

XOR2x2_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_104),
.Y(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_132),
.B(n_141),
.C(n_154),
.D(n_161),
.Y(n_198)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_171),
.Y(n_214)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_169),
.B(n_159),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_114),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_117),
.B1(n_125),
.B2(n_116),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_173),
.A2(n_175),
.B1(n_141),
.B2(n_132),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_138),
.A2(n_112),
.B1(n_104),
.B2(n_115),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_104),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_178),
.Y(n_205)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_134),
.A2(n_123),
.B1(n_107),
.B2(n_120),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_151),
.Y(n_213)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_186),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_162),
.A2(n_120),
.B1(n_105),
.B2(n_121),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_155),
.B(n_133),
.Y(n_202)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_121),
.B1(n_120),
.B2(n_6),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_5),
.B(n_6),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_121),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_161),
.Y(n_220)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_157),
.B(n_105),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_145),
.B(n_11),
.Y(n_190)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_160),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_197),
.A2(n_198),
.B(n_202),
.Y(n_235)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_204),
.A2(n_207),
.B1(n_219),
.B2(n_222),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_147),
.B1(n_141),
.B2(n_134),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_218),
.C(n_223),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_167),
.A2(n_142),
.B(n_139),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_212),
.A2(n_225),
.B(n_178),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_220),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_217),
.Y(n_227)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_156),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_175),
.B1(n_194),
.B2(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_169),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_139),
.B1(n_6),
.B2(n_7),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_5),
.C(n_7),
.Y(n_223)
);

A2O1A1O1Ixp25_ASAP7_75t_L g224 ( 
.A1(n_164),
.A2(n_12),
.B(n_15),
.C(n_14),
.D(n_10),
.Y(n_224)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_7),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_228),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_185),
.B1(n_186),
.B2(n_163),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_229),
.A2(n_243),
.B1(n_245),
.B2(n_247),
.Y(n_254)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_232),
.Y(n_258)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_172),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_236),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_206),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_238),
.B(n_241),
.Y(n_265)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_196),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_168),
.Y(n_241)
);

OAI31xp33_ASAP7_75t_L g269 ( 
.A1(n_242),
.A2(n_215),
.A3(n_224),
.B(n_199),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_197),
.A2(n_185),
.B1(n_163),
.B2(n_192),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_197),
.A2(n_191),
.B1(n_183),
.B2(n_180),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_181),
.C(n_193),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_210),
.C(n_204),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_183),
.B1(n_179),
.B2(n_195),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_166),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_248),
.B(n_171),
.Y(n_268)
);

OAI22x1_ASAP7_75t_L g249 ( 
.A1(n_202),
.A2(n_183),
.B1(n_195),
.B2(n_193),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_249),
.A2(n_250),
.B1(n_211),
.B2(n_223),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_189),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_251),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_263),
.C(n_264),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_219),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_257),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_207),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_261),
.A2(n_230),
.B1(n_227),
.B2(n_232),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_198),
.C(n_220),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_214),
.C(n_211),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_222),
.C(n_195),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_271),
.C(n_226),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_267),
.Y(n_282)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_242),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_215),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_272),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_8),
.C(n_9),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_10),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_244),
.B1(n_238),
.B2(n_247),
.Y(n_273)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_273),
.Y(n_303)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_275),
.A2(n_288),
.B(n_289),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_267),
.A2(n_243),
.B1(n_245),
.B2(n_229),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_276),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_248),
.B1(n_236),
.B2(n_241),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_278),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_268),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_265),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_281),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_264),
.C(n_266),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_285),
.B(n_286),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_8),
.B(n_12),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_257),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_291),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_255),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_263),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_299),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_253),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_297),
.C(n_298),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_271),
.C(n_270),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_252),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_260),
.C(n_259),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_301),
.A2(n_289),
.B(n_287),
.Y(n_306)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_301),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_302),
.B(n_275),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_309),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_259),
.Y(n_308)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_281),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_295),
.B(n_273),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_294),
.A2(n_282),
.B(n_276),
.C(n_284),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_293),
.Y(n_315)
);

MAJx2_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_296),
.C(n_290),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_288),
.Y(n_316)
);

A2O1A1O1Ixp25_ASAP7_75t_L g329 ( 
.A1(n_316),
.A2(n_8),
.B(n_13),
.C(n_15),
.D(n_16),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_321),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_312),
.C(n_311),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_310),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_297),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_324),
.B(n_13),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_328),
.C(n_330),
.Y(n_333)
);

O2A1O1Ixp5_ASAP7_75t_L g327 ( 
.A1(n_316),
.A2(n_282),
.B(n_315),
.C(n_312),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_329),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_298),
.C(n_13),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_327),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_317),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_323),
.B1(n_322),
.B2(n_331),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_333),
.C(n_326),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);


endmodule