module fake_jpeg_51_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx16_ASAP7_75t_R g6 ( 
.A(n_1),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_SL g7 ( 
.A(n_5),
.B(n_1),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_4),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_15),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_10),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_18),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_10),
.A2(n_7),
.B1(n_11),
.B2(n_8),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_23),
.A2(n_18),
.B1(n_16),
.B2(n_14),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_15),
.B(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_22),
.B(n_13),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_23),
.B(n_21),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_17),
.B(n_8),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_17),
.C(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_6),
.C(n_20),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_31),
.B(n_24),
.Y(n_32)
);

AOI21x1_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_34),
.B(n_27),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_8),
.C(n_19),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.C(n_19),
.Y(n_37)
);


endmodule