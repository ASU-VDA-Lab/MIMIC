module fake_jpeg_3060_n_288 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_42),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_44),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_0),
.C(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_29),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_39),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_64),
.B(n_78),
.Y(n_129)
);

CKINVDCx6p67_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

INVxp67_ASAP7_75t_SL g127 ( 
.A(n_65),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_67),
.A2(n_95),
.B1(n_102),
.B2(n_88),
.Y(n_130)
);

BUFx2_ASAP7_75t_SL g68 ( 
.A(n_57),
.Y(n_68)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

HAxp5_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_28),
.CON(n_71),
.SN(n_71)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_76),
.Y(n_117)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_37),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_33),
.C(n_36),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_33),
.C(n_36),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_37),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_80),
.B(n_84),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_21),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_23),
.B1(n_18),
.B2(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_53),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_41),
.B(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_98),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_43),
.A2(n_24),
.B1(n_35),
.B2(n_50),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_21),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_40),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_101),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_40),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_41),
.A2(n_24),
.B1(n_35),
.B2(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_56),
.B(n_38),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_106),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_77),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_124),
.Y(n_152)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_125),
.Y(n_140)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_132),
.B1(n_72),
.B2(n_65),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_67),
.A2(n_38),
.B(n_32),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_107),
.B(n_88),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_86),
.A2(n_32),
.B1(n_30),
.B2(n_27),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_97),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_85),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_30),
.B1(n_27),
.B2(n_22),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_135),
.A2(n_22),
.B1(n_34),
.B2(n_74),
.Y(n_162)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_85),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_137),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_165),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_150),
.Y(n_180)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_148),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_149),
.A2(n_164),
.B(n_3),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_109),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_71),
.C(n_79),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_90),
.C(n_87),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_159),
.B1(n_3),
.B2(n_5),
.Y(n_196)
);

NOR2x1_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_65),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_13),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_103),
.B1(n_93),
.B2(n_75),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_66),
.Y(n_173)
);

OR2x4_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_66),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_103),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_108),
.B(n_24),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_166),
.B(n_167),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_35),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_34),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_168),
.B(n_1),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_110),
.B(n_93),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_114),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_122),
.B1(n_121),
.B2(n_120),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_173),
.A2(n_196),
.B1(n_162),
.B2(n_161),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_139),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_106),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_175),
.A2(n_183),
.B(n_184),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_112),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_115),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_135),
.B(n_116),
.C(n_126),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_179),
.B(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_126),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_188),
.C(n_193),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_90),
.B(n_128),
.C(n_81),
.D(n_4),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_81),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_87),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_192),
.C(n_194),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_1),
.C(n_2),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_142),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_7),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_160),
.C(n_163),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_197),
.B1(n_183),
.B2(n_173),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_219),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_147),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_210),
.C(n_175),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_209),
.B(n_213),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_157),
.C(n_163),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_186),
.B(n_160),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_212),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_156),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_156),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_174),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_215),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_142),
.B(n_139),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_153),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_216),
.B(n_189),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_200),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_177),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_231),
.C(n_235),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_219),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_229),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_225),
.Y(n_243)
);

AOI221xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_176),
.B1(n_188),
.B2(n_187),
.C(n_171),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_203),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_179),
.B1(n_170),
.B2(n_173),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_228),
.A2(n_201),
.B1(n_217),
.B2(n_218),
.Y(n_241)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_151),
.B(n_141),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_175),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_184),
.B(n_181),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_237),
.B(n_218),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_178),
.C(n_184),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_157),
.C(n_141),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_217),
.C(n_199),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_151),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_244),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_240),
.A2(n_223),
.B(n_236),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_241),
.A2(n_245),
.B1(n_248),
.B2(n_224),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_232),
.A2(n_224),
.B1(n_228),
.B2(n_237),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_200),
.C(n_209),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_247),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_198),
.B1(n_203),
.B2(n_207),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_224),
.A2(n_198),
.B(n_142),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_227),
.B(n_235),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_234),
.B1(n_227),
.B2(n_233),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_239),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_251),
.B(n_260),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_253),
.A2(n_240),
.B1(n_249),
.B2(n_241),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_261),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_257),
.A2(n_258),
.B(n_247),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_221),
.B(n_220),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_259),
.A2(n_246),
.B(n_238),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_193),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_148),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_267),
.B(n_260),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_248),
.B1(n_243),
.B2(n_245),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_264),
.A2(n_256),
.B1(n_252),
.B2(n_153),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_261),
.Y(n_267)
);

AOI31xp33_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_10),
.A3(n_11),
.B(n_12),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_272),
.B(n_275),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_271),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_269),
.A2(n_252),
.B(n_256),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_273),
.Y(n_277)
);

NAND4xp25_ASAP7_75t_SL g274 ( 
.A(n_268),
.B(n_7),
.C(n_9),
.D(n_10),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_10),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_266),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_279),
.A2(n_268),
.B(n_263),
.Y(n_282)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_280),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_282),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

AOI21x1_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_276),
.B(n_277),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_286),
.B(n_284),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_267),
.Y(n_288)
);


endmodule