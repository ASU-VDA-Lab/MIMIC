module fake_netlist_5_1202_n_1602 (n_137, n_91, n_82, n_122, n_10, n_140, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_1602);

input n_137;
input n_91;
input n_82;
input n_122;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1602;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_150;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_144;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1565;
wire n_182;
wire n_143;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_142;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_146;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_149;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_148;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_147;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_141;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_145;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_78),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_23),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_81),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_68),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_19),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_74),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_13),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_48),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_17),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_49),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_17),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_66),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_110),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_124),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_76),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_33),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_51),
.Y(n_163)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_32),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_31),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_24),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_96),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_12),
.Y(n_170)
);

BUFx2_ASAP7_75t_SL g171 ( 
.A(n_49),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_89),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_4),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_56),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_139),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_58),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_107),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_63),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_36),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_9),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_75),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_32),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_61),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_26),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_55),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_93),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_84),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_36),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_7),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_5),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_1),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_113),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_100),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_30),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_5),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_41),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_119),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_80),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_104),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_123),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_131),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_54),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_77),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_69),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_48),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_0),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_79),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_109),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_25),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_71),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_10),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_34),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_73),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_31),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_20),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_137),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_118),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_70),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_127),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_33),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_129),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_0),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_53),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_41),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_112),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_35),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_115),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_16),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_16),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_7),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_34),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_23),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_35),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_86),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_30),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_122),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_57),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_19),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_98),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_24),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_12),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_18),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_4),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_20),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_14),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_90),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_8),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_39),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_40),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_26),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_28),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_39),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_2),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_64),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_138),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_136),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_2),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_28),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_45),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_18),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_11),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_67),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_85),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_38),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_29),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_59),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_50),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_42),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_83),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_44),
.Y(n_275)
);

HB1xp67_ASAP7_75t_SL g276 ( 
.A(n_128),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_120),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_133),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_6),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_46),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_151),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_163),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_168),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_188),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_214),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_214),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_172),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_214),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_214),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_174),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_241),
.Y(n_292)
);

INVxp33_ASAP7_75t_SL g293 ( 
.A(n_254),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_164),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_142),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_267),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_175),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_142),
.Y(n_299)
);

INVxp33_ASAP7_75t_SL g300 ( 
.A(n_146),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_160),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_239),
.B(n_274),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_177),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_231),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_146),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_231),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_178),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_185),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_231),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_187),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_231),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_179),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_182),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_264),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_145),
.B(n_1),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_142),
.B(n_3),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_187),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_189),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_264),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_264),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_197),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_144),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_202),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_264),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_203),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_164),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_164),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_204),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_180),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_205),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_145),
.B(n_3),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_206),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_180),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_208),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_148),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_276),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_209),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_212),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_184),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_184),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_211),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_278),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_211),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_213),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_273),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_221),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_318),
.B(n_229),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_332),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_284),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_283),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_288),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_283),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_337),
.B(n_278),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_281),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_291),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_297),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_286),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_287),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_305),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_287),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_289),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_289),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_290),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_290),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_298),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_282),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_298),
.B(n_161),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_304),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_304),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_306),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_306),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_303),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_309),
.B(n_161),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_311),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_311),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_314),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_337),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_314),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_315),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_307),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_315),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_301),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_312),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_313),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_310),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_293),
.A2(n_196),
.B1(n_165),
.B2(n_181),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_321),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_325),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_325),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_319),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_334),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_323),
.B(n_242),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_334),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_295),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_295),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_299),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_341),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_299),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_322),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_323),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_323),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_343),
.B(n_278),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_343),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_349),
.B(n_329),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_390),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_349),
.B(n_331),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

BUFx10_ASAP7_75t_L g415 ( 
.A(n_350),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_407),
.B(n_228),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_348),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_407),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_407),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_398),
.B(n_300),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_338),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_361),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_407),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_398),
.A2(n_302),
.B(n_317),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_355),
.A2(n_347),
.B1(n_324),
.B2(n_339),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_336),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_361),
.B(n_345),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_353),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_403),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_408),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_310),
.Y(n_433)
);

OR2x6_ASAP7_75t_L g434 ( 
.A(n_369),
.B(n_171),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_207),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_359),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_380),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_380),
.B(n_294),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_359),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_362),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_408),
.Y(n_441)
);

INVx4_ASAP7_75t_SL g442 ( 
.A(n_408),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_408),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_352),
.B(n_228),
.Y(n_444)
);

BUFx10_ASAP7_75t_L g445 ( 
.A(n_357),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_358),
.B(n_244),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_362),
.B(n_310),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

AND2x2_ASAP7_75t_SL g449 ( 
.A(n_410),
.B(n_244),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_403),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_363),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_375),
.B(n_326),
.Y(n_452)
);

BUFx4f_ASAP7_75t_L g453 ( 
.A(n_403),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_365),
.Y(n_454)
);

NAND3xp33_ASAP7_75t_L g455 ( 
.A(n_391),
.B(n_328),
.C(n_327),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_354),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_383),
.B(n_333),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_365),
.B(n_242),
.Y(n_458)
);

OR2x6_ASAP7_75t_L g459 ( 
.A(n_369),
.B(n_186),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_356),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_387),
.B(n_335),
.Y(n_462)
);

OR2x6_ASAP7_75t_L g463 ( 
.A(n_376),
.B(n_186),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_403),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_403),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_388),
.B(n_207),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_371),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_371),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_403),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_373),
.Y(n_470)
);

INVxp33_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_363),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_373),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_354),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_400),
.B(n_207),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_374),
.B(n_224),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_354),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_363),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_396),
.B(n_308),
.Y(n_479)
);

INVx5_ASAP7_75t_L g480 ( 
.A(n_363),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_363),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_367),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_360),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_406),
.Y(n_484)
);

BUFx6f_ASAP7_75t_SL g485 ( 
.A(n_410),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_386),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_400),
.A2(n_273),
.B1(n_229),
.B2(n_240),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_381),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_376),
.B(n_207),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_397),
.B(n_330),
.Y(n_490)
);

AO21x2_ASAP7_75t_L g491 ( 
.A1(n_381),
.A2(n_156),
.B(n_149),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_367),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_400),
.A2(n_240),
.B1(n_191),
.B2(n_190),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_360),
.Y(n_494)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_367),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_386),
.A2(n_285),
.B1(n_296),
.B2(n_292),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_367),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_384),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_397),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_402),
.A2(n_200),
.B1(n_280),
.B2(n_263),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_402),
.A2(n_217),
.B1(n_236),
.B2(n_201),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_399),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_367),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_368),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_399),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_402),
.A2(n_253),
.B1(n_250),
.B2(n_216),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_405),
.B(n_207),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_401),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_405),
.A2(n_248),
.B1(n_261),
.B2(n_230),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_360),
.Y(n_510)
);

BUFx8_ASAP7_75t_SL g511 ( 
.A(n_405),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_367),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_401),
.B(n_255),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_378),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_378),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_404),
.B(n_234),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_378),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_385),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_385),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_378),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_392),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_366),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_366),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_378),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_392),
.B(n_393),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_393),
.A2(n_215),
.B1(n_261),
.B2(n_230),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_SL g527 ( 
.A(n_351),
.B(n_243),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_378),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_379),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_351),
.B(n_330),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_366),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_372),
.B(n_158),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_351),
.B(n_226),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_351),
.B(n_269),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_364),
.B(n_227),
.C(n_195),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_364),
.B(n_395),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_364),
.B(n_141),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_L g538 ( 
.A(n_379),
.B(n_215),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_372),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_379),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_372),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_379),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_379),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_379),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_395),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_377),
.B(n_340),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_395),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_394),
.A2(n_147),
.B1(n_159),
.B2(n_277),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_394),
.A2(n_147),
.B1(n_159),
.B2(n_277),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_394),
.B(n_141),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_411),
.B(n_394),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_508),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_413),
.B(n_143),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_420),
.B(n_394),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_530),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_420),
.B(n_394),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_530),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_412),
.B(n_143),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_425),
.B(n_537),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_530),
.Y(n_560)
);

AND2x6_ASAP7_75t_SL g561 ( 
.A(n_427),
.B(n_340),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_460),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_519),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_537),
.B(n_395),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_526),
.A2(n_249),
.B1(n_262),
.B2(n_230),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_525),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_414),
.B(n_155),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_516),
.A2(n_232),
.B1(n_272),
.B2(n_271),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_437),
.B(n_167),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_438),
.B(n_155),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_534),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_449),
.B(n_157),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_513),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_505),
.B(n_157),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_449),
.B(n_268),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_421),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_527),
.A2(n_268),
.B1(n_272),
.B2(n_271),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_527),
.A2(n_218),
.B1(n_176),
.B2(n_260),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_496),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_430),
.Y(n_580)
);

INVx8_ASAP7_75t_L g581 ( 
.A(n_485),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_434),
.A2(n_169),
.B1(n_192),
.B2(n_193),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_436),
.B(n_395),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_439),
.B(n_440),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_454),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_461),
.B(n_183),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_423),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_456),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_467),
.B(n_194),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_456),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_468),
.B(n_198),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_470),
.B(n_473),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_488),
.B(n_222),
.Y(n_593)
);

OR2x6_ASAP7_75t_L g594 ( 
.A(n_434),
.B(n_223),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_474),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_486),
.B(n_434),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_434),
.B(n_150),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_498),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_474),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_518),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_521),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_531),
.B(n_251),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_428),
.B(n_259),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_499),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_502),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_539),
.B(n_377),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_444),
.A2(n_261),
.B1(n_230),
.B2(n_215),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_477),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_541),
.B(n_377),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_444),
.B(n_166),
.Y(n_610)
);

O2A1O1Ixp5_ASAP7_75t_L g611 ( 
.A1(n_416),
.A2(n_389),
.B(n_382),
.C(n_346),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_415),
.B(n_256),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_446),
.B(n_170),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_550),
.B(n_422),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_466),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_446),
.B(n_173),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_504),
.B(n_150),
.Y(n_617)
);

NAND3xp33_ASAP7_75t_L g618 ( 
.A(n_535),
.B(n_245),
.C(n_199),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_L g619 ( 
.A(n_426),
.B(n_52),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_543),
.B(n_389),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_433),
.B(n_389),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_490),
.Y(n_622)
);

CKINVDCx11_ASAP7_75t_R g623 ( 
.A(n_415),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_476),
.B(n_215),
.Y(n_624)
);

NOR2xp67_ASAP7_75t_SL g625 ( 
.A(n_526),
.B(n_215),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_466),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_455),
.B(n_152),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_548),
.B(n_230),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_477),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_452),
.B(n_246),
.C(n_210),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_429),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_471),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_447),
.Y(n_633)
);

OAI21xp33_ASAP7_75t_L g634 ( 
.A1(n_471),
.A2(n_153),
.B(n_154),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_533),
.A2(n_261),
.B1(n_220),
.B2(n_225),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_429),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_459),
.B(n_162),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_549),
.B(n_238),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_459),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_415),
.B(n_256),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_432),
.B(n_257),
.Y(n_641)
);

BUFx5_ASAP7_75t_L g642 ( 
.A(n_418),
.Y(n_642)
);

AND2x2_ASAP7_75t_SL g643 ( 
.A(n_509),
.B(n_346),
.Y(n_643)
);

AOI221xp5_ASAP7_75t_L g644 ( 
.A1(n_500),
.A2(n_162),
.B1(n_219),
.B2(n_279),
.C(n_275),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_511),
.B(n_459),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_441),
.B(n_258),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_431),
.B(n_252),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_483),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_445),
.B(n_233),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_511),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_431),
.B(n_235),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_R g652 ( 
.A(n_445),
.B(n_237),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_459),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_431),
.B(n_247),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_L g655 ( 
.A1(n_463),
.A2(n_270),
.B1(n_265),
.B2(n_279),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_484),
.B(n_452),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_450),
.B(n_344),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_450),
.B(n_344),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_450),
.B(n_342),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_464),
.B(n_342),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_464),
.B(n_465),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_484),
.B(n_256),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_464),
.B(n_465),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_484),
.B(n_275),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_483),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_463),
.B(n_266),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_463),
.B(n_266),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_457),
.B(n_265),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_491),
.A2(n_219),
.B1(n_8),
.B2(n_9),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_SL g670 ( 
.A(n_485),
.B(n_6),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_463),
.B(n_10),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_491),
.A2(n_82),
.B1(n_134),
.B2(n_130),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_462),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_429),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_465),
.B(n_65),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_469),
.B(n_72),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_453),
.A2(n_60),
.B(n_125),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_546),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_494),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_532),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_462),
.B(n_11),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_479),
.B(n_13),
.Y(n_682)
);

BUFx5_ASAP7_75t_L g683 ( 
.A(n_418),
.Y(n_683)
);

O2A1O1Ixp5_ASAP7_75t_L g684 ( 
.A1(n_416),
.A2(n_14),
.B(n_15),
.C(n_21),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_479),
.B(n_15),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_478),
.B(n_497),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_509),
.A2(n_21),
.B1(n_22),
.B2(n_27),
.Y(n_687)
);

NOR3xp33_ASAP7_75t_L g688 ( 
.A(n_458),
.B(n_22),
.C(n_27),
.Y(n_688)
);

NOR2xp67_ASAP7_75t_L g689 ( 
.A(n_489),
.B(n_92),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_487),
.B(n_37),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_532),
.B(n_37),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_532),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_472),
.Y(n_693)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_451),
.Y(n_694)
);

NAND2x1p5_ASAP7_75t_L g695 ( 
.A(n_419),
.B(n_88),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_472),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_493),
.B(n_487),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_493),
.B(n_40),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_544),
.B(n_42),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_478),
.B(n_514),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_497),
.B(n_517),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_510),
.Y(n_702)
);

OAI321xp33_ASAP7_75t_L g703 ( 
.A1(n_669),
.A2(n_500),
.A3(n_501),
.B1(n_506),
.B2(n_489),
.C(n_507),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_560),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_573),
.B(n_506),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_555),
.Y(n_706)
);

O2A1O1Ixp5_ASAP7_75t_L g707 ( 
.A1(n_559),
.A2(n_507),
.B(n_453),
.C(n_536),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_R g708 ( 
.A(n_579),
.B(n_529),
.Y(n_708)
);

O2A1O1Ixp5_ASAP7_75t_L g709 ( 
.A1(n_554),
.A2(n_443),
.B(n_424),
.C(n_419),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_614),
.A2(n_419),
.B(n_424),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_551),
.A2(n_424),
.B(n_443),
.Y(n_711)
);

AND2x2_ASAP7_75t_SL g712 ( 
.A(n_565),
.B(n_501),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_560),
.Y(n_713)
);

AOI21xp33_ASAP7_75t_L g714 ( 
.A1(n_553),
.A2(n_435),
.B(n_547),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_553),
.B(n_443),
.Y(n_715)
);

AO21x1_ASAP7_75t_L g716 ( 
.A1(n_628),
.A2(n_435),
.B(n_538),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_564),
.A2(n_448),
.B(n_542),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_560),
.B(n_615),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_626),
.A2(n_545),
.B1(n_515),
.B2(n_482),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_633),
.A2(n_492),
.B1(n_515),
.B2(n_482),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_571),
.B(n_451),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_610),
.A2(n_514),
.B(n_540),
.C(n_517),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_694),
.A2(n_542),
.B(n_448),
.Y(n_723)
);

AOI21x1_ASAP7_75t_L g724 ( 
.A1(n_556),
.A2(n_522),
.B(n_523),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_557),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_678),
.B(n_574),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_697),
.A2(n_523),
.B1(n_522),
.B2(n_492),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_565),
.A2(n_540),
.B1(n_529),
.B2(n_497),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_588),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_693),
.Y(n_730)
);

INVx3_ASAP7_75t_SL g731 ( 
.A(n_581),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_694),
.A2(n_542),
.B(n_448),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_613),
.A2(n_529),
.B(n_514),
.C(n_512),
.Y(n_733)
);

BUFx12f_ASAP7_75t_L g734 ( 
.A(n_623),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_621),
.A2(n_524),
.B(n_528),
.Y(n_735)
);

AOI21x1_ASAP7_75t_L g736 ( 
.A1(n_624),
.A2(n_442),
.B(n_524),
.Y(n_736)
);

NAND3xp33_ASAP7_75t_L g737 ( 
.A(n_570),
.B(n_528),
.C(n_481),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_693),
.A2(n_528),
.B(n_481),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_566),
.B(n_528),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_696),
.A2(n_663),
.B(n_661),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_576),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_587),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_696),
.A2(n_451),
.B(n_481),
.Y(n_743)
);

CKINVDCx8_ASAP7_75t_R g744 ( 
.A(n_581),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_686),
.A2(n_701),
.B(n_700),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_673),
.B(n_481),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_580),
.B(n_451),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_562),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_585),
.B(n_442),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_598),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_616),
.A2(n_520),
.B(n_503),
.C(n_495),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_590),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_687),
.A2(n_520),
.B1(n_503),
.B2(n_495),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_595),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_668),
.B(n_43),
.C(n_44),
.Y(n_755)
);

CKINVDCx10_ASAP7_75t_R g756 ( 
.A(n_569),
.Y(n_756)
);

O2A1O1Ixp5_ASAP7_75t_L g757 ( 
.A1(n_584),
.A2(n_475),
.B(n_503),
.C(n_495),
.Y(n_757)
);

INVx3_ASAP7_75t_SL g758 ( 
.A(n_581),
.Y(n_758)
);

AND2x6_ASAP7_75t_L g759 ( 
.A(n_690),
.B(n_672),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_643),
.B(n_520),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_SL g761 ( 
.A(n_685),
.B(n_475),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_599),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_L g763 ( 
.A1(n_611),
.A2(n_475),
.B(n_495),
.Y(n_763)
);

BUFx2_ASAP7_75t_SL g764 ( 
.A(n_650),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_578),
.A2(n_503),
.B(n_480),
.C(n_46),
.Y(n_765)
);

AOI21x1_ASAP7_75t_L g766 ( 
.A1(n_583),
.A2(n_480),
.B(n_475),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_569),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_643),
.B(n_480),
.Y(n_768)
);

A2O1A1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_558),
.A2(n_43),
.B(n_45),
.C(n_47),
.Y(n_769)
);

O2A1O1Ixp5_ASAP7_75t_L g770 ( 
.A1(n_592),
.A2(n_103),
.B(n_87),
.C(n_94),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_636),
.A2(n_97),
.B(n_101),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_631),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_656),
.B(n_106),
.Y(n_773)
);

BUFx4f_ASAP7_75t_L g774 ( 
.A(n_596),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_600),
.B(n_47),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_558),
.A2(n_111),
.B(n_114),
.C(n_121),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_601),
.B(n_622),
.Y(n_777)
);

BUFx10_ASAP7_75t_L g778 ( 
.A(n_645),
.Y(n_778)
);

OR2x6_ASAP7_75t_SL g779 ( 
.A(n_698),
.B(n_627),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_604),
.B(n_605),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_657),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_563),
.B(n_612),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_569),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_702),
.B(n_608),
.Y(n_784)
);

OAI21xp33_ASAP7_75t_L g785 ( 
.A1(n_634),
.A2(n_567),
.B(n_644),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_640),
.B(n_567),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_682),
.B(n_619),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_681),
.A2(n_638),
.B(n_669),
.C(n_572),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_674),
.A2(n_620),
.B(n_641),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_629),
.B(n_648),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_664),
.B(n_568),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_674),
.A2(n_646),
.B(n_631),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_552),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_665),
.B(n_679),
.Y(n_794)
);

O2A1O1Ixp5_ASAP7_75t_L g795 ( 
.A1(n_647),
.A2(n_651),
.B(n_654),
.C(n_603),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_631),
.A2(n_606),
.B(n_609),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_658),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_630),
.A2(n_639),
.B1(n_653),
.B2(n_575),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_617),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_SL g800 ( 
.A(n_625),
.B(n_671),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_695),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_659),
.Y(n_802)
);

OA22x2_ASAP7_75t_L g803 ( 
.A1(n_632),
.A2(n_594),
.B1(n_577),
.B2(n_692),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_692),
.B(n_680),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_684),
.A2(n_676),
.B(n_675),
.Y(n_805)
);

BUFx12f_ASAP7_75t_L g806 ( 
.A(n_561),
.Y(n_806)
);

NAND2x1p5_ASAP7_75t_L g807 ( 
.A(n_689),
.B(n_677),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_586),
.B(n_591),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_594),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_589),
.B(n_593),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_642),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_660),
.A2(n_602),
.B(n_683),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_594),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_642),
.A2(n_683),
.B(n_618),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_667),
.A2(n_635),
.B(n_691),
.C(n_644),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_699),
.A2(n_667),
.B(n_607),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_687),
.A2(n_597),
.B1(n_666),
.B2(n_637),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_683),
.B(n_655),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_652),
.B(n_649),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_662),
.B(n_655),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_670),
.A2(n_645),
.B(n_688),
.Y(n_821)
);

AND2x2_ASAP7_75t_SL g822 ( 
.A(n_688),
.B(n_565),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_560),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_614),
.A2(n_551),
.B(n_564),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_614),
.A2(n_551),
.B(n_564),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_565),
.A2(n_687),
.B1(n_559),
.B2(n_669),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_559),
.B(n_411),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_555),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_560),
.B(n_417),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_555),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_553),
.B(n_411),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_614),
.A2(n_551),
.B(n_564),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_555),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_559),
.B(n_614),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_614),
.A2(n_551),
.B(n_564),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_614),
.A2(n_551),
.B(n_564),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_614),
.A2(n_551),
.B(n_564),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_614),
.A2(n_551),
.B(n_564),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_560),
.B(n_417),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_614),
.A2(n_551),
.B(n_564),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_614),
.A2(n_551),
.B(n_564),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_559),
.B(n_411),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_555),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_555),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_566),
.B(n_639),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_559),
.A2(n_614),
.B(n_697),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_614),
.A2(n_551),
.B(n_564),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_560),
.B(n_417),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_555),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_559),
.A2(n_553),
.B(n_613),
.C(n_610),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_560),
.B(n_417),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_694),
.Y(n_852)
);

O2A1O1Ixp5_ASAP7_75t_L g853 ( 
.A1(n_559),
.A2(n_349),
.B(n_556),
.C(n_554),
.Y(n_853)
);

A2O1A1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_559),
.A2(n_553),
.B(n_613),
.C(n_610),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_559),
.B(n_614),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_555),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_559),
.B(n_614),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_559),
.B(n_411),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_SL g859 ( 
.A1(n_685),
.A2(n_516),
.B1(n_656),
.B2(n_449),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_614),
.A2(n_551),
.B(n_564),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_559),
.B(n_411),
.Y(n_861)
);

AO32x2_ASAP7_75t_L g862 ( 
.A1(n_615),
.A2(n_626),
.A3(n_582),
.B1(n_653),
.B2(n_639),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_562),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_555),
.Y(n_864)
);

OAI21xp33_ASAP7_75t_L g865 ( 
.A1(n_570),
.A2(n_302),
.B(n_349),
.Y(n_865)
);

INVx5_ASAP7_75t_L g866 ( 
.A(n_631),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_623),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_741),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_850),
.B(n_854),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_824),
.A2(n_832),
.B(n_825),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_853),
.A2(n_842),
.B(n_827),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_834),
.B(n_855),
.Y(n_872)
);

BUFx12f_ASAP7_75t_L g873 ( 
.A(n_748),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_858),
.A2(n_861),
.B(n_855),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_750),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_831),
.B(n_834),
.Y(n_876)
);

OAI21x1_ASAP7_75t_L g877 ( 
.A1(n_745),
.A2(n_740),
.B(n_724),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_865),
.B(n_726),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_857),
.A2(n_846),
.B(n_707),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_742),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_704),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_782),
.B(n_786),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_835),
.A2(n_837),
.B(n_836),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_784),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_736),
.A2(n_711),
.B(n_717),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_857),
.B(n_715),
.Y(n_886)
);

CKINVDCx6p67_ASAP7_75t_R g887 ( 
.A(n_731),
.Y(n_887)
);

OAI21x1_ASAP7_75t_L g888 ( 
.A1(n_814),
.A2(n_735),
.B(n_792),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_723),
.A2(n_732),
.B(n_812),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_852),
.B(n_826),
.Y(n_890)
);

NAND2x1p5_ASAP7_75t_L g891 ( 
.A(n_713),
.B(n_866),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_826),
.B(n_785),
.Y(n_892)
);

AO31x2_ASAP7_75t_L g893 ( 
.A1(n_722),
.A2(n_733),
.A3(n_716),
.B(n_860),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_712),
.A2(n_788),
.B(n_703),
.C(n_815),
.Y(n_894)
);

AND2x6_ASAP7_75t_L g895 ( 
.A(n_801),
.B(n_811),
.Y(n_895)
);

O2A1O1Ixp5_ASAP7_75t_L g896 ( 
.A1(n_805),
.A2(n_816),
.B(n_847),
.C(n_840),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_808),
.B(n_810),
.Y(n_897)
);

AOI21x1_ASAP7_75t_L g898 ( 
.A1(n_838),
.A2(n_841),
.B(n_789),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_784),
.Y(n_899)
);

NOR2xp67_ASAP7_75t_SL g900 ( 
.A(n_744),
.B(n_703),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_828),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_709),
.A2(n_811),
.B(n_796),
.Y(n_902)
);

NOR2xp67_ASAP7_75t_L g903 ( 
.A(n_799),
.B(n_819),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_822),
.B(n_777),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_863),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_781),
.B(n_797),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_705),
.B(n_774),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_802),
.B(n_746),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_833),
.Y(n_909)
);

OAI21x1_ASAP7_75t_L g910 ( 
.A1(n_710),
.A2(n_738),
.B(n_743),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_845),
.B(n_804),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_845),
.B(n_804),
.Y(n_912)
);

OAI21x1_ASAP7_75t_SL g913 ( 
.A1(n_760),
.A2(n_768),
.B(n_771),
.Y(n_913)
);

NAND2x1p5_ASAP7_75t_L g914 ( 
.A(n_713),
.B(n_866),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_843),
.B(n_849),
.Y(n_915)
);

OAI21x1_ASAP7_75t_L g916 ( 
.A1(n_766),
.A2(n_757),
.B(n_763),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_856),
.Y(n_917)
);

BUFx10_ASAP7_75t_L g918 ( 
.A(n_820),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_706),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_759),
.B(n_725),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_758),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_704),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_759),
.B(n_830),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_759),
.B(n_844),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_SL g925 ( 
.A1(n_859),
.A2(n_817),
.B(n_821),
.Y(n_925)
);

OAI21x1_ASAP7_75t_L g926 ( 
.A1(n_763),
.A2(n_727),
.B(n_795),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_807),
.A2(n_787),
.B(n_714),
.Y(n_927)
);

NAND2x1p5_ASAP7_75t_L g928 ( 
.A(n_866),
.B(n_704),
.Y(n_928)
);

OAI22x1_ASAP7_75t_L g929 ( 
.A1(n_798),
.A2(n_791),
.B1(n_767),
.B2(n_783),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_818),
.A2(n_816),
.B1(n_760),
.B2(n_768),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_793),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_790),
.A2(n_794),
.B(n_747),
.Y(n_932)
);

NOR2xp67_ASAP7_75t_L g933 ( 
.A(n_780),
.B(n_734),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_759),
.B(n_864),
.Y(n_934)
);

AO31x2_ASAP7_75t_L g935 ( 
.A1(n_751),
.A2(n_728),
.A3(n_769),
.B(n_765),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_729),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_708),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_714),
.A2(n_800),
.B(n_753),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_823),
.B(n_739),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_866),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_752),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_774),
.B(n_779),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_823),
.B(n_775),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_800),
.A2(n_753),
.B(n_801),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_749),
.A2(n_737),
.B(n_728),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_755),
.A2(n_761),
.B(n_776),
.C(n_770),
.Y(n_946)
);

O2A1O1Ixp5_ASAP7_75t_L g947 ( 
.A1(n_773),
.A2(n_718),
.B(n_730),
.C(n_721),
.Y(n_947)
);

AO31x2_ASAP7_75t_L g948 ( 
.A1(n_862),
.A2(n_762),
.A3(n_754),
.B(n_809),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_761),
.B(n_730),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_829),
.B(n_839),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_848),
.B(n_851),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_720),
.B(n_772),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_764),
.B(n_813),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_772),
.B(n_719),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_813),
.B(n_803),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_813),
.B(n_778),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_778),
.B(n_862),
.Y(n_957)
);

OAI21x1_ASAP7_75t_SL g958 ( 
.A1(n_862),
.A2(n_756),
.B(n_806),
.Y(n_958)
);

NAND2x1p5_ASAP7_75t_L g959 ( 
.A(n_867),
.B(n_713),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_850),
.A2(n_854),
.B(n_853),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_831),
.B(n_827),
.Y(n_961)
);

NOR2xp67_ASAP7_75t_L g962 ( 
.A(n_799),
.B(n_573),
.Y(n_962)
);

AOI21x1_ASAP7_75t_SL g963 ( 
.A1(n_827),
.A2(n_559),
.B(n_842),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_L g964 ( 
.A(n_831),
.B(n_685),
.C(n_859),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_799),
.B(n_573),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_824),
.A2(n_832),
.B(n_825),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_831),
.B(n_827),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_742),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_730),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_831),
.B(n_827),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_866),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_831),
.B(n_827),
.Y(n_972)
);

AO221x1_ASAP7_75t_L g973 ( 
.A1(n_826),
.A2(n_655),
.B1(n_632),
.B2(n_817),
.C(n_801),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_831),
.B(n_827),
.Y(n_974)
);

AOI21x1_ASAP7_75t_L g975 ( 
.A1(n_736),
.A2(n_724),
.B(n_564),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_704),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_745),
.A2(n_740),
.B(n_724),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_845),
.B(n_804),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_745),
.A2(n_740),
.B(n_724),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_831),
.B(n_861),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_850),
.A2(n_854),
.B(n_853),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_706),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_745),
.A2(n_740),
.B(n_724),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_850),
.B(n_854),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_745),
.A2(n_740),
.B(n_724),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_706),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_831),
.B(n_827),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_745),
.A2(n_740),
.B(n_724),
.Y(n_988)
);

OA22x2_ASAP7_75t_L g989 ( 
.A1(n_785),
.A2(n_391),
.B1(n_826),
.B2(n_865),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_831),
.B(n_827),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_748),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_826),
.A2(n_831),
.B(n_785),
.C(n_850),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_870),
.A2(n_966),
.B(n_883),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_882),
.B(n_907),
.Y(n_994)
);

NAND3xp33_ASAP7_75t_L g995 ( 
.A(n_964),
.B(n_980),
.C(n_992),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_980),
.A2(n_925),
.B1(n_904),
.B2(n_987),
.Y(n_996)
);

INVx5_ASAP7_75t_L g997 ( 
.A(n_971),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_870),
.A2(n_966),
.B(n_883),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_961),
.A2(n_972),
.B1(n_990),
.B2(n_974),
.Y(n_999)
);

OAI21xp33_ASAP7_75t_L g1000 ( 
.A1(n_967),
.A2(n_970),
.B(n_897),
.Y(n_1000)
);

OR2x6_ASAP7_75t_L g1001 ( 
.A(n_873),
.B(n_921),
.Y(n_1001)
);

INVx6_ASAP7_75t_SL g1002 ( 
.A(n_911),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_887),
.Y(n_1003)
);

BUFx10_ASAP7_75t_L g1004 ( 
.A(n_911),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_991),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_905),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_971),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_953),
.Y(n_1008)
);

OA21x2_ASAP7_75t_L g1009 ( 
.A1(n_938),
.A2(n_879),
.B(n_960),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_884),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_876),
.B(n_905),
.Y(n_1011)
);

OR2x6_ASAP7_75t_L g1012 ( 
.A(n_921),
.B(n_931),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_971),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_874),
.B(n_886),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_878),
.B(n_872),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_878),
.B(n_872),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_906),
.B(n_899),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_912),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_903),
.A2(n_989),
.B1(n_962),
.B2(n_965),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_912),
.B(n_978),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_908),
.B(n_992),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_978),
.B(n_942),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_928),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_968),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_989),
.B(n_871),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_868),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_956),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_973),
.A2(n_918),
.B1(n_900),
.B2(n_892),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_937),
.B(n_880),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_955),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_976),
.B(n_881),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_895),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_875),
.B(n_901),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_918),
.B(n_894),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_915),
.B(n_909),
.Y(n_1035)
);

OAI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_920),
.A2(n_934),
.B1(n_924),
.B2(n_923),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_917),
.B(n_890),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_869),
.A2(n_984),
.B1(n_929),
.B2(n_957),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_880),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_R g1040 ( 
.A(n_881),
.B(n_922),
.Y(n_1040)
);

OA21x2_ASAP7_75t_L g1041 ( 
.A1(n_938),
.A2(n_981),
.B(n_926),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_950),
.B(n_919),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_982),
.B(n_986),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_950),
.B(n_951),
.Y(n_1044)
);

OAI221xp5_ASAP7_75t_L g1045 ( 
.A1(n_933),
.A2(n_869),
.B1(n_984),
.B2(n_946),
.C(n_943),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_936),
.B(n_941),
.Y(n_1046)
);

INVxp67_ASAP7_75t_SL g1047 ( 
.A(n_928),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_959),
.B(n_914),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_976),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_944),
.A2(n_946),
.B(n_927),
.C(n_896),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_895),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_927),
.B(n_959),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_930),
.B(n_969),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_922),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_891),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_939),
.B(n_969),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_891),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_948),
.B(n_952),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_949),
.B(n_954),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_914),
.Y(n_1060)
);

INVx5_ASAP7_75t_SL g1061 ( 
.A(n_958),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_949),
.B(n_932),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_895),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_948),
.B(n_935),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_940),
.B(n_895),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_948),
.B(n_935),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_940),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_L g1068 ( 
.A(n_895),
.B(n_963),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_948),
.Y(n_1069)
);

AND2x2_ASAP7_75t_SL g1070 ( 
.A(n_947),
.B(n_963),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_935),
.B(n_888),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_935),
.B(n_893),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_945),
.B(n_910),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_893),
.B(n_902),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_893),
.Y(n_1075)
);

AND2x6_ASAP7_75t_L g1076 ( 
.A(n_947),
.B(n_896),
.Y(n_1076)
);

NOR2x1_ASAP7_75t_SL g1077 ( 
.A(n_898),
.B(n_975),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_893),
.B(n_889),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_877),
.B(n_979),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_977),
.A2(n_983),
.B(n_985),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_916),
.B(n_988),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_885),
.B(n_882),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_868),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_980),
.A2(n_961),
.B1(n_970),
.B2(n_967),
.Y(n_1084)
);

BUFx10_ASAP7_75t_L g1085 ( 
.A(n_911),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_905),
.Y(n_1086)
);

INVx4_ASAP7_75t_L g1087 ( 
.A(n_971),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_980),
.A2(n_961),
.B1(n_970),
.B2(n_967),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_873),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_882),
.B(n_907),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_911),
.B(n_912),
.Y(n_1091)
);

OAI21xp33_ASAP7_75t_L g1092 ( 
.A1(n_980),
.A2(n_865),
.B(n_831),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_905),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_884),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_882),
.B(n_907),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_980),
.B(n_961),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_980),
.A2(n_854),
.B(n_850),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_887),
.Y(n_1098)
);

AND2x6_ASAP7_75t_L g1099 ( 
.A(n_971),
.B(n_801),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_980),
.B(n_831),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_897),
.B(n_859),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_980),
.A2(n_961),
.B1(n_970),
.B2(n_967),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_911),
.B(n_912),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_971),
.Y(n_1104)
);

NOR2xp67_ASAP7_75t_L g1105 ( 
.A(n_931),
.B(n_573),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_873),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_991),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_980),
.A2(n_831),
.B(n_854),
.C(n_850),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_980),
.B(n_961),
.Y(n_1109)
);

INVx5_ASAP7_75t_L g1110 ( 
.A(n_971),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_980),
.A2(n_831),
.B(n_854),
.C(n_850),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_868),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_868),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_884),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_980),
.A2(n_961),
.B1(n_970),
.B2(n_967),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_980),
.A2(n_831),
.B(n_854),
.C(n_850),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_884),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_868),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_884),
.Y(n_1119)
);

AO21x2_ASAP7_75t_L g1120 ( 
.A1(n_1080),
.A2(n_998),
.B(n_993),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1100),
.A2(n_1092),
.B1(n_995),
.B2(n_1101),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1026),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_996),
.B(n_1034),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_1065),
.B(n_1048),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1028),
.B(n_1097),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1000),
.A2(n_1045),
.B1(n_1115),
.B2(n_1102),
.Y(n_1126)
);

BUFx2_ASAP7_75t_SL g1127 ( 
.A(n_997),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1026),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_SL g1129 ( 
.A1(n_1084),
.A2(n_1088),
.B1(n_1061),
.B2(n_999),
.Y(n_1129)
);

BUFx2_ASAP7_75t_R g1130 ( 
.A(n_1003),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_1005),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1065),
.B(n_1048),
.Y(n_1132)
);

BUFx2_ASAP7_75t_SL g1133 ( 
.A(n_1098),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1083),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_1058),
.B(n_1025),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1118),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_1086),
.Y(n_1137)
);

NAND2x1p5_ASAP7_75t_L g1138 ( 
.A(n_1052),
.B(n_1071),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1112),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1113),
.Y(n_1140)
);

BUFx12f_ASAP7_75t_L g1141 ( 
.A(n_1106),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1046),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1010),
.Y(n_1143)
);

AOI22x1_ASAP7_75t_L g1144 ( 
.A1(n_1119),
.A2(n_1117),
.B1(n_1114),
.B2(n_1094),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1094),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_1093),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1039),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1082),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1096),
.B(n_1109),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_1071),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_1072),
.B(n_1064),
.Y(n_1151)
);

AOI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1079),
.A2(n_1053),
.B(n_1073),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1063),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1108),
.A2(n_1111),
.B(n_1116),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1119),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1033),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1063),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1017),
.A2(n_1019),
.B1(n_1014),
.B2(n_1038),
.Y(n_1158)
);

OAI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1030),
.A2(n_1015),
.B1(n_1016),
.B2(n_1011),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_1006),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1107),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_994),
.B(n_1090),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_SL g1163 ( 
.A1(n_1061),
.A2(n_1095),
.B1(n_1021),
.B2(n_1059),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1033),
.Y(n_1164)
);

BUFx2_ASAP7_75t_R g1165 ( 
.A(n_1089),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1001),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1035),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_1018),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1029),
.B(n_1044),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1043),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1042),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1037),
.B(n_1008),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1056),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1024),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1027),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1069),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1075),
.B(n_1009),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1032),
.B(n_1051),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1067),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1105),
.Y(n_1180)
);

AOI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1073),
.A2(n_1062),
.B(n_1078),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1054),
.Y(n_1182)
);

AO21x2_ASAP7_75t_L g1183 ( 
.A1(n_1077),
.A2(n_1050),
.B(n_1081),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1041),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1009),
.B(n_1066),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1104),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1104),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1007),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_SL g1189 ( 
.A1(n_1022),
.A2(n_1103),
.B1(n_1091),
.B2(n_1020),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1012),
.A2(n_1036),
.B1(n_1047),
.B2(n_1002),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1074),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1070),
.B(n_1078),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1007),
.Y(n_1193)
);

AO21x2_ASAP7_75t_L g1194 ( 
.A1(n_1068),
.A2(n_1076),
.B(n_1040),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1032),
.Y(n_1195)
);

INVx6_ASAP7_75t_L g1196 ( 
.A(n_1110),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1020),
.B(n_1091),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1076),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1007),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1103),
.A2(n_1076),
.B1(n_1002),
.B2(n_1001),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1060),
.B(n_1031),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1076),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1110),
.A2(n_1055),
.B1(n_1057),
.B2(n_1023),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1055),
.A2(n_1057),
.B1(n_1023),
.B2(n_1087),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1004),
.A2(n_1085),
.B1(n_1057),
.B2(n_1055),
.Y(n_1205)
);

BUFx2_ASAP7_75t_R g1206 ( 
.A(n_1085),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1099),
.Y(n_1207)
);

INVx4_ASAP7_75t_SL g1208 ( 
.A(n_1099),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1099),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1099),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1049),
.A2(n_831),
.B1(n_859),
.B2(n_964),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1013),
.Y(n_1212)
);

OAI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1049),
.A2(n_685),
.B1(n_964),
.B2(n_656),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1026),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1086),
.Y(n_1215)
);

NAND2x1_ASAP7_75t_L g1216 ( 
.A(n_1071),
.B(n_913),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1098),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1005),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1100),
.A2(n_980),
.B1(n_961),
.B2(n_970),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1063),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1100),
.A2(n_980),
.B1(n_961),
.B2(n_970),
.Y(n_1221)
);

NAND2x1p5_ASAP7_75t_L g1222 ( 
.A(n_1052),
.B(n_1071),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1026),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_1098),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1005),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1026),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1100),
.A2(n_831),
.B1(n_859),
.B2(n_964),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1086),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1176),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1192),
.B(n_1148),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1227),
.A2(n_1121),
.B1(n_1211),
.B2(n_1149),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1146),
.Y(n_1232)
);

INVx6_ASAP7_75t_L g1233 ( 
.A(n_1208),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1150),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1124),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1184),
.Y(n_1236)
);

INVx5_ASAP7_75t_L g1237 ( 
.A(n_1198),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1192),
.B(n_1148),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1219),
.B(n_1221),
.Y(n_1239)
);

OR2x6_ASAP7_75t_L g1240 ( 
.A(n_1216),
.B(n_1138),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1181),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1144),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1215),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1185),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1123),
.B(n_1135),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1124),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_1131),
.Y(n_1247)
);

AOI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1181),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1124),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1171),
.B(n_1167),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1125),
.A2(n_1123),
.B1(n_1154),
.B2(n_1163),
.Y(n_1251)
);

BUFx4f_ASAP7_75t_SL g1252 ( 
.A(n_1141),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1150),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1228),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1135),
.B(n_1177),
.Y(n_1255)
);

INVxp67_ASAP7_75t_SL g1256 ( 
.A(n_1172),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1185),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1191),
.B(n_1132),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1138),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1196),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1160),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1143),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1138),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_1175),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1145),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1182),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1173),
.B(n_1169),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1151),
.B(n_1177),
.Y(n_1268)
);

AO21x2_ASAP7_75t_L g1269 ( 
.A1(n_1120),
.A2(n_1202),
.B(n_1183),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_1142),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1222),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1159),
.B(n_1126),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1125),
.B(n_1151),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1161),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1155),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1122),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1128),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1214),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1194),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1223),
.B(n_1226),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1194),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1139),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1208),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1137),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1183),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1194),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1183),
.B(n_1140),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1170),
.B(n_1134),
.Y(n_1288)
);

AO21x2_ASAP7_75t_L g1289 ( 
.A1(n_1213),
.A2(n_1190),
.B(n_1195),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1131),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1136),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1156),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1162),
.B(n_1129),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1209),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1178),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1209),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1210),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1164),
.B(n_1225),
.Y(n_1298)
);

NAND2x1p5_ASAP7_75t_L g1299 ( 
.A(n_1132),
.B(n_1207),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1186),
.B(n_1187),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1287),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1232),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1287),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1278),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1273),
.B(n_1200),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1237),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1231),
.A2(n_1189),
.B1(n_1168),
.B2(n_1225),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1273),
.B(n_1179),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1245),
.B(n_1218),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1259),
.B(n_1208),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1244),
.B(n_1218),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1262),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1272),
.A2(n_1168),
.B1(n_1166),
.B2(n_1197),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1265),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1257),
.B(n_1188),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1257),
.B(n_1193),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1268),
.B(n_1212),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1255),
.B(n_1212),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1241),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1299),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1255),
.B(n_1236),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1268),
.B(n_1199),
.Y(n_1322)
);

AOI221xp5_ASAP7_75t_L g1323 ( 
.A1(n_1239),
.A2(n_1174),
.B1(n_1180),
.B2(n_1166),
.C(n_1147),
.Y(n_1323)
);

NOR2x1_ASAP7_75t_L g1324 ( 
.A(n_1242),
.B(n_1127),
.Y(n_1324)
);

NOR2x1_ASAP7_75t_L g1325 ( 
.A(n_1242),
.B(n_1127),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1256),
.B(n_1220),
.Y(n_1326)
);

AOI21xp33_ASAP7_75t_L g1327 ( 
.A1(n_1251),
.A2(n_1203),
.B(n_1204),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1279),
.B(n_1157),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1281),
.B(n_1153),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1281),
.B(n_1153),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1286),
.B(n_1269),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1286),
.B(n_1153),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1269),
.B(n_1153),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1275),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1275),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1269),
.B(n_1220),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1241),
.B(n_1201),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_L g1338 ( 
.A(n_1323),
.B(n_1293),
.C(n_1267),
.Y(n_1338)
);

NAND3xp33_ASAP7_75t_L g1339 ( 
.A(n_1323),
.B(n_1261),
.C(n_1250),
.Y(n_1339)
);

AOI221xp5_ASAP7_75t_L g1340 ( 
.A1(n_1302),
.A2(n_1264),
.B1(n_1243),
.B2(n_1254),
.C(n_1266),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1321),
.B(n_1230),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1313),
.B(n_1247),
.Y(n_1342)
);

NAND3xp33_ASAP7_75t_L g1343 ( 
.A(n_1307),
.B(n_1284),
.C(n_1274),
.Y(n_1343)
);

OAI221xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1313),
.A2(n_1298),
.B1(n_1290),
.B2(n_1205),
.C(n_1242),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1302),
.A2(n_1233),
.B1(n_1283),
.B2(n_1270),
.Y(n_1345)
);

AOI221xp5_ASAP7_75t_L g1346 ( 
.A1(n_1305),
.A2(n_1292),
.B1(n_1291),
.B2(n_1282),
.C(n_1294),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1312),
.Y(n_1347)
);

AOI221xp5_ASAP7_75t_L g1348 ( 
.A1(n_1327),
.A2(n_1291),
.B1(n_1297),
.B2(n_1296),
.C(n_1294),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1321),
.B(n_1238),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1309),
.B(n_1238),
.Y(n_1350)
);

NAND3xp33_ASAP7_75t_L g1351 ( 
.A(n_1326),
.B(n_1288),
.C(n_1297),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1309),
.B(n_1295),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1310),
.B(n_1258),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1329),
.B(n_1285),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1308),
.B(n_1147),
.Y(n_1355)
);

NAND3xp33_ASAP7_75t_L g1356 ( 
.A(n_1326),
.B(n_1288),
.C(n_1296),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1329),
.B(n_1285),
.Y(n_1357)
);

NOR3xp33_ASAP7_75t_L g1358 ( 
.A(n_1324),
.B(n_1248),
.C(n_1260),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1308),
.B(n_1295),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1312),
.Y(n_1360)
);

NAND3xp33_ASAP7_75t_L g1361 ( 
.A(n_1324),
.B(n_1300),
.C(n_1229),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1310),
.A2(n_1233),
.B1(n_1289),
.B2(n_1283),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1318),
.B(n_1276),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_L g1364 ( 
.A(n_1325),
.B(n_1300),
.C(n_1229),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1329),
.B(n_1234),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1330),
.B(n_1234),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1311),
.B(n_1276),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1330),
.B(n_1253),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1311),
.B(n_1277),
.Y(n_1369)
);

OAI221xp5_ASAP7_75t_SL g1370 ( 
.A1(n_1337),
.A2(n_1322),
.B1(n_1331),
.B2(n_1317),
.C(n_1240),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1322),
.B(n_1280),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1317),
.A2(n_1233),
.B1(n_1206),
.B2(n_1283),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1332),
.B(n_1263),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1328),
.B(n_1271),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1310),
.B(n_1258),
.Y(n_1375)
);

OAI221xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1337),
.A2(n_1240),
.B1(n_1246),
.B2(n_1249),
.C(n_1235),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1371),
.B(n_1301),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1353),
.B(n_1306),
.Y(n_1378)
);

NAND2x1p5_ASAP7_75t_L g1379 ( 
.A(n_1375),
.B(n_1306),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1347),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1360),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1363),
.B(n_1303),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1373),
.B(n_1333),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1360),
.Y(n_1384)
);

AOI33xp33_ASAP7_75t_L g1385 ( 
.A1(n_1340),
.A2(n_1316),
.A3(n_1315),
.B1(n_1314),
.B2(n_1335),
.B3(n_1334),
.Y(n_1385)
);

INVx4_ASAP7_75t_L g1386 ( 
.A(n_1365),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1367),
.Y(n_1387)
);

INVxp33_ASAP7_75t_L g1388 ( 
.A(n_1355),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1338),
.B(n_1133),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1369),
.B(n_1359),
.Y(n_1390)
);

NOR2xp67_ASAP7_75t_L g1391 ( 
.A(n_1361),
.B(n_1319),
.Y(n_1391)
);

INVxp67_ASAP7_75t_L g1392 ( 
.A(n_1361),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1354),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1357),
.B(n_1320),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1338),
.B(n_1252),
.Y(n_1395)
);

AND2x4_ASAP7_75t_SL g1396 ( 
.A(n_1374),
.B(n_1310),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1357),
.B(n_1333),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1351),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1342),
.B(n_1165),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1352),
.B(n_1370),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1351),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1356),
.B(n_1304),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1356),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1341),
.B(n_1336),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1349),
.B(n_1350),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1391),
.A2(n_1339),
.B(n_1364),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1386),
.B(n_1365),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1398),
.B(n_1346),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1391),
.B(n_1364),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1398),
.B(n_1348),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1401),
.B(n_1358),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1380),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1393),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1401),
.B(n_1403),
.Y(n_1414)
);

INVxp67_ASAP7_75t_L g1415 ( 
.A(n_1389),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1396),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1403),
.B(n_1366),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1388),
.B(n_1339),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1392),
.B(n_1368),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1380),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1393),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1381),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1381),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1384),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1392),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1384),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1402),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1396),
.B(n_1362),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1402),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1393),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1394),
.B(n_1320),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1377),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1394),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1412),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1412),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1428),
.B(n_1394),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1425),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1418),
.B(n_1400),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1428),
.B(n_1404),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1416),
.B(n_1404),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1416),
.B(n_1383),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1408),
.B(n_1400),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1408),
.B(n_1385),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1420),
.Y(n_1444)
);

INVxp67_ASAP7_75t_L g1445 ( 
.A(n_1411),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1420),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1415),
.B(n_1395),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1433),
.B(n_1383),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1414),
.B(n_1382),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1422),
.Y(n_1450)
);

INVxp67_ASAP7_75t_SL g1451 ( 
.A(n_1409),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1414),
.B(n_1382),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1422),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1423),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1413),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1423),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1424),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1432),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1411),
.B(n_1387),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1409),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1424),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1410),
.B(n_1390),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1410),
.A2(n_1344),
.B(n_1399),
.C(n_1343),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1413),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1433),
.B(n_1397),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1419),
.B(n_1141),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1417),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1431),
.B(n_1397),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1426),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1419),
.B(n_1417),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_SL g1471 ( 
.A(n_1406),
.B(n_1376),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1426),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1406),
.B(n_1427),
.Y(n_1473)
);

INVxp67_ASAP7_75t_SL g1474 ( 
.A(n_1409),
.Y(n_1474)
);

OAI21xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1407),
.A2(n_1405),
.B(n_1390),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1438),
.A2(n_1343),
.B1(n_1409),
.B2(n_1429),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1460),
.B(n_1413),
.Y(n_1477)
);

AOI22x1_ASAP7_75t_L g1478 ( 
.A1(n_1437),
.A2(n_1378),
.B1(n_1379),
.B2(n_1130),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1460),
.B(n_1421),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1451),
.B(n_1421),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_1458),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1474),
.B(n_1421),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1434),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1436),
.B(n_1430),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1455),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1455),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1464),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1434),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1464),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1435),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1473),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1435),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1445),
.B(n_1427),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1444),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1436),
.B(n_1430),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1439),
.B(n_1430),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1444),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1446),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_1447),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1471),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1449),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1449),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1452),
.Y(n_1503)
);

INVx3_ASAP7_75t_SL g1504 ( 
.A(n_1452),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1466),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1446),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1450),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1450),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1442),
.B(n_1429),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1453),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1500),
.A2(n_1463),
.B(n_1443),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1477),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1476),
.A2(n_1462),
.B1(n_1467),
.B2(n_1470),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1500),
.A2(n_1475),
.B(n_1459),
.C(n_1372),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1476),
.A2(n_1439),
.B1(n_1440),
.B2(n_1441),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1480),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1499),
.B(n_1468),
.Y(n_1517)
);

OAI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1491),
.A2(n_1345),
.B1(n_1379),
.B2(n_1378),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1491),
.B(n_1468),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1510),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1510),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1499),
.A2(n_1509),
.B(n_1481),
.C(n_1505),
.Y(n_1522)
);

AOI21xp33_ASAP7_75t_L g1523 ( 
.A1(n_1481),
.A2(n_1454),
.B(n_1453),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1483),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1509),
.A2(n_1456),
.B1(n_1472),
.B2(n_1461),
.C(n_1457),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1504),
.B(n_1440),
.Y(n_1526)
);

OAI211xp5_ASAP7_75t_L g1527 ( 
.A1(n_1493),
.A2(n_1472),
.B(n_1469),
.C(n_1454),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1478),
.A2(n_1379),
.B1(n_1378),
.B2(n_1441),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1480),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1483),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1504),
.B(n_1448),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1488),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1488),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1490),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1480),
.Y(n_1535)
);

NOR2x1_ASAP7_75t_L g1536 ( 
.A(n_1522),
.B(n_1490),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1517),
.B(n_1504),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1512),
.Y(n_1538)
);

INVxp33_ASAP7_75t_L g1539 ( 
.A(n_1526),
.Y(n_1539)
);

INVx4_ASAP7_75t_L g1540 ( 
.A(n_1516),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1512),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1519),
.B(n_1504),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1511),
.B(n_1501),
.Y(n_1543)
);

INVx1_ASAP7_75t_SL g1544 ( 
.A(n_1531),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1520),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1516),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1515),
.B(n_1529),
.Y(n_1547)
);

NOR3xp33_ASAP7_75t_L g1548 ( 
.A(n_1522),
.B(n_1505),
.C(n_1493),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1513),
.B(n_1501),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1514),
.B(n_1502),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1521),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1529),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1535),
.B(n_1502),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1535),
.B(n_1503),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1514),
.B(n_1503),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1544),
.B(n_1525),
.Y(n_1556)
);

OAI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1548),
.A2(n_1523),
.B1(n_1528),
.B2(n_1478),
.C(n_1527),
.Y(n_1557)
);

O2A1O1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1550),
.A2(n_1518),
.B(n_1534),
.C(n_1524),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1543),
.A2(n_1518),
.B1(n_1532),
.B2(n_1530),
.Y(n_1559)
);

AOI221xp5_ASAP7_75t_L g1560 ( 
.A1(n_1555),
.A2(n_1533),
.B1(n_1508),
.B2(n_1492),
.C(n_1494),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1538),
.Y(n_1561)
);

AOI211xp5_ASAP7_75t_L g1562 ( 
.A1(n_1555),
.A2(n_1482),
.B(n_1480),
.C(n_1477),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1546),
.B(n_1484),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1536),
.A2(n_1448),
.B1(n_1465),
.B2(n_1484),
.Y(n_1564)
);

OAI31xp33_ASAP7_75t_L g1565 ( 
.A1(n_1549),
.A2(n_1482),
.A3(n_1480),
.B(n_1477),
.Y(n_1565)
);

NAND5xp2_ASAP7_75t_SL g1566 ( 
.A(n_1565),
.B(n_1547),
.C(n_1554),
.D(n_1539),
.E(n_1537),
.Y(n_1566)
);

NOR2x1p5_ASAP7_75t_L g1567 ( 
.A(n_1556),
.B(n_1542),
.Y(n_1567)
);

AOI211x1_ASAP7_75t_L g1568 ( 
.A1(n_1557),
.A2(n_1547),
.B(n_1551),
.C(n_1554),
.Y(n_1568)
);

NOR3xp33_ASAP7_75t_L g1569 ( 
.A(n_1558),
.B(n_1545),
.C(n_1540),
.Y(n_1569)
);

NOR2x1p5_ASAP7_75t_L g1570 ( 
.A(n_1563),
.B(n_1553),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1561),
.B(n_1539),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_L g1572 ( 
.A(n_1560),
.B(n_1541),
.C(n_1553),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1559),
.B(n_1540),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1564),
.B(n_1540),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1571),
.B(n_1562),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1574),
.B(n_1552),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1570),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1569),
.B(n_1552),
.Y(n_1578)
);

OAI211xp5_ASAP7_75t_SL g1579 ( 
.A1(n_1573),
.A2(n_1508),
.B(n_1492),
.C(n_1494),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1576),
.A2(n_1567),
.B1(n_1572),
.B2(n_1566),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1577),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1578),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1575),
.B(n_1482),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1579),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1577),
.Y(n_1585)
);

NAND3x1_ASAP7_75t_L g1586 ( 
.A(n_1580),
.B(n_1568),
.C(n_1479),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1583),
.Y(n_1587)
);

NOR2x1_ASAP7_75t_SL g1588 ( 
.A(n_1581),
.B(n_1479),
.Y(n_1588)
);

NAND3xp33_ASAP7_75t_L g1589 ( 
.A(n_1584),
.B(n_1479),
.C(n_1497),
.Y(n_1589)
);

OAI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1585),
.A2(n_1497),
.B1(n_1498),
.B2(n_1506),
.C(n_1507),
.Y(n_1590)
);

NOR2xp67_ASAP7_75t_L g1591 ( 
.A(n_1589),
.B(n_1583),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1587),
.B(n_1582),
.Y(n_1592)
);

XNOR2xp5_ASAP7_75t_L g1593 ( 
.A(n_1586),
.B(n_1217),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1592),
.Y(n_1594)
);

NAND5xp2_ASAP7_75t_L g1595 ( 
.A(n_1594),
.B(n_1593),
.C(n_1590),
.D(n_1591),
.E(n_1588),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1595),
.B(n_1498),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1596),
.A2(n_1224),
.B(n_1217),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1597),
.A2(n_1224),
.B(n_1506),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1598),
.B(n_1507),
.Y(n_1599)
);

OAI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1599),
.A2(n_1487),
.B1(n_1486),
.B2(n_1489),
.Y(n_1600)
);

AOI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1600),
.A2(n_1486),
.B1(n_1485),
.B2(n_1484),
.C(n_1495),
.Y(n_1601)
);

AOI211xp5_ASAP7_75t_L g1602 ( 
.A1(n_1601),
.A2(n_1485),
.B(n_1495),
.C(n_1496),
.Y(n_1602)
);


endmodule