module fake_jpeg_32080_n_183 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_183);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_43),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_21),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_79),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_0),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_84),
.Y(n_90)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp67_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_3),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_4),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_75),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_SL g89 ( 
.A(n_80),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_56),
.B1(n_73),
.B2(n_71),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_62),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_60),
.B1(n_65),
.B2(n_75),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_56),
.B1(n_73),
.B2(n_71),
.Y(n_96)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_108),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_53),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_115),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_59),
.B1(n_66),
.B2(n_60),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_116),
.B1(n_5),
.B2(n_6),
.Y(n_131)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_113),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_67),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_77),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_58),
.B1(n_70),
.B2(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_111),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_91),
.B1(n_58),
.B2(n_76),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_91),
.B(n_57),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_31),
.B(n_34),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_55),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_54),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_127),
.B(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_4),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_91),
.C(n_27),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_136),
.C(n_123),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_137),
.B1(n_8),
.B2(n_9),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_7),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_132),
.B(n_13),
.Y(n_144)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_29),
.C(n_49),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_142),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_133),
.B1(n_135),
.B2(n_44),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_149),
.B1(n_157),
.B2(n_158),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_35),
.B(n_47),
.C(n_16),
.D(n_19),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_148),
.B(n_153),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_14),
.B1(n_15),
.B2(n_20),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_23),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_26),
.Y(n_155)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_36),
.B(n_38),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_150),
.B1(n_154),
.B2(n_120),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_161),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_160),
.B(n_165),
.C(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_173),
.A2(n_174),
.B1(n_159),
.B2(n_171),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_167),
.C(n_163),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_166),
.Y(n_176)
);

OAI21x1_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_164),
.B(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_155),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_158),
.B(n_40),
.Y(n_179)
);

AOI321xp33_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_39),
.A3(n_45),
.B1(n_46),
.B2(n_51),
.C(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_145),
.B(n_146),
.Y(n_182)
);

BUFx24_ASAP7_75t_SL g183 ( 
.A(n_182),
.Y(n_183)
);


endmodule