module fake_jpeg_18807_n_260 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_38),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_44),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_54),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_49),
.B(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_31),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_26),
.B1(n_33),
.B2(n_18),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_58),
.B1(n_65),
.B2(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_67),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_26),
.B1(n_33),
.B2(n_18),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_26),
.B1(n_28),
.B2(n_19),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_45),
.B1(n_28),
.B2(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_20),
.B1(n_31),
.B2(n_27),
.Y(n_65)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_40),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_27),
.B1(n_20),
.B2(n_29),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_74),
.B(n_100),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_21),
.B1(n_32),
.B2(n_29),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_75),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_78),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_77),
.A2(n_5),
.B1(n_6),
.B2(n_10),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_17),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_45),
.B1(n_40),
.B2(n_37),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_84),
.B1(n_87),
.B2(n_93),
.Y(n_107)
);

BUFx2_ASAP7_75t_SL g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_21),
.B1(n_32),
.B2(n_45),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_82),
.A2(n_97),
.B(n_99),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_51),
.B1(n_46),
.B2(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_35),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_105),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_23),
.B1(n_22),
.B2(n_30),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_90),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_35),
.C(n_34),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_25),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_30),
.B1(n_22),
.B2(n_34),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_67),
.A2(n_22),
.B1(n_34),
.B2(n_30),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_96),
.B1(n_102),
.B2(n_0),
.Y(n_119)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_35),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_30),
.B(n_40),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_35),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_40),
.B1(n_11),
.B2(n_15),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_43),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_66),
.B1(n_40),
.B2(n_43),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_121),
.B1(n_124),
.B2(n_129),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_40),
.B1(n_37),
.B2(n_43),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_113),
.B1(n_116),
.B2(n_119),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_43),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_99),
.B1(n_91),
.B2(n_71),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_60),
.B(n_62),
.C(n_25),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_131),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_76),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_0),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_125),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_86),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

AO22x1_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_72),
.B(n_1),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_130),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_75),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_4),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_82),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_SL g142 ( 
.A1(n_133),
.A2(n_102),
.B(n_94),
.Y(n_142)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_145),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_140),
.A2(n_144),
.B(n_112),
.Y(n_171)
);

OAI22x1_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_126),
.B1(n_116),
.B2(n_119),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_142),
.B1(n_107),
.B2(n_110),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_108),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_148),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_97),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_121),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_95),
.B1(n_88),
.B2(n_92),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_152),
.B1(n_154),
.B2(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_115),
.A2(n_92),
.B1(n_73),
.B2(n_98),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_107),
.A2(n_104),
.B1(n_101),
.B2(n_103),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_104),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_156),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_101),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_101),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_120),
.Y(n_180)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_160),
.Y(n_170)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_118),
.C(n_109),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_165),
.C(n_172),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_126),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_168),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_140),
.C(n_160),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_123),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_149),
.B1(n_137),
.B2(n_134),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_177),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_150),
.C(n_139),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_154),
.B1(n_158),
.B2(n_138),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_159),
.B(n_128),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_176),
.B(n_145),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_124),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_136),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_120),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_164),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_131),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_125),
.C(n_11),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_187),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_188),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_138),
.B1(n_149),
.B2(n_144),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_176),
.B(n_145),
.Y(n_189)
);

AOI321xp33_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_177),
.A3(n_169),
.B1(n_125),
.B2(n_182),
.C(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_106),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_193),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_106),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_196),
.A2(n_167),
.B1(n_199),
.B2(n_197),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_175),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_198),
.B(n_199),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_151),
.B1(n_146),
.B2(n_136),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_175),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_161),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_183),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_209),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_205),
.B(n_215),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_206),
.A2(n_198),
.B1(n_196),
.B2(n_190),
.Y(n_220)
);

NOR2x1_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_163),
.Y(n_207)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_162),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_201),
.B(n_165),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_213),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_168),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_171),
.C(n_163),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_217),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_182),
.C(n_179),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_218),
.B(n_103),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_222),
.Y(n_236)
);

INVxp33_ASAP7_75t_SL g221 ( 
.A(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_221),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_192),
.B1(n_187),
.B2(n_186),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_189),
.B(n_200),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_225),
.B(n_207),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_202),
.B1(n_167),
.B2(n_12),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_231),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_10),
.B(n_11),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_209),
.Y(n_240)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_210),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_237),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_218),
.B(n_215),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_223),
.B(n_219),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_213),
.C(n_205),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_226),
.B(n_204),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_238),
.B(n_240),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_235),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_233),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_219),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_234),
.A2(n_221),
.B(n_217),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_248),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_242),
.B(n_239),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_250),
.A2(n_251),
.B(n_232),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_236),
.Y(n_251)
);

AOI21x1_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_232),
.B(n_243),
.Y(n_252)
);

OAI21x1_ASAP7_75t_SL g256 ( 
.A1(n_252),
.A2(n_247),
.B(n_237),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_244),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_255),
.A2(n_256),
.B(n_12),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_253),
.C(n_103),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_258),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_14),
.Y(n_260)
);


endmodule