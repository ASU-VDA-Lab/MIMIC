module fake_jpeg_2214_n_83 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_37),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_0),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_31),
.B1(n_26),
.B2(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_33),
.B(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_1),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_27),
.B1(n_29),
.B2(n_3),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_1),
.Y(n_52)
);

A2O1A1O1Ixp25_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_29),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

AOI32xp33_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_45),
.A3(n_29),
.B1(n_27),
.B2(n_4),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_61),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_5),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_69),
.B1(n_12),
.B2(n_15),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_46),
.B1(n_45),
.B2(n_57),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_64),
.B1(n_66),
.B2(n_63),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.C(n_11),
.Y(n_74)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_6),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_74),
.B1(n_75),
.B2(n_17),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_8),
.B(n_9),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_72),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_76),
.B(n_73),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_18),
.C(n_19),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_20),
.C(n_21),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_22),
.Y(n_83)
);


endmodule