module real_jpeg_29743_n_17 (n_8, n_0, n_93, n_95, n_2, n_91, n_10, n_9, n_12, n_92, n_97, n_6, n_11, n_14, n_90, n_7, n_3, n_5, n_4, n_98, n_94, n_1, n_96, n_89, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_93;
input n_95;
input n_2;
input n_91;
input n_10;
input n_9;
input n_12;
input n_92;
input n_97;
input n_6;
input n_11;
input n_14;
input n_90;
input n_7;
input n_3;
input n_5;
input n_4;
input n_98;
input n_94;
input n_1;
input n_96;
input n_89;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_1),
.B(n_26),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_1),
.B(n_26),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_3),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_3),
.B(n_84),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_4),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_5),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_6),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_6),
.B(n_58),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_7),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

FAx1_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_18),
.CI(n_22),
.CON(n_17),
.SN(n_17)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_10),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_11),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_11),
.B(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_12),
.B(n_50),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_12),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_13),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_13),
.B(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_14),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_15),
.B(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_16),
.B(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_20),
.B(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_83),
.B(n_86),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_78),
.B(n_82),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_29),
.B(n_74),
.C(n_77),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_27),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_73),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_35),
.B(n_72),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_33),
.B(n_76),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_33),
.B(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_67),
.B(n_71),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B(n_66),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_61),
.B(n_65),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_57),
.B(n_60),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_52),
.B(n_56),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_48),
.B(n_51),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_59),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_62),
.B(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_81),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_89),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_90),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_91),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_92),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_93),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_94),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_95),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_96),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_97),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_98),
.Y(n_76)
);


endmodule