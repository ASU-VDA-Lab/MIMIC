module fake_jpeg_30713_n_547 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_547);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_547;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_6),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_54),
.Y(n_158)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_31),
.B(n_10),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_66),
.Y(n_108)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_10),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_69),
.B(n_84),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

CKINVDCx6p67_ASAP7_75t_R g142 ( 
.A(n_77),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_25),
.B(n_9),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_78),
.B(n_85),
.Y(n_148)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_9),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_27),
.B(n_11),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_27),
.B(n_8),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_89),
.B(n_94),
.Y(n_165)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_32),
.B(n_8),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_32),
.B(n_12),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_45),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_36),
.B(n_12),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_45),
.Y(n_146)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

BUFx4f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

BUFx8_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_106),
.B(n_146),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_56),
.B(n_17),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_109),
.B(n_7),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_61),
.A2(n_51),
.B1(n_36),
.B2(n_40),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_111),
.A2(n_118),
.B1(n_127),
.B2(n_14),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_51),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_113),
.B(n_157),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_77),
.A2(n_87),
.B1(n_71),
.B2(n_88),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_117),
.A2(n_128),
.B1(n_130),
.B2(n_135),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_63),
.A2(n_40),
.B1(n_29),
.B2(n_46),
.Y(n_118)
);

AND2x4_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_24),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_24),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_65),
.A2(n_70),
.B1(n_68),
.B2(n_59),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_77),
.A2(n_43),
.B1(n_41),
.B2(n_49),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_86),
.B1(n_82),
.B2(n_83),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_53),
.A2(n_43),
.B1(n_41),
.B2(n_49),
.Y(n_135)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_57),
.Y(n_156)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_101),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_90),
.A2(n_43),
.B1(n_41),
.B2(n_49),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_128),
.B1(n_135),
.B2(n_117),
.Y(n_199)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_64),
.Y(n_163)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_60),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_132),
.A2(n_52),
.B1(n_62),
.B2(n_75),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_169),
.A2(n_181),
.B1(n_197),
.B2(n_211),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_171),
.B(n_190),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_142),
.Y(n_172)
);

INVx11_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_76),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_174),
.B(n_178),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_132),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_175),
.B(n_205),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_180),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_143),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_140),
.A2(n_92),
.B1(n_74),
.B2(n_73),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_182),
.A2(n_199),
.B1(n_202),
.B2(n_204),
.Y(n_269)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_142),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_224),
.Y(n_241)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_185),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_187),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_189),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_162),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_108),
.B(n_95),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_191),
.Y(n_235)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_192),
.Y(n_249)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_106),
.A2(n_46),
.B1(n_28),
.B2(n_39),
.Y(n_195)
);

A2O1A1O1Ixp25_ASAP7_75t_L g266 ( 
.A1(n_195),
.A2(n_206),
.B(n_218),
.C(n_220),
.D(n_14),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_168),
.A2(n_54),
.B1(n_99),
.B2(n_103),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_134),
.Y(n_198)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_198),
.Y(n_271)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_200),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_152),
.B1(n_149),
.B2(n_136),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_123),
.A2(n_102),
.B1(n_50),
.B2(n_21),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_203),
.Y(n_281)
);

AO22x2_ASAP7_75t_L g204 ( 
.A1(n_120),
.A2(n_41),
.B1(n_50),
.B2(n_21),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_108),
.B(n_50),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_109),
.A2(n_50),
.B1(n_21),
.B2(n_19),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_207),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_148),
.B(n_50),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_208),
.B(n_225),
.Y(n_253)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_137),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_209),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_21),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_210),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_139),
.A2(n_21),
.B1(n_19),
.B2(n_2),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_114),
.Y(n_212)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_212),
.Y(n_276)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_116),
.Y(n_213)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_112),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_107),
.Y(n_215)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_148),
.B(n_19),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_221),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_129),
.A2(n_19),
.B1(n_12),
.B2(n_2),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_151),
.A2(n_141),
.B(n_138),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_125),
.B(n_13),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_159),
.A2(n_123),
.B1(n_124),
.B2(n_152),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_222),
.A2(n_223),
.B1(n_7),
.B2(n_17),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_124),
.A2(n_19),
.B1(n_13),
.B2(n_2),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_130),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_125),
.Y(n_226)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_115),
.B(n_7),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_151),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_228),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_131),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_229),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

BUFx16f_ASAP7_75t_L g272 ( 
.A(n_230),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_232),
.A2(n_256),
.B1(n_258),
.B2(n_178),
.Y(n_294)
);

AND2x6_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_237),
.B(n_255),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_186),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_242),
.B(n_261),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_263),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_191),
.B(n_225),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_275),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_170),
.B(n_158),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_201),
.A2(n_136),
.B1(n_149),
.B2(n_150),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_224),
.A2(n_150),
.B1(n_158),
.B2(n_164),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_207),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_177),
.B(n_161),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_195),
.B(n_131),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_270),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_266),
.B(n_173),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_210),
.B(n_119),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_217),
.B(n_160),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_274),
.B(n_190),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_191),
.B(n_160),
.Y(n_275)
);

OA22x2_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_218),
.B1(n_206),
.B2(n_216),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_196),
.B1(n_222),
.B2(n_182),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_283),
.A2(n_296),
.B1(n_298),
.B2(n_299),
.Y(n_338)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_280),
.Y(n_286)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_243),
.A2(n_229),
.B1(n_193),
.B2(n_172),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_287),
.A2(n_291),
.B1(n_294),
.B2(n_324),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_171),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_288),
.B(n_290),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_171),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_289),
.B(n_317),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_238),
.B(n_204),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_257),
.A2(n_187),
.B1(n_173),
.B2(n_220),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_239),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_292),
.B(n_304),
.Y(n_334)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_293),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_233),
.Y(n_295)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_279),
.B1(n_235),
.B2(n_265),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_235),
.A2(n_204),
.B1(n_198),
.B2(n_194),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_300),
.Y(n_353)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_275),
.A2(n_204),
.B(n_176),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_302),
.A2(n_327),
.B(n_234),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_238),
.B(n_189),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_253),
.B(n_180),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_305),
.B(n_309),
.Y(n_347)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_306),
.Y(n_358)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_307),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_321),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_255),
.B(n_179),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_256),
.A2(n_215),
.B1(n_228),
.B2(n_226),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_310),
.A2(n_323),
.B1(n_328),
.B2(n_267),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_253),
.B(n_200),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_311),
.B(n_312),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_241),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_249),
.B(n_185),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_313),
.B(n_326),
.Y(n_364)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_254),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_316),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_248),
.B(n_212),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_272),
.Y(n_339)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_250),
.Y(n_319)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_251),
.Y(n_320)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_248),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_272),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_330),
.Y(n_343)
);

OA22x2_ASAP7_75t_L g323 ( 
.A1(n_232),
.A2(n_183),
.B1(n_219),
.B2(n_214),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_258),
.A2(n_230),
.B1(n_188),
.B2(n_4),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_248),
.B(n_0),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_236),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_249),
.B(n_6),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_266),
.B(n_0),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_237),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_272),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_297),
.A2(n_236),
.B(n_242),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_331),
.A2(n_339),
.B(n_349),
.Y(n_387)
);

AOI32xp33_ASAP7_75t_L g333 ( 
.A1(n_303),
.A2(n_234),
.A3(n_261),
.B1(n_268),
.B2(n_278),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_333),
.B(n_298),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_337),
.A2(n_341),
.B(n_346),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_302),
.A2(n_262),
.B(n_240),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_329),
.A2(n_262),
.B(n_240),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_348),
.B(n_362),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_290),
.A2(n_281),
.B(n_245),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_318),
.A2(n_281),
.B(n_233),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_350),
.A2(n_355),
.B(n_357),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_285),
.B(n_276),
.C(n_271),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_361),
.C(n_370),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_318),
.A2(n_276),
.B(n_231),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_309),
.A2(n_231),
.B(n_257),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_312),
.A2(n_285),
.B(n_288),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_360),
.A2(n_369),
.B(n_301),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_305),
.B(n_271),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_289),
.B(n_259),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_365),
.A2(n_324),
.B1(n_329),
.B2(n_298),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_311),
.B(n_259),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_368),
.B(n_260),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_321),
.A2(n_327),
.B(n_317),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_304),
.B(n_296),
.C(n_292),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_352),
.A2(n_283),
.B1(n_328),
.B2(n_299),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_372),
.A2(n_373),
.B1(n_393),
.B2(n_400),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_341),
.A2(n_310),
.B1(n_294),
.B2(n_298),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_284),
.C(n_327),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_374),
.B(n_395),
.Y(n_413)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_363),
.Y(n_375)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_376),
.A2(n_385),
.B1(n_390),
.B2(n_394),
.Y(n_408)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_336),
.Y(n_377)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_377),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_335),
.B(n_329),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_379),
.B(n_381),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_343),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_382),
.A2(n_406),
.B1(n_360),
.B2(n_369),
.Y(n_417)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_336),
.Y(n_383)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_383),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_334),
.B(n_286),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_388),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_338),
.A2(n_323),
.B1(n_325),
.B2(n_300),
.Y(n_385)
);

OAI21xp33_ASAP7_75t_L g386 ( 
.A1(n_332),
.A2(n_316),
.B(n_322),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_SL g423 ( 
.A(n_386),
.B(n_404),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_323),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_364),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_389),
.B(n_401),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_338),
.A2(n_323),
.B1(n_293),
.B2(n_316),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_397),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_337),
.A2(n_254),
.B1(n_320),
.B2(n_319),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_365),
.A2(n_247),
.B1(n_246),
.B2(n_306),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_335),
.B(n_330),
.Y(n_396)
);

XNOR2x1_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_361),
.Y(n_422)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_353),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_315),
.C(n_251),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_398),
.B(n_354),
.C(n_340),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_339),
.A2(n_247),
.B1(n_246),
.B2(n_314),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_399),
.A2(n_345),
.B1(n_342),
.B2(n_344),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_351),
.A2(n_247),
.B1(n_246),
.B2(n_307),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_346),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_403),
.B(n_340),
.Y(n_407)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_331),
.B(n_6),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_405),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_368),
.A2(n_260),
.B1(n_1),
.B2(n_0),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_407),
.B(n_422),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_429),
.C(n_431),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_410),
.A2(n_412),
.B1(n_427),
.B2(n_393),
.Y(n_438)
);

OAI22x1_ASAP7_75t_L g412 ( 
.A1(n_373),
.A2(n_355),
.B1(n_350),
.B2(n_357),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_417),
.A2(n_385),
.B1(n_394),
.B2(n_372),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_380),
.A2(n_349),
.B(n_344),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_419),
.A2(n_412),
.B(n_423),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_379),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_425),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_384),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_426),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_376),
.A2(n_348),
.B1(n_345),
.B2(n_371),
.Y(n_427)
);

OA22x2_ASAP7_75t_L g428 ( 
.A1(n_390),
.A2(n_359),
.B1(n_371),
.B2(n_358),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_433),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_378),
.B(n_367),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_380),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_430),
.B(n_432),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_378),
.B(n_402),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_400),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_381),
.A2(n_342),
.B1(n_366),
.B2(n_358),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_367),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_434),
.B(n_374),
.C(n_398),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_401),
.A2(n_405),
.B(n_395),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_437),
.A2(n_392),
.B(n_387),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_438),
.A2(n_420),
.B1(n_419),
.B2(n_408),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_409),
.Y(n_471)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_418),
.Y(n_441)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_441),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_404),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_450),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_444),
.A2(n_356),
.B(n_359),
.Y(n_484)
);

OAI21xp33_ASAP7_75t_L g447 ( 
.A1(n_436),
.A2(n_387),
.B(n_396),
.Y(n_447)
);

OAI21xp33_ASAP7_75t_L g477 ( 
.A1(n_447),
.A2(n_413),
.B(n_422),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_414),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_448),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_449),
.A2(n_408),
.B1(n_427),
.B2(n_420),
.Y(n_475)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_403),
.C(n_392),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_458),
.C(n_413),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_452),
.B(n_437),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_415),
.B(n_421),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_453),
.B(n_455),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_377),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_454),
.B(n_464),
.Y(n_486)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_416),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_415),
.B(n_397),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_457),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_429),
.B(n_406),
.C(n_391),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_411),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_459),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_410),
.Y(n_461)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_461),
.Y(n_467)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_416),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_462),
.B(n_463),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_435),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_435),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_465),
.B(n_477),
.Y(n_488)
);

INVxp33_ASAP7_75t_SL g470 ( 
.A(n_443),
.Y(n_470)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_470),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_478),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_474),
.A2(n_459),
.B1(n_441),
.B2(n_450),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_475),
.A2(n_445),
.B1(n_454),
.B2(n_446),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_407),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_480),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_451),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_439),
.B(n_434),
.C(n_428),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_483),
.C(n_458),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_449),
.A2(n_383),
.B1(n_428),
.B2(n_411),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_484),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_439),
.B(n_375),
.C(n_366),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_467),
.A2(n_461),
.B1(n_456),
.B2(n_453),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_496),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_491),
.A2(n_486),
.B1(n_476),
.B2(n_455),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_481),
.A2(n_456),
.B(n_444),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_492),
.B(n_499),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_495),
.B(n_468),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_467),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_440),
.C(n_446),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_497),
.B(n_499),
.C(n_501),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_498),
.A2(n_474),
.B1(n_484),
.B2(n_472),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_452),
.C(n_445),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_485),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_469),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_479),
.B(n_445),
.C(n_442),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_454),
.C(n_457),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_502),
.B(n_503),
.C(n_485),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_478),
.B(n_464),
.C(n_462),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_505),
.B(n_506),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_498),
.A2(n_472),
.B(n_486),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_510),
.Y(n_519)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_509),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_494),
.A2(n_486),
.B(n_476),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_511),
.B(n_512),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_466),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_513),
.A2(n_496),
.B1(n_488),
.B2(n_487),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_501),
.A2(n_468),
.B1(n_473),
.B2(n_465),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_514),
.A2(n_5),
.B1(n_15),
.B2(n_16),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_517),
.C(n_5),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_497),
.B(n_473),
.C(n_363),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_516),
.B(n_495),
.C(n_493),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_502),
.A2(n_342),
.B(n_4),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_520),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_515),
.B(n_487),
.C(n_489),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_521),
.B(n_524),
.C(n_504),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_506),
.B(n_489),
.C(n_488),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_525),
.B(n_514),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_527),
.B(n_507),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_529),
.B(n_518),
.C(n_523),
.Y(n_536)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_522),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_530),
.B(n_531),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_504),
.C(n_509),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_532),
.B(n_533),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_536),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_529),
.B(n_526),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_537),
.A2(n_524),
.B1(n_535),
.B2(n_528),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_538),
.B(n_523),
.Y(n_540)
);

A2O1A1O1Ixp25_ASAP7_75t_L g542 ( 
.A1(n_540),
.A2(n_541),
.B(n_507),
.C(n_508),
.D(n_510),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_539),
.A2(n_534),
.B(n_538),
.Y(n_541)
);

AOI322xp5_ASAP7_75t_L g543 ( 
.A1(n_542),
.A2(n_519),
.A3(n_517),
.B1(n_511),
.B2(n_516),
.C1(n_513),
.C2(n_505),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_543),
.A2(n_15),
.B(n_16),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_544),
.A2(n_15),
.B(n_18),
.Y(n_545)
);

AO21x1_ASAP7_75t_L g546 ( 
.A1(n_545),
.A2(n_18),
.B(n_1),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_18),
.Y(n_547)
);


endmodule