module fake_jpeg_15404_n_155 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_155);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_15),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_35),
.B1(n_28),
.B2(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_24),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_14),
.B1(n_17),
.B2(n_25),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_17),
.B1(n_14),
.B2(n_25),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_56),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_53),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_54),
.B(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_19),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_35),
.B1(n_36),
.B2(n_33),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_28),
.B1(n_43),
.B2(n_27),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_43),
.B1(n_37),
.B2(n_31),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_22),
.B(n_16),
.C(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_23),
.B(n_16),
.C(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx2_ASAP7_75t_SL g81 ( 
.A(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_78),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_44),
.B1(n_16),
.B2(n_26),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_75),
.B1(n_82),
.B2(n_84),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_22),
.B1(n_20),
.B2(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_48),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_59),
.B1(n_62),
.B2(n_53),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_26),
.B1(n_14),
.B2(n_25),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_57),
.A2(n_28),
.B1(n_31),
.B2(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_58),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g115 ( 
.A(n_92),
.B(n_93),
.C(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_53),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_100),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_55),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_18),
.C(n_1),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_86),
.B1(n_71),
.B2(n_73),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_59),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_85),
.B(n_68),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_103),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_27),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_13),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_104),
.Y(n_106)
);

AOI322xp5_ASAP7_75t_SL g105 ( 
.A1(n_99),
.A2(n_86),
.A3(n_74),
.B1(n_80),
.B2(n_81),
.C1(n_72),
.C2(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_114),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_77),
.B(n_84),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_110),
.Y(n_119)
);

AOI221xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_88),
.B1(n_27),
.B2(n_18),
.C(n_15),
.Y(n_111)
);

AOI322xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_113),
.A3(n_118),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_123)
);

AOI221xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_95),
.B1(n_94),
.B2(n_98),
.C(n_97),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_18),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_117),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_93),
.B1(n_98),
.B2(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_128),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_127),
.A3(n_115),
.B1(n_121),
.B2(n_7),
.C1(n_8),
.C2(n_5),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_110),
.Y(n_128)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_120),
.B(n_107),
.CI(n_116),
.CON(n_129),
.SN(n_129)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_130),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_106),
.Y(n_130)
);

OAI322xp33_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_115),
.A3(n_106),
.B1(n_118),
.B2(n_114),
.C1(n_108),
.C2(n_11),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_133),
.B(n_127),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_124),
.B(n_126),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_139),
.B1(n_132),
.B2(n_136),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_134),
.A2(n_124),
.B(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_140),
.Y(n_143)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_10),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_6),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_147),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_129),
.Y(n_145)
);

NAND2x1p5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_130),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_146),
.A2(n_129),
.B1(n_7),
.B2(n_8),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_136),
.B(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_150),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_143),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_151),
.Y(n_153)
);

AOI21x1_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_152),
.B(n_145),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_148),
.Y(n_155)
);


endmodule