module fake_jpeg_6414_n_251 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_20),
.B(n_12),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_16),
.B1(n_15),
.B2(n_25),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_13),
.B1(n_19),
.B2(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_25),
.B1(n_15),
.B2(n_18),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_19),
.B1(n_22),
.B2(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_16),
.B1(n_26),
.B2(n_13),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_51),
.B1(n_58),
.B2(n_59),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_35),
.B1(n_28),
.B2(n_37),
.Y(n_71)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_30),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_61),
.Y(n_70)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_31),
.B1(n_32),
.B2(n_40),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_71),
.B1(n_77),
.B2(n_80),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_65),
.B(n_47),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_39),
.C(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_73),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_39),
.C(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_45),
.B1(n_36),
.B2(n_43),
.Y(n_80)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_82),
.Y(n_101)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_84),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_87),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_89),
.B(n_96),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_59),
.B1(n_58),
.B2(n_49),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_91),
.B1(n_95),
.B2(n_66),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_48),
.B1(n_50),
.B2(n_45),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_63),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_73),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_61),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_55),
.B1(n_43),
.B2(n_62),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_97),
.A2(n_55),
.B1(n_69),
.B2(n_79),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_64),
.B(n_78),
.C(n_76),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_90),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_73),
.B(n_76),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_108),
.B(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_17),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_92),
.B(n_95),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_79),
.B1(n_71),
.B2(n_64),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_56),
.B1(n_82),
.B2(n_72),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_70),
.C(n_43),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_115),
.C(n_116),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_17),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_61),
.C(n_67),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_119),
.B(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_81),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_97),
.B1(n_84),
.B2(n_83),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_134),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_126),
.B(n_114),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_125),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_112),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_96),
.B(n_87),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_133),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_81),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_116),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_132),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_17),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_82),
.B1(n_86),
.B2(n_27),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_103),
.B1(n_100),
.B2(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_152),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_114),
.B1(n_107),
.B2(n_109),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_144),
.B1(n_14),
.B2(n_18),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_148),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_115),
.C(n_104),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_128),
.C(n_132),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_104),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_127),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_136),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_151),
.B(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_117),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_104),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_155),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_122),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_23),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_15),
.B1(n_25),
.B2(n_14),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_158),
.A2(n_13),
.B1(n_14),
.B2(n_23),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_130),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_162),
.B1(n_153),
.B2(n_138),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_172),
.C(n_175),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_163),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_106),
.B1(n_22),
.B2(n_19),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_146),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_176),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_106),
.C(n_88),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_17),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_141),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_88),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_177),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_156),
.B1(n_144),
.B2(n_137),
.Y(n_178)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_113),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_SL g195 ( 
.A(n_182),
.B(n_188),
.C(n_191),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_168),
.B1(n_164),
.B2(n_145),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_185),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_142),
.C(n_143),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_190),
.C(n_23),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_141),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_152),
.C(n_157),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_138),
.Y(n_192)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_158),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g207 ( 
.A(n_193),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_167),
.A2(n_88),
.B1(n_113),
.B2(n_23),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_170),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_204),
.Y(n_209)
);

OAI322xp33_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_159),
.A3(n_177),
.B1(n_172),
.B2(n_10),
.C1(n_11),
.C2(n_9),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_203),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_183),
.C(n_187),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_185),
.A2(n_11),
.B(n_9),
.C(n_2),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_201),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_23),
.B(n_21),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_0),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_206),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_208),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_211),
.A2(n_214),
.B(n_216),
.Y(n_224)
);

OAI321xp33_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_181),
.A3(n_193),
.B1(n_189),
.B2(n_180),
.C(n_182),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_188),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_183),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_113),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_201),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_218),
.A2(n_4),
.B(n_5),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_1),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_21),
.B1(n_29),
.B2(n_27),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_34),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_225),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_207),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_195),
.B(n_3),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_226),
.A2(n_230),
.B(n_4),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_34),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_229),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_228),
.B(n_222),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_233),
.B(n_5),
.Y(n_241)
);

INVx11_ASAP7_75t_L g232 ( 
.A(n_221),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_237),
.Y(n_239)
);

OAI21x1_ASAP7_75t_SL g233 ( 
.A1(n_226),
.A2(n_220),
.B(n_210),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_228),
.A2(n_213),
.B1(n_219),
.B2(n_21),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_34),
.C(n_29),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_234),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_241),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_243),
.C(n_244),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_235),
.A2(n_29),
.B(n_27),
.Y(n_244)
);

AOI321xp33_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_238),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C(n_5),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_248)
);

AOI321xp33_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_249),
.A3(n_246),
.B1(n_8),
.B2(n_7),
.C(n_21),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_247),
.B(n_7),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_8),
.Y(n_251)
);


endmodule