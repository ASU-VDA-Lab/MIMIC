module fake_jpeg_3115_n_616 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_616);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_616;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_32),
.A2(n_49),
.B1(n_36),
.B2(n_25),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_63),
.A2(n_55),
.B1(n_30),
.B2(n_20),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_72),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_22),
.B(n_9),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_81),
.Y(n_118)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_76),
.Y(n_169)
);

BUFx24_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_77),
.Y(n_164)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_80),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_22),
.B(n_9),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_82),
.Y(n_177)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_49),
.Y(n_85)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_31),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_111),
.Y(n_116)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_94),
.Y(n_176)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_96),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_106),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_39),
.B(n_9),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_108),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_31),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_107),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_34),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_109),
.B(n_110),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_35),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_29),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_121),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_46),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_125),
.B(n_173),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_41),
.B1(n_40),
.B2(n_52),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_126),
.B(n_150),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_63),
.A2(n_48),
.B1(n_40),
.B2(n_52),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_127),
.A2(n_139),
.B1(n_145),
.B2(n_161),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_24),
.B1(n_53),
.B2(n_20),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_132),
.A2(n_166),
.B1(n_77),
.B2(n_107),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_61),
.A2(n_24),
.B1(n_44),
.B2(n_43),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_58),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_82),
.B1(n_80),
.B2(n_72),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_85),
.A2(n_24),
.B1(n_44),
.B2(n_43),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_111),
.B(n_79),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_94),
.A2(n_45),
.B1(n_39),
.B2(n_51),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_151),
.Y(n_195)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_55),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_154),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_103),
.B1(n_90),
.B2(n_30),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_76),
.A2(n_48),
.B1(n_45),
.B2(n_51),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_62),
.A2(n_53),
.B1(n_20),
.B2(n_26),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_69),
.A2(n_44),
.B1(n_26),
.B2(n_43),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_172),
.A2(n_55),
.B1(n_30),
.B2(n_28),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_77),
.B(n_26),
.Y(n_173)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_178),
.Y(n_267)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_179),
.Y(n_276)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_181),
.Y(n_273)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_182),
.Y(n_266)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_183),
.Y(n_245)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_184),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_108),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_185),
.B(n_198),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_186),
.A2(n_205),
.B1(n_208),
.B2(n_212),
.Y(n_256)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_187),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_116),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g263 ( 
.A(n_189),
.B(n_210),
.C(n_225),
.Y(n_263)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_190),
.Y(n_252)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_191),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_192),
.A2(n_139),
.B1(n_126),
.B2(n_166),
.Y(n_244)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_193),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_118),
.B(n_89),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_194),
.B(n_203),
.Y(n_281)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_197),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_110),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_199),
.Y(n_282)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_137),
.Y(n_200)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_200),
.Y(n_286)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_201),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_123),
.B(n_67),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_141),
.A2(n_50),
.B1(n_42),
.B2(n_46),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_207),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_164),
.A2(n_28),
.B1(n_50),
.B2(n_42),
.Y(n_208)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_124),
.Y(n_209)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_209),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_122),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_146),
.B(n_117),
.C(n_143),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_211),
.B(n_226),
.C(n_229),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_157),
.A2(n_28),
.B1(n_156),
.B2(n_144),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_213),
.Y(n_275)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_137),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_215),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_173),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_217),
.A2(n_227),
.B1(n_155),
.B2(n_104),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_140),
.B(n_109),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_218),
.B(n_223),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_168),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_219),
.B(n_231),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_220),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_172),
.A2(n_84),
.B1(n_102),
.B2(n_96),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_221),
.A2(n_78),
.B1(n_68),
.B2(n_175),
.Y(n_284)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_135),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_222),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_150),
.B(n_86),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_133),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_228),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_150),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_119),
.B(n_98),
.C(n_97),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_157),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_136),
.B(n_74),
.C(n_70),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_115),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_230),
.Y(n_285)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_167),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_130),
.B(n_92),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_232),
.B(n_113),
.Y(n_283)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_237),
.Y(n_255)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_147),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_236),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_151),
.B(n_0),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_235),
.B(n_240),
.Y(n_246)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_148),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_129),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_160),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_145),
.B(n_0),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_130),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_241),
.B(n_181),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_244),
.A2(n_182),
.B1(n_165),
.B2(n_226),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_207),
.A2(n_134),
.B1(n_147),
.B2(n_174),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_249),
.A2(n_258),
.B1(n_259),
.B2(n_278),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_185),
.B(n_153),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_251),
.B(n_257),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_196),
.A2(n_171),
.B(n_156),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_253),
.A2(n_229),
.B(n_193),
.Y(n_310)
);

AO21x2_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_177),
.B(n_175),
.Y(n_254)
);

AO21x2_ASAP7_75t_L g306 ( 
.A1(n_254),
.A2(n_238),
.B(n_237),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_204),
.B(n_131),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_195),
.A2(n_174),
.B1(n_159),
.B2(n_163),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_SL g261 ( 
.A(n_199),
.B(n_131),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_261),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_202),
.A2(n_169),
.B1(n_158),
.B2(n_163),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_265),
.A2(n_270),
.B1(n_254),
.B2(n_259),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_235),
.A2(n_113),
.B1(n_135),
.B2(n_158),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_230),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_271),
.B(n_283),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_201),
.A2(n_159),
.B1(n_169),
.B2(n_93),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_284),
.A2(n_288),
.B1(n_219),
.B2(n_241),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_216),
.B(n_88),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_287),
.B(n_291),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_196),
.A2(n_177),
.B1(n_73),
.B2(n_165),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_216),
.B(n_71),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_209),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_222),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_188),
.B(n_73),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_295),
.B(n_220),
.Y(n_327)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_298),
.Y(n_361)
);

AO22x1_ASAP7_75t_L g299 ( 
.A1(n_244),
.A2(n_227),
.B1(n_196),
.B2(n_198),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_299),
.B(n_301),
.Y(n_393)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_243),
.Y(n_300)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_300),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_223),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_273),
.Y(n_302)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_263),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g394 ( 
.A(n_305),
.Y(n_394)
);

AO21x2_ASAP7_75t_L g358 ( 
.A1(n_306),
.A2(n_314),
.B(n_331),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_218),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_307),
.B(n_312),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_253),
.A2(n_228),
.B1(n_180),
.B2(n_234),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_309),
.A2(n_333),
.B1(n_336),
.B2(n_258),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_310),
.A2(n_315),
.B(n_320),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_211),
.Y(n_312)
);

OAI32xp33_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_191),
.A3(n_183),
.B1(n_231),
.B2(n_184),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_329),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_239),
.C(n_233),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_316),
.B(n_318),
.C(n_262),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_246),
.A2(n_190),
.B1(n_197),
.B2(n_224),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_317),
.A2(n_332),
.B1(n_260),
.B2(n_255),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_272),
.B(n_214),
.C(n_200),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_319),
.A2(n_345),
.B1(n_294),
.B2(n_252),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_246),
.A2(n_219),
.B(n_187),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_281),
.B(n_206),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_321),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_254),
.Y(n_322)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_322),
.Y(n_366)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_282),
.B(n_178),
.CI(n_112),
.CON(n_324),
.SN(n_324)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_324),
.B(n_339),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_325),
.B(n_327),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_254),
.A2(n_181),
.B(n_179),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_326),
.A2(n_278),
.B(n_267),
.Y(n_349)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_243),
.Y(n_328)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_328),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_0),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_245),
.Y(n_330)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

O2A1O1Ixp33_ASAP7_75t_SL g331 ( 
.A1(n_254),
.A2(n_293),
.B(n_256),
.C(n_282),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_293),
.A2(n_265),
.B1(n_251),
.B2(n_289),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_254),
.A2(n_289),
.B1(n_257),
.B2(n_242),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_274),
.B(n_0),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_334),
.B(n_343),
.Y(n_386)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_245),
.Y(n_335)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_242),
.A2(n_120),
.B1(n_181),
.B2(n_35),
.Y(n_336)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_338),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_11),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_269),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_340),
.B(n_341),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_269),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_273),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_342),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_274),
.B(n_1),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_287),
.B(n_11),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_344),
.B(n_347),
.Y(n_372)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_250),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_291),
.B(n_35),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_346),
.B(n_269),
.Y(n_378)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_260),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_SL g348 ( 
.A(n_288),
.B(n_10),
.C(n_18),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g368 ( 
.A(n_348),
.B(n_267),
.CI(n_14),
.CON(n_368),
.SN(n_368)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_349),
.A2(n_357),
.B(n_365),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_354),
.C(n_374),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_332),
.A2(n_262),
.B1(n_255),
.B2(n_292),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_351),
.A2(n_360),
.B1(n_379),
.B2(n_389),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_373),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_275),
.C(n_264),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_311),
.A2(n_283),
.B(n_255),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_359),
.A2(n_370),
.B1(n_381),
.B2(n_385),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_310),
.A2(n_248),
.B1(n_247),
.B2(n_249),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_311),
.A2(n_267),
.B(n_271),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_SL g401 ( 
.A(n_368),
.B(n_383),
.C(n_301),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_299),
.A2(n_248),
.B1(n_247),
.B2(n_294),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_324),
.B(n_269),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_275),
.C(n_264),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_378),
.B(n_313),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_312),
.A2(n_307),
.B1(n_322),
.B2(n_299),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_337),
.A2(n_297),
.B(n_266),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_382),
.Y(n_400)
);

A2O1A1O1Ixp25_ASAP7_75t_L g383 ( 
.A1(n_301),
.A2(n_279),
.B(n_252),
.C(n_286),
.D(n_266),
.Y(n_383)
);

OAI31xp33_ASAP7_75t_SL g384 ( 
.A1(n_320),
.A2(n_279),
.A3(n_285),
.B(n_250),
.Y(n_384)
);

OA21x2_ASAP7_75t_L g422 ( 
.A1(n_384),
.A2(n_336),
.B(n_328),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_322),
.A2(n_290),
.B1(n_250),
.B2(n_276),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_327),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_387),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_334),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_388),
.B(n_391),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_308),
.A2(n_290),
.B1(n_286),
.B2(n_268),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_308),
.A2(n_268),
.B1(n_276),
.B2(n_285),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_390),
.A2(n_342),
.B1(n_302),
.B2(n_1),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_343),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_304),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_396),
.B(n_423),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_367),
.B(n_323),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_397),
.Y(n_462)
);

FAx1_ASAP7_75t_SL g399 ( 
.A(n_379),
.B(n_333),
.CI(n_309),
.CON(n_399),
.SN(n_399)
);

XOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_399),
.B(n_355),
.Y(n_464)
);

OR2x6_ASAP7_75t_L g446 ( 
.A(n_401),
.B(n_412),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_403),
.B(n_351),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_372),
.B(n_323),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_404),
.B(n_416),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_371),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_405),
.B(n_413),
.Y(n_448)
);

OAI21xp33_ASAP7_75t_L g407 ( 
.A1(n_394),
.A2(n_325),
.B(n_303),
.Y(n_407)
);

BUFx5_ASAP7_75t_L g465 ( 
.A(n_407),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_364),
.A2(n_306),
.B1(n_319),
.B2(n_326),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_408),
.A2(n_422),
.B1(n_429),
.B2(n_366),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_358),
.A2(n_306),
.B1(n_331),
.B2(n_341),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_409),
.A2(n_411),
.B1(n_415),
.B2(n_418),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_358),
.A2(n_306),
.B1(n_331),
.B2(n_340),
.Y(n_411)
);

XOR2x2_ASAP7_75t_L g412 ( 
.A(n_356),
.B(n_329),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_371),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_358),
.A2(n_306),
.B1(n_314),
.B2(n_303),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_356),
.B(n_300),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_362),
.Y(n_417)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_417),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_358),
.A2(n_324),
.B1(n_317),
.B2(n_347),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_372),
.B(n_335),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_419),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_374),
.B(n_346),
.C(n_330),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_430),
.C(n_433),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_361),
.B(n_345),
.Y(n_421)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_421),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_354),
.B(n_348),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_365),
.Y(n_424)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_424),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_361),
.B(n_338),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_425),
.Y(n_441)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_362),
.Y(n_427)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_427),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_385),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_428),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_378),
.B(n_342),
.C(n_3),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_364),
.B(n_393),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_433),
.Y(n_459)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_376),
.Y(n_432)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_432),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_393),
.B(n_19),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_434),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_406),
.A2(n_358),
.B1(n_373),
.B2(n_393),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_437),
.A2(n_451),
.B1(n_458),
.B2(n_463),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_439),
.B(n_427),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_395),
.B(n_353),
.C(n_369),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_444),
.C(n_453),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_417),
.Y(n_443)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_443),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_395),
.B(n_353),
.C(n_369),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_445),
.B(n_423),
.Y(n_479)
);

AO22x1_ASAP7_75t_L g449 ( 
.A1(n_418),
.A2(n_360),
.B1(n_366),
.B2(n_352),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_449),
.B(n_399),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_406),
.A2(n_358),
.B1(n_373),
.B2(n_359),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_400),
.A2(n_355),
.B1(n_387),
.B2(n_388),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_452),
.A2(n_454),
.B1(n_466),
.B2(n_467),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_396),
.B(n_357),
.C(n_391),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_402),
.A2(n_370),
.B1(n_349),
.B2(n_384),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_420),
.B(n_382),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_403),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_402),
.A2(n_413),
.B1(n_405),
.B2(n_400),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_431),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_410),
.A2(n_380),
.B1(n_392),
.B2(n_386),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_428),
.A2(n_380),
.B1(n_392),
.B2(n_386),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_426),
.A2(n_383),
.B(n_390),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_468),
.A2(n_422),
.B(n_383),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_415),
.A2(n_389),
.B1(n_375),
.B2(n_363),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_470),
.A2(n_435),
.B1(n_461),
.B2(n_468),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_414),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_471),
.B(n_434),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_473),
.B(n_477),
.Y(n_515)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_474),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_476),
.A2(n_498),
.B1(n_449),
.B2(n_495),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_412),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_478),
.B(n_480),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_479),
.B(n_446),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_363),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_426),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_481),
.B(n_486),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_430),
.C(n_424),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_485),
.C(n_488),
.Y(n_504)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_448),
.Y(n_483)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_483),
.Y(n_516)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_443),
.Y(n_484)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_484),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_444),
.B(n_447),
.C(n_439),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_453),
.B(n_447),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_443),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_487),
.B(n_489),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_445),
.B(n_401),
.C(n_432),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_436),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_462),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_490),
.B(n_496),
.Y(n_525)
);

CKINVDCx14_ASAP7_75t_R g517 ( 
.A(n_491),
.Y(n_517)
);

AOI21x1_ASAP7_75t_L g492 ( 
.A1(n_450),
.A2(n_398),
.B(n_465),
.Y(n_492)
);

OAI21x1_ASAP7_75t_SL g513 ( 
.A1(n_492),
.A2(n_494),
.B(n_495),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_463),
.A2(n_411),
.B(n_409),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_436),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_497),
.B(n_503),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_435),
.A2(n_399),
.B1(n_422),
.B2(n_429),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_456),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_499),
.A2(n_500),
.B1(n_469),
.B2(n_438),
.Y(n_521)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_456),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_501),
.A2(n_446),
.B1(n_465),
.B2(n_368),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_459),
.B(n_375),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_505),
.A2(n_8),
.B1(n_17),
.B2(n_4),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_459),
.C(n_464),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_507),
.B(n_519),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_486),
.B(n_497),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_511),
.B(n_514),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_493),
.A2(n_457),
.B1(n_452),
.B2(n_470),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_512),
.B(n_531),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_481),
.B(n_458),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_475),
.B(n_440),
.C(n_437),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_SL g520 ( 
.A(n_477),
.B(n_446),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_520),
.B(n_5),
.Y(n_553)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_521),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_522),
.B(n_524),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_472),
.A2(n_451),
.B1(n_449),
.B2(n_469),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_523),
.A2(n_531),
.B1(n_8),
.B2(n_16),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_503),
.B(n_446),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_475),
.B(n_377),
.Y(n_526)
);

CKINVDCx14_ASAP7_75t_R g540 ( 
.A(n_526),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_528),
.A2(n_474),
.B1(n_476),
.B2(n_494),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_488),
.B(n_446),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_529),
.B(n_530),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_482),
.B(n_368),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_498),
.A2(n_377),
.B1(n_368),
.B2(n_4),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_535),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_511),
.B(n_479),
.C(n_484),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_536),
.B(n_538),
.Y(n_560)
);

OAI221xp5_ASAP7_75t_L g539 ( 
.A1(n_506),
.A2(n_501),
.B1(n_493),
.B2(n_487),
.C(n_502),
.Y(n_539)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_539),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_519),
.B(n_504),
.C(n_527),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_541),
.B(n_543),
.Y(n_564)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_525),
.Y(n_542)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_542),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_517),
.B(n_500),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_529),
.A2(n_492),
.B(n_502),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_544),
.A2(n_510),
.B1(n_523),
.B2(n_509),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_516),
.B(n_499),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_545),
.A2(n_7),
.B(n_10),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_504),
.B(n_1),
.C(n_3),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_546),
.B(n_551),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_SL g554 ( 
.A1(n_547),
.A2(n_549),
.B1(n_528),
.B2(n_518),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_527),
.B(n_10),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_550),
.B(n_5),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_508),
.B(n_1),
.C(n_3),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_508),
.B(n_5),
.C(n_6),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_552),
.B(n_507),
.C(n_522),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_553),
.A2(n_513),
.B1(n_530),
.B2(n_524),
.Y(n_557)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_554),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_556),
.B(n_570),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_557),
.B(n_572),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_558),
.B(n_559),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_541),
.B(n_514),
.C(n_505),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_545),
.B(n_520),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_561),
.B(n_563),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_SL g563 ( 
.A(n_537),
.B(n_515),
.C(n_6),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_548),
.B(n_515),
.C(n_7),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_565),
.B(n_550),
.C(n_546),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_566),
.B(n_568),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_567),
.A2(n_547),
.B(n_534),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_540),
.B(n_7),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_533),
.B(n_19),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_535),
.Y(n_572)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_573),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_564),
.B(n_536),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_574),
.B(n_580),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_555),
.A2(n_537),
.B(n_532),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_576),
.B(n_581),
.Y(n_595)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_579),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_559),
.B(n_532),
.C(n_534),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g581 ( 
.A1(n_561),
.A2(n_552),
.B(n_551),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_560),
.B(n_562),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_582),
.B(n_583),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_572),
.B(n_10),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_571),
.B(n_11),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_586),
.B(n_588),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_558),
.B(n_11),
.C(n_15),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_577),
.B(n_580),
.C(n_578),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_589),
.B(n_593),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_585),
.A2(n_571),
.B1(n_570),
.B2(n_557),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_587),
.B(n_565),
.C(n_563),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_594),
.B(n_596),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_587),
.B(n_584),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_584),
.B(n_567),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_599),
.A2(n_581),
.B(n_579),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_590),
.Y(n_600)
);

AO21x1_ASAP7_75t_L g610 ( 
.A1(n_600),
.A2(n_603),
.B(n_606),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_592),
.B(n_575),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_601),
.B(n_604),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_595),
.B(n_596),
.C(n_598),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_597),
.B(n_588),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_605),
.B(n_591),
.Y(n_609)
);

A2O1A1Ixp33_ASAP7_75t_L g607 ( 
.A1(n_602),
.A2(n_599),
.B(n_591),
.C(n_573),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_607),
.B(n_609),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_SL g612 ( 
.A1(n_610),
.A2(n_569),
.B(n_16),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_612),
.B(n_15),
.Y(n_613)
);

OAI211xp5_ASAP7_75t_L g614 ( 
.A1(n_613),
.A2(n_608),
.B(n_611),
.C(n_19),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_614),
.A2(n_15),
.B(n_16),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_615),
.B(n_15),
.Y(n_616)
);


endmodule