module fake_jpeg_1430_n_195 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_195);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_20),
.B(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_19),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_1),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_63),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_75),
.A2(n_64),
.B1(n_53),
.B2(n_61),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_83),
.B1(n_58),
.B2(n_68),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_64),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_81),
.B(n_55),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_64),
.B1(n_61),
.B2(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_88),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_89),
.B(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_89),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_107),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_72),
.B1(n_69),
.B2(n_60),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_101),
.B1(n_63),
.B2(n_80),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_102),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_68),
.B1(n_77),
.B2(n_67),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_58),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_67),
.B(n_54),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_51),
.Y(n_110)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_108),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_57),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_2),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_126),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_80),
.B1(n_90),
.B2(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_117),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_102),
.B1(n_95),
.B2(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_1),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_3),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_125),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_55),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

AO22x1_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_3),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_4),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_5),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_49),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_23),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_6),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_133),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_147),
.B1(n_149),
.B2(n_124),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_105),
.B1(n_99),
.B2(n_108),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_131),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_163)
);

AOI21x1_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_102),
.B(n_96),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_136),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_22),
.C(n_46),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_137),
.C(n_40),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_140),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_115),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_21),
.C(n_42),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_128),
.Y(n_141)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_27),
.B(n_39),
.C(n_36),
.D(n_35),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_143),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_7),
.B(n_9),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_152),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_157),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_163),
.B1(n_148),
.B2(n_165),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_160),
.A2(n_165),
.B(n_129),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_134),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_31),
.C(n_29),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_149),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_144),
.A2(n_26),
.B1(n_12),
.B2(n_13),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_11),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_137),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_170),
.B1(n_173),
.B2(n_176),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_139),
.B1(n_155),
.B2(n_164),
.Y(n_180)
);

INVxp33_ASAP7_75t_SL g170 ( 
.A(n_154),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_160),
.B(n_159),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_155),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_146),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_181),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_156),
.B1(n_147),
.B2(n_161),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_179),
.A2(n_183),
.B1(n_175),
.B2(n_172),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_182),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_162),
.B(n_13),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_185),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_181),
.B(n_174),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_182),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_191),
.B1(n_186),
.B2(n_184),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_192),
.Y(n_193)
);

AOI221xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_189),
.B1(n_190),
.B2(n_18),
.C(n_16),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_17),
.Y(n_195)
);


endmodule