module fake_ariane_1297_n_1180 (n_295, n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_289, n_288, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_294, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_269, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_274, n_115, n_272, n_133, n_66, n_205, n_236, n_265, n_71, n_267, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_281, n_209, n_49, n_262, n_291, n_20, n_292, n_174, n_275, n_100, n_17, n_283, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_297, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_271, n_46, n_290, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_286, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_287, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_284, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_278, n_122, n_268, n_257, n_266, n_198, n_282, n_148, n_232, n_164, n_52, n_277, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_293, n_171, n_228, n_15, n_118, n_93, n_121, n_276, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_279, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_270, n_194, n_97, n_154, n_280, n_215, n_252, n_142, n_251, n_161, n_285, n_14, n_163, n_88, n_186, n_141, n_296, n_298, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_273, n_54, n_25, n_1180);

input n_295;
input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_289;
input n_288;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_294;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_269;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_274;
input n_115;
input n_272;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_267;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_281;
input n_209;
input n_49;
input n_262;
input n_291;
input n_20;
input n_292;
input n_174;
input n_275;
input n_100;
input n_17;
input n_283;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_297;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_271;
input n_46;
input n_290;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_286;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_287;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_284;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_278;
input n_122;
input n_268;
input n_257;
input n_266;
input n_198;
input n_282;
input n_148;
input n_232;
input n_164;
input n_52;
input n_277;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_293;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_276;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_279;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_270;
input n_194;
input n_97;
input n_154;
input n_280;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_285;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_296;
input n_298;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_273;
input n_54;
input n_25;

output n_1180;

wire n_356;
wire n_556;
wire n_1127;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_1020;
wire n_1137;
wire n_646;
wire n_1174;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_423;
wire n_347;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_479;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_690;
wire n_416;
wire n_969;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_679;
wire n_643;
wire n_924;
wire n_927;
wire n_781;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_586;
wire n_952;
wire n_864;
wire n_443;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_1154;
wire n_1166;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_1138;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_670;
wire n_607;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_1131;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1167;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_945;
wire n_702;
wire n_905;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_779;
wire n_336;
wire n_731;
wire n_754;
wire n_903;
wire n_871;
wire n_315;
wire n_1073;
wire n_594;
wire n_1173;
wire n_311;
wire n_402;
wire n_1052;
wire n_1068;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_553;
wire n_446;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_557;
wire n_405;
wire n_1107;
wire n_858;
wire n_645;
wire n_989;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_1134;
wire n_485;
wire n_401;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_822;
wire n_1143;
wire n_344;
wire n_795;
wire n_381;
wire n_721;
wire n_433;
wire n_481;
wire n_600;
wire n_840;
wire n_426;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_561;
wire n_770;
wire n_821;
wire n_928;
wire n_839;
wire n_1099;
wire n_1153;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_369;
wire n_894;
wire n_787;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_604;
wire n_677;
wire n_614;
wire n_439;
wire n_1172;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_1160;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_689;
wire n_694;
wire n_400;
wire n_884;
wire n_1116;
wire n_983;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1085;
wire n_467;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_1080;
wire n_576;
wire n_843;
wire n_1148;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_728;
wire n_388;
wire n_449;
wire n_333;
wire n_612;
wire n_957;
wire n_392;
wire n_376;
wire n_413;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_685;
wire n_459;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_1142;
wire n_617;
wire n_616;
wire n_705;
wire n_630;
wire n_658;
wire n_1140;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_1089;
wire n_565;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_1135;
wire n_918;
wire n_639;
wire n_673;
wire n_452;
wire n_1114;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_571;
wire n_680;
wire n_414;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_534;
wire n_1108;
wire n_355;
wire n_609;
wire n_851;
wire n_444;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_947;
wire n_409;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_774;
wire n_872;
wire n_933;
wire n_407;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_1157;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_982;
wire n_915;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_1178;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_666;
wire n_306;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_622;
wire n_697;
wire n_998;
wire n_967;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_746;
wire n_456;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_751;
wire n_1027;
wire n_615;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_1139;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_580;
wire n_358;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1129;
wire n_1102;
wire n_563;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_972;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_782;
wire n_856;
wire n_1161;
wire n_425;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_1164;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_23),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_238),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_17),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_29),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_80),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_191),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_89),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_68),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_20),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_142),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_163),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_130),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_216),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_176),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_217),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_124),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_297),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_40),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_256),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_140),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_283),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_31),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_278),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_8),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_245),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_188),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_147),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_10),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_166),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_189),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_5),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_175),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_22),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_90),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_87),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_199),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_282),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_125),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_103),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_219),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_44),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_231),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_160),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_20),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_150),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_192),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_27),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_4),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_279),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_215),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_234),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_229),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_10),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_255),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_50),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_154),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_200),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_146),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_11),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_289),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_11),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_91),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_72),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_78),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_57),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_37),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_23),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_129),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_246),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_134),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_14),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_290),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_66),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_43),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_208),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_148),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_45),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_46),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_252),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_17),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_156),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_119),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_165),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_19),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_184),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_288),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_260),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_116),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_143),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_95),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_114),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_269),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_110),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_295),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_32),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_104),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_12),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_86),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_58),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_190),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_61),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_25),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_55),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_98),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_75),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_202),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_38),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_159),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_242),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_185),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_172),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_21),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_6),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_179),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_213),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_79),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_296),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_162),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_5),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_128),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_137),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_247),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_101),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_100),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_7),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_180),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_233),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_51),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_212),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_267),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_65),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_123),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_177),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_183),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_205),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_249),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_15),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_155),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_228),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_271),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_121),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_149),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_250),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_181),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_263),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_164),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_139),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_69),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_285),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_158),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_14),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_21),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_24),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_151),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_251),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_286),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_60),
.Y(n_455)
);

BUFx10_ASAP7_75t_L g456 ( 
.A(n_298),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_284),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_42),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_226),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_222),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_7),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_178),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_194),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_211),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_39),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_161),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_240),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_225),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_67),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_102),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_266),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_28),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_26),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_126),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_274),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_272),
.Y(n_476)
);

BUFx4f_ASAP7_75t_SL g477 ( 
.A(n_15),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_127),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_292),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_81),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_169),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_153),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_56),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_84),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_52),
.Y(n_485)
);

BUFx10_ASAP7_75t_L g486 ( 
.A(n_171),
.Y(n_486)
);

BUFx8_ASAP7_75t_SL g487 ( 
.A(n_281),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_112),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_141),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_97),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_111),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_76),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_182),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_77),
.Y(n_494)
);

BUFx10_ASAP7_75t_L g495 ( 
.A(n_265),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_210),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_293),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_254),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_326),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_367),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_346),
.Y(n_501)
);

NOR2xp67_ASAP7_75t_L g502 ( 
.A(n_299),
.B(n_301),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_487),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_375),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_425),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_351),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_445),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_L g508 ( 
.A(n_365),
.B(n_0),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_L g509 ( 
.A(n_369),
.B(n_0),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_L g510 ( 
.A(n_417),
.B(n_1),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_465),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_307),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_326),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_482),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_488),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_382),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_382),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g518 ( 
.A(n_423),
.B(n_1),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_410),
.B(n_327),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_331),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_449),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_357),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_329),
.B(n_2),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_451),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_378),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_461),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_435),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_450),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_300),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_304),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_395),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_308),
.Y(n_533)
);

INVxp67_ASAP7_75t_SL g534 ( 
.A(n_314),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_350),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_455),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_322),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_359),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_455),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_342),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_456),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_309),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_310),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_456),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_312),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_486),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_486),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_315),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_495),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_316),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_495),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_314),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_303),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_305),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_311),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_334),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_411),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_319),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_338),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_320),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_313),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_317),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_338),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_323),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_477),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_387),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_318),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_477),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_328),
.Y(n_569)
);

NOR2xp67_ASAP7_75t_L g570 ( 
.A(n_330),
.B(n_2),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_324),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_332),
.B(n_339),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_356),
.B(n_361),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_362),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_363),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_333),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_335),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_364),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_371),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_334),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_376),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_379),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_337),
.Y(n_583)
);

INVxp33_ASAP7_75t_SL g584 ( 
.A(n_340),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_343),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_344),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_384),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_388),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_390),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_457),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_345),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_393),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_347),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_391),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_348),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_399),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_416),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_349),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_418),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_352),
.Y(n_600)
);

INVxp67_ASAP7_75t_SL g601 ( 
.A(n_393),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_354),
.Y(n_602)
);

NOR2xp67_ASAP7_75t_L g603 ( 
.A(n_424),
.B(n_3),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_408),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_429),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_430),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_408),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_447),
.Y(n_608)
);

INVxp67_ASAP7_75t_SL g609 ( 
.A(n_447),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_433),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_437),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_355),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_504),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_552),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_505),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_556),
.B(n_440),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_507),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_521),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_556),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_511),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_523),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_526),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_580),
.B(n_458),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_514),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_520),
.B(n_453),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_580),
.B(n_460),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_SL g627 ( 
.A(n_559),
.B(n_321),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_538),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_528),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_552),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_530),
.B(n_325),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_503),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_500),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_499),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_529),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_515),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_531),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_533),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_584),
.B(n_462),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_513),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_542),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_517),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_543),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_540),
.B(n_453),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_519),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_537),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_516),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_573),
.B(n_463),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_553),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_554),
.Y(n_650)
);

NOR2xp67_ASAP7_75t_L g651 ( 
.A(n_546),
.B(n_360),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_573),
.B(n_466),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_532),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_555),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_R g655 ( 
.A(n_545),
.B(n_498),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_561),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_612),
.B(n_468),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_538),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_611),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_562),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_610),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_563),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_548),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_567),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_569),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_574),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_590),
.Y(n_667)
);

OA21x2_ASAP7_75t_L g668 ( 
.A1(n_572),
.A2(n_481),
.B(n_480),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_575),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_550),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_558),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_578),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_579),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_560),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_564),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_581),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_571),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_582),
.Y(n_678)
);

CKINVDCx16_ASAP7_75t_R g679 ( 
.A(n_590),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_587),
.B(n_491),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_588),
.Y(n_681)
);

NOR2xp67_ASAP7_75t_L g682 ( 
.A(n_547),
.B(n_438),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_506),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_534),
.B(n_492),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_589),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_594),
.B(n_493),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_596),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_576),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_597),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_577),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_599),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_583),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_566),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_605),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_606),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_585),
.B(n_341),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_586),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_591),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_593),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_604),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_613),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_619),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_625),
.B(n_595),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_614),
.Y(n_704)
);

AND2x2_ASAP7_75t_SL g705 ( 
.A(n_679),
.B(n_501),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_614),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_639),
.B(n_598),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_633),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_630),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_657),
.B(n_600),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_614),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_636),
.Y(n_712)
);

AND2x6_ASAP7_75t_L g713 ( 
.A(n_677),
.B(n_475),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_625),
.A2(n_602),
.B1(n_525),
.B2(n_527),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_634),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_660),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_625),
.B(n_601),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_660),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_700),
.B(n_536),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_640),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_693),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_660),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_649),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_632),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_668),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_692),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_642),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_644),
.B(n_646),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_650),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_637),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_655),
.B(n_638),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_645),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_618),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_621),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_641),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_643),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_622),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_663),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_672),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_625),
.B(n_609),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_665),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_670),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_683),
.B(n_557),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_665),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_629),
.Y(n_745)
);

NOR2x1p5_ASAP7_75t_L g746 ( 
.A(n_671),
.B(n_522),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_651),
.B(n_539),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_615),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_666),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_635),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_666),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_647),
.B(n_535),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_674),
.B(n_506),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_678),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_681),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_685),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_653),
.B(n_541),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_682),
.B(n_544),
.Y(n_758)
);

AND2x6_ASAP7_75t_L g759 ( 
.A(n_669),
.B(n_475),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_669),
.B(n_654),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_689),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_656),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_659),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_675),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_688),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_648),
.B(n_608),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_648),
.B(n_549),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_690),
.B(n_568),
.Y(n_768)
);

AND2x6_ASAP7_75t_L g769 ( 
.A(n_661),
.B(n_478),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_631),
.B(n_551),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_664),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_673),
.Y(n_772)
);

AND2x2_ASAP7_75t_SL g773 ( 
.A(n_652),
.B(n_592),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_676),
.B(n_592),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_687),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_696),
.B(n_607),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_668),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_684),
.B(n_512),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_697),
.Y(n_779)
);

BUFx6f_ASAP7_75t_SL g780 ( 
.A(n_667),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_691),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_652),
.B(n_607),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_698),
.B(n_502),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_710),
.B(n_699),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_707),
.B(n_694),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_728),
.B(n_617),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_720),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_767),
.A2(n_695),
.B(n_686),
.C(n_680),
.Y(n_788)
);

AND2x6_ASAP7_75t_SL g789 ( 
.A(n_753),
.B(n_524),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_721),
.B(n_620),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_727),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_743),
.B(n_624),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_732),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_724),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_733),
.Y(n_795)
);

NAND2x1p5_ASAP7_75t_L g796 ( 
.A(n_726),
.B(n_735),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_714),
.B(n_764),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_708),
.B(n_627),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_766),
.A2(n_686),
.B(n_680),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_709),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_764),
.B(n_565),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_782),
.A2(n_603),
.B1(n_570),
.B2(n_616),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_765),
.B(n_662),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_773),
.A2(n_623),
.B1(n_626),
.B2(n_616),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_765),
.B(n_565),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_744),
.B(n_623),
.Y(n_806)
);

INVx8_ASAP7_75t_L g807 ( 
.A(n_780),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_SL g808 ( 
.A1(n_705),
.A2(n_658),
.B1(n_628),
.B2(n_730),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_738),
.B(n_508),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_768),
.B(n_626),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_706),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_702),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_744),
.B(n_302),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_771),
.A2(n_763),
.B1(n_737),
.B2(n_745),
.Y(n_814)
);

OR2x6_ASAP7_75t_L g815 ( 
.A(n_742),
.B(n_509),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_SL g816 ( 
.A1(n_776),
.A2(n_478),
.B1(n_336),
.B2(n_442),
.Y(n_816)
);

BUFx5_ASAP7_75t_L g817 ( 
.A(n_725),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_703),
.A2(n_510),
.B1(n_518),
.B2(n_497),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_779),
.B(n_3),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_774),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_734),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_741),
.B(n_306),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_741),
.B(n_472),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_736),
.B(n_783),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_770),
.B(n_749),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_749),
.B(n_474),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_751),
.B(n_476),
.Y(n_827)
);

AOI22x1_ASAP7_75t_L g828 ( 
.A1(n_751),
.A2(n_762),
.B1(n_772),
.B2(n_750),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_723),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_760),
.B(n_358),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_760),
.B(n_366),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_775),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_778),
.B(n_496),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_781),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_778),
.B(n_368),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_731),
.B(n_370),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_748),
.B(n_4),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_718),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_748),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_771),
.A2(n_420),
.B1(n_392),
.B2(n_400),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_729),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_771),
.A2(n_353),
.B1(n_446),
.B2(n_484),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_757),
.A2(n_467),
.B(n_8),
.C(n_9),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_747),
.B(n_758),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_774),
.B(n_372),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_747),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_759),
.A2(n_494),
.B1(n_490),
.B2(n_489),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_713),
.B(n_373),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_739),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_756),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_725),
.A2(n_383),
.B1(n_397),
.B2(n_479),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_758),
.B(n_374),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_717),
.A2(n_6),
.B(n_9),
.C(n_12),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_754),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_754),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_715),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_712),
.B(n_13),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_754),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_755),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_701),
.B(n_746),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_759),
.A2(n_485),
.B1(n_483),
.B2(n_473),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_711),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_759),
.A2(n_471),
.B1(n_470),
.B2(n_469),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_787),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_800),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_794),
.B(n_704),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_791),
.Y(n_867)
);

AO22x1_ASAP7_75t_L g868 ( 
.A1(n_784),
.A2(n_713),
.B1(n_769),
.B2(n_719),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_839),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_793),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_786),
.B(n_719),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_795),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_821),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_832),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_829),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_849),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_846),
.B(n_704),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_785),
.B(n_713),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_834),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_825),
.B(n_810),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_799),
.B(n_740),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_813),
.B(n_706),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_812),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_804),
.B(n_755),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_856),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_807),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_841),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_820),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_807),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_850),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_R g891 ( 
.A(n_790),
.B(n_769),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_796),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_803),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_792),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_837),
.B(n_706),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_838),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_803),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_828),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_844),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_808),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_788),
.B(n_755),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_798),
.B(n_718),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_806),
.B(n_761),
.Y(n_903)
);

INVxp67_ASAP7_75t_SL g904 ( 
.A(n_817),
.Y(n_904)
);

BUFx8_ASAP7_75t_L g905 ( 
.A(n_860),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_797),
.B(n_761),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_819),
.Y(n_907)
);

BUFx12f_ASAP7_75t_L g908 ( 
.A(n_789),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_862),
.Y(n_909)
);

NOR3xp33_ASAP7_75t_SL g910 ( 
.A(n_801),
.B(n_380),
.C(n_377),
.Y(n_910)
);

NOR3xp33_ASAP7_75t_SL g911 ( 
.A(n_805),
.B(n_385),
.C(n_381),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_857),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_R g913 ( 
.A(n_838),
.B(n_769),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_811),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_833),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_847),
.B(n_718),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_809),
.Y(n_917)
);

NOR3xp33_ASAP7_75t_SL g918 ( 
.A(n_824),
.B(n_389),
.C(n_386),
.Y(n_918)
);

CKINVDCx11_ASAP7_75t_R g919 ( 
.A(n_815),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_828),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_815),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_904),
.A2(n_823),
.B(n_822),
.Y(n_922)
);

OAI21x1_ASAP7_75t_L g923 ( 
.A1(n_898),
.A2(n_777),
.B(n_854),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_892),
.B(n_809),
.Y(n_924)
);

AOI21xp33_ASAP7_75t_L g925 ( 
.A1(n_915),
.A2(n_816),
.B(n_835),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_904),
.A2(n_814),
.B1(n_827),
.B2(n_826),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_880),
.B(n_802),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_901),
.A2(n_863),
.B(n_861),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_881),
.A2(n_831),
.B(n_830),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_915),
.B(n_845),
.Y(n_930)
);

OAI21x1_ASAP7_75t_L g931 ( 
.A1(n_920),
.A2(n_777),
.B(n_855),
.Y(n_931)
);

AO31x2_ASAP7_75t_L g932 ( 
.A1(n_906),
.A2(n_859),
.A3(n_858),
.B(n_716),
.Y(n_932)
);

OA22x2_ASAP7_75t_L g933 ( 
.A1(n_894),
.A2(n_852),
.B1(n_818),
.B2(n_848),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_871),
.B(n_899),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_909),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_884),
.A2(n_722),
.B(n_851),
.Y(n_936)
);

NAND3xp33_ASAP7_75t_L g937 ( 
.A(n_878),
.B(n_843),
.C(n_836),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_903),
.A2(n_811),
.B(n_853),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_864),
.A2(n_811),
.B1(n_842),
.B2(n_840),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_867),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_890),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_882),
.A2(n_817),
.B(n_752),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_899),
.B(n_870),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_891),
.B(n_817),
.Y(n_944)
);

OAI21x1_ASAP7_75t_L g945 ( 
.A1(n_916),
.A2(n_817),
.B(n_761),
.Y(n_945)
);

OAI22x1_ASAP7_75t_L g946 ( 
.A1(n_900),
.A2(n_422),
.B1(n_464),
.B2(n_459),
.Y(n_946)
);

NOR2xp67_ASAP7_75t_SL g947 ( 
.A(n_889),
.B(n_394),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_906),
.A2(n_817),
.B(n_33),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_869),
.B(n_396),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_897),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_897),
.B(n_912),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_907),
.B(n_398),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_895),
.A2(n_34),
.B(n_30),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_912),
.B(n_13),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_866),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_872),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_896),
.A2(n_36),
.B(n_35),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_907),
.B(n_16),
.Y(n_958)
);

INVx5_ASAP7_75t_L g959 ( 
.A(n_886),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_873),
.B(n_16),
.Y(n_960)
);

AOI221x1_ASAP7_75t_L g961 ( 
.A1(n_885),
.A2(n_397),
.B1(n_383),
.B2(n_22),
.C(n_24),
.Y(n_961)
);

AO21x1_ASAP7_75t_L g962 ( 
.A1(n_902),
.A2(n_397),
.B(n_383),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_874),
.A2(n_402),
.B(n_401),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_886),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_868),
.A2(n_404),
.B(n_403),
.Y(n_965)
);

AO21x2_ASAP7_75t_L g966 ( 
.A1(n_923),
.A2(n_931),
.B(n_936),
.Y(n_966)
);

INVxp67_ASAP7_75t_SL g967 ( 
.A(n_943),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_940),
.Y(n_968)
);

INVx6_ASAP7_75t_L g969 ( 
.A(n_959),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_956),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_929),
.A2(n_879),
.B(n_887),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_948),
.A2(n_875),
.B(n_865),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_941),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_955),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_945),
.A2(n_957),
.B(n_938),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_935),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_953),
.A2(n_883),
.B(n_876),
.Y(n_977)
);

OAI222xp33_ASAP7_75t_L g978 ( 
.A1(n_933),
.A2(n_921),
.B1(n_917),
.B2(n_893),
.C1(n_888),
.C2(n_877),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_922),
.A2(n_914),
.B(n_888),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_932),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_942),
.A2(n_914),
.B(n_913),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_962),
.A2(n_918),
.B(n_911),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_951),
.B(n_866),
.Y(n_983)
);

OA21x2_ASAP7_75t_L g984 ( 
.A1(n_961),
.A2(n_911),
.B(n_910),
.Y(n_984)
);

NOR2xp67_ASAP7_75t_L g985 ( 
.A(n_959),
.B(n_908),
.Y(n_985)
);

BUFx2_ASAP7_75t_R g986 ( 
.A(n_934),
.Y(n_986)
);

OA21x2_ASAP7_75t_L g987 ( 
.A1(n_928),
.A2(n_910),
.B(n_918),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_950),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_926),
.A2(n_877),
.B(n_47),
.Y(n_989)
);

NOR2xp67_ASAP7_75t_SL g990 ( 
.A(n_959),
.B(n_905),
.Y(n_990)
);

CKINVDCx6p67_ASAP7_75t_R g991 ( 
.A(n_935),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_924),
.B(n_905),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_960),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_944),
.A2(n_48),
.B(n_41),
.Y(n_994)
);

AOI21x1_ASAP7_75t_L g995 ( 
.A1(n_937),
.A2(n_397),
.B(n_383),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_939),
.A2(n_220),
.B(n_294),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_958),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_927),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_965),
.A2(n_218),
.B(n_291),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_924),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_932),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_963),
.A2(n_214),
.B(n_287),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_930),
.B(n_18),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_991),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_974),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_968),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_988),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_998),
.A2(n_925),
.B1(n_946),
.B2(n_919),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_970),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_976),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_1003),
.A2(n_954),
.B1(n_952),
.B2(n_955),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_969),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_983),
.B(n_955),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_987),
.A2(n_949),
.B1(n_947),
.B2(n_964),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_973),
.Y(n_1015)
);

AND2x6_ASAP7_75t_L g1016 ( 
.A(n_980),
.B(n_1001),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_967),
.B(n_971),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_1003),
.A2(n_993),
.B1(n_988),
.B2(n_967),
.Y(n_1018)
);

BUFx12f_ASAP7_75t_L g1019 ( 
.A(n_992),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_987),
.A2(n_428),
.B1(n_454),
.B2(n_452),
.Y(n_1020)
);

CKINVDCx16_ASAP7_75t_R g1021 ( 
.A(n_992),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_986),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_997),
.B(n_18),
.Y(n_1023)
);

OAI221xp5_ASAP7_75t_L g1024 ( 
.A1(n_987),
.A2(n_426),
.B1(n_448),
.B2(n_444),
.C(n_443),
.Y(n_1024)
);

BUFx8_ASAP7_75t_L g1025 ( 
.A(n_974),
.Y(n_1025)
);

NAND3xp33_ASAP7_75t_L g1026 ( 
.A(n_984),
.B(n_419),
.C(n_441),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_974),
.Y(n_1027)
);

OAI221xp5_ASAP7_75t_L g1028 ( 
.A1(n_984),
.A2(n_415),
.B1(n_439),
.B2(n_436),
.C(n_434),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_1000),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_984),
.A2(n_413),
.B1(n_432),
.B2(n_431),
.Y(n_1030)
);

OAI221xp5_ASAP7_75t_L g1031 ( 
.A1(n_971),
.A2(n_412),
.B1(n_427),
.B2(n_421),
.C(n_414),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_986),
.B(n_19),
.Y(n_1032)
);

CKINVDCx11_ASAP7_75t_R g1033 ( 
.A(n_974),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_979),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_979),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_972),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_980),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_SL g1038 ( 
.A1(n_978),
.A2(n_409),
.B1(n_407),
.B2(n_406),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1001),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_989),
.A2(n_932),
.B(n_405),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_977),
.Y(n_1041)
);

AO21x2_ASAP7_75t_L g1042 ( 
.A1(n_1040),
.A2(n_995),
.B(n_966),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_1019),
.Y(n_1043)
);

AOI211xp5_ASAP7_75t_L g1044 ( 
.A1(n_1011),
.A2(n_978),
.B(n_990),
.C(n_985),
.Y(n_1044)
);

CKINVDCx14_ASAP7_75t_R g1045 ( 
.A(n_1004),
.Y(n_1045)
);

OAI221xp5_ASAP7_75t_L g1046 ( 
.A1(n_1008),
.A2(n_969),
.B1(n_982),
.B2(n_1002),
.C(n_996),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_1011),
.A2(n_977),
.B1(n_981),
.B2(n_969),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_1024),
.A2(n_966),
.B1(n_994),
.B2(n_999),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1020),
.A2(n_975),
.B(n_53),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1015),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1006),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_1010),
.B(n_49),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1009),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1032),
.A2(n_54),
.B1(n_59),
.B2(n_62),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1013),
.B(n_63),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1007),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1018),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1037),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1018),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_1029),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1017),
.A2(n_64),
.B(n_70),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1021),
.B(n_71),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1017),
.B(n_73),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1026),
.A2(n_1028),
.B(n_1030),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1023),
.B(n_1027),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1022),
.A2(n_74),
.B1(n_82),
.B2(n_83),
.Y(n_1066)
);

AOI21xp33_ASAP7_75t_L g1067 ( 
.A1(n_1038),
.A2(n_85),
.B(n_88),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_1022),
.A2(n_1031),
.B1(n_1014),
.B2(n_1033),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1005),
.B(n_92),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1039),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1012),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1012),
.A2(n_99),
.B1(n_105),
.B2(n_106),
.Y(n_1072)
);

OAI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1005),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_1073)
);

AOI221xp5_ASAP7_75t_SL g1074 ( 
.A1(n_1034),
.A2(n_113),
.B1(n_115),
.B2(n_117),
.C(n_118),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1035),
.A2(n_120),
.B(n_122),
.C(n_131),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1016),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1005),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_1043),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1051),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1056),
.B(n_1036),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1057),
.B(n_1059),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1053),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1076),
.B(n_1041),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1050),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1058),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1070),
.Y(n_1086)
);

INVxp67_ASAP7_75t_SL g1087 ( 
.A(n_1063),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_1042),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1042),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1065),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1043),
.B(n_1062),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1043),
.B(n_1016),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1046),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1052),
.B(n_1044),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1047),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_1055),
.B(n_136),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1045),
.B(n_1016),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1060),
.B(n_1016),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1069),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1049),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1061),
.B(n_138),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1061),
.B(n_144),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1097),
.B(n_1098),
.Y(n_1103)
);

OAI33xp33_ASAP7_75t_L g1104 ( 
.A1(n_1081),
.A2(n_1073),
.A3(n_1077),
.B1(n_1072),
.B2(n_1071),
.B3(n_1064),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1087),
.A2(n_1073),
.B(n_1075),
.Y(n_1105)
);

NAND2xp33_ASAP7_75t_R g1106 ( 
.A(n_1094),
.B(n_1091),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1079),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_1080),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1101),
.A2(n_1068),
.B1(n_1054),
.B2(n_1066),
.Y(n_1109)
);

NAND4xp25_ASAP7_75t_L g1110 ( 
.A(n_1093),
.B(n_1074),
.C(n_1068),
.D(n_1054),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1095),
.A2(n_1067),
.B1(n_1066),
.B2(n_1048),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_1090),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1093),
.A2(n_1025),
.B1(n_152),
.B2(n_157),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1085),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1105),
.B(n_1087),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1108),
.B(n_1090),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1103),
.B(n_1107),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_1112),
.B(n_1082),
.Y(n_1118)
);

AND2x4_ASAP7_75t_SL g1119 ( 
.A(n_1113),
.B(n_1078),
.Y(n_1119)
);

INVxp67_ASAP7_75t_L g1120 ( 
.A(n_1106),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1114),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_1105),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_1109),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1111),
.B(n_1078),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_1122),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_1116),
.B(n_1086),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1117),
.B(n_1078),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1120),
.B(n_1092),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1118),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1115),
.Y(n_1130)
);

NAND2x1_ASAP7_75t_SL g1131 ( 
.A(n_1124),
.B(n_1101),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1125),
.A2(n_1123),
.B(n_1110),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_SL g1133 ( 
.A1(n_1125),
.A2(n_1123),
.B(n_1100),
.C(n_1096),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1129),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1127),
.B(n_1119),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_R g1136 ( 
.A(n_1130),
.B(n_1102),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_SL g1137 ( 
.A(n_1128),
.B(n_1102),
.C(n_1100),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_1126),
.B(n_1084),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1131),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_1129),
.B(n_1121),
.Y(n_1140)
);

OAI33xp33_ASAP7_75t_L g1141 ( 
.A1(n_1125),
.A2(n_1104),
.A3(n_1089),
.B1(n_1099),
.B2(n_1085),
.B3(n_1088),
.Y(n_1141)
);

OAI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1132),
.A2(n_1099),
.B1(n_1088),
.B2(n_1089),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1134),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1138),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1140),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1136),
.B(n_1083),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1139),
.A2(n_1083),
.B1(n_1025),
.B2(n_168),
.Y(n_1147)
);

OAI31xp33_ASAP7_75t_L g1148 ( 
.A1(n_1142),
.A2(n_1133),
.A3(n_1145),
.B(n_1141),
.Y(n_1148)
);

OAI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1147),
.A2(n_1137),
.B1(n_1135),
.B2(n_1083),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1143),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1144),
.Y(n_1151)
);

NAND2x1_ASAP7_75t_SL g1152 ( 
.A(n_1146),
.B(n_145),
.Y(n_1152)
);

AOI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_1143),
.A2(n_167),
.B(n_170),
.Y(n_1153)
);

NAND2xp33_ASAP7_75t_L g1154 ( 
.A(n_1151),
.B(n_173),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1150),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1148),
.B(n_174),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1152),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1157),
.B(n_1149),
.Y(n_1158)
);

NOR3xp33_ASAP7_75t_L g1159 ( 
.A(n_1156),
.B(n_1153),
.C(n_187),
.Y(n_1159)
);

NAND4xp25_ASAP7_75t_L g1160 ( 
.A(n_1155),
.B(n_186),
.C(n_193),
.D(n_195),
.Y(n_1160)
);

AND4x1_ASAP7_75t_L g1161 ( 
.A(n_1159),
.B(n_1154),
.C(n_197),
.D(n_198),
.Y(n_1161)
);

AOI21xp33_ASAP7_75t_L g1162 ( 
.A1(n_1158),
.A2(n_196),
.B(n_201),
.Y(n_1162)
);

OAI221xp5_ASAP7_75t_L g1163 ( 
.A1(n_1160),
.A2(n_203),
.B1(n_204),
.B2(n_206),
.C(n_207),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1161),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1162),
.A2(n_209),
.B1(n_221),
.B2(n_223),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1164),
.B(n_1163),
.Y(n_1166)
);

NOR2x1_ASAP7_75t_L g1167 ( 
.A(n_1166),
.B(n_1165),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1166),
.A2(n_224),
.B1(n_227),
.B2(n_230),
.Y(n_1168)
);

NOR2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1167),
.B(n_232),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1168),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1170),
.A2(n_1169),
.B(n_236),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1170),
.B(n_235),
.Y(n_1172)
);

OAI22x1_ASAP7_75t_L g1173 ( 
.A1(n_1169),
.A2(n_237),
.B1(n_239),
.B2(n_241),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1173),
.Y(n_1174)
);

XOR2x1_ASAP7_75t_L g1175 ( 
.A(n_1174),
.B(n_1172),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1175),
.A2(n_1171),
.B1(n_244),
.B2(n_248),
.Y(n_1176)
);

AOI21xp33_ASAP7_75t_L g1177 ( 
.A1(n_1176),
.A2(n_243),
.B(n_253),
.Y(n_1177)
);

AOI322xp5_ASAP7_75t_L g1178 ( 
.A1(n_1177),
.A2(n_257),
.A3(n_258),
.B1(n_259),
.B2(n_261),
.C1(n_262),
.C2(n_264),
.Y(n_1178)
);

AOI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_1178),
.A2(n_268),
.B1(n_270),
.B2(n_273),
.C(n_275),
.Y(n_1179)
);

AOI211xp5_ASAP7_75t_L g1180 ( 
.A1(n_1179),
.A2(n_276),
.B(n_277),
.C(n_280),
.Y(n_1180)
);


endmodule