module fake_netlist_6_1135_n_5869 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_706, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_5869);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_706;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_5869;

wire n_5643;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_741;
wire n_1351;
wire n_5254;
wire n_1212;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4395;
wire n_4388;
wire n_1061;
wire n_3089;
wire n_783;
wire n_5653;
wire n_4978;
wire n_5409;
wire n_5301;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_5524;
wire n_5345;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_5818;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5548;
wire n_5057;
wire n_3030;
wire n_830;
wire n_5838;
wire n_5725;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_4273;
wire n_5545;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_5598;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_5819;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_5279;
wire n_2786;
wire n_5239;
wire n_1781;
wire n_1971;
wire n_5354;
wire n_5332;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_5420;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_5638;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_5684;
wire n_5729;
wire n_5680;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_5522;
wire n_5828;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_5493;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_5452;
wire n_3888;
wire n_764;
wire n_5476;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_5536;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_5532;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_5609;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_5658;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_5667;
wire n_780;
wire n_2624;
wire n_5865;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_5281;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_5314;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_5795;
wire n_4473;
wire n_5552;
wire n_5226;
wire n_890;
wire n_5457;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_2712;
wire n_5529;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_925;
wire n_1932;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_5787;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_5445;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5501;
wire n_5342;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_5748;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_5636;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_989;
wire n_2689;
wire n_1473;
wire n_5286;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_5811;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_1004;
wire n_1529;
wire n_5530;
wire n_2473;
wire n_5397;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_5595;
wire n_3119;
wire n_5427;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_5388;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_5599;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_5326;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_1398;
wire n_1201;
wire n_884;
wire n_5394;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_5359;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_5741;
wire n_2773;
wire n_5405;
wire n_5288;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_5761;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_5760;
wire n_2146;
wire n_2131;
wire n_5472;
wire n_3547;
wire n_5679;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_5688;
wire n_5740;
wire n_1731;
wire n_5820;
wire n_5648;
wire n_2135;
wire n_5745;
wire n_4707;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_5180;
wire n_858;
wire n_2049;
wire n_5182;
wire n_956;
wire n_5534;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_5660;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_5334;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_5783;
wire n_3120;
wire n_5821;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_5556;
wire n_4932;
wire n_5456;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_5500;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_5433;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_5618;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_5689;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_5641;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_5731;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_5754;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_5629;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_5434;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_5852;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_5358;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_5571;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_5512;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_5607;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_5562;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_5622;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_5577;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_5413;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_5779;
wire n_2020;
wire n_1643;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_4027;
wire n_763;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_5591;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_5518;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_5847;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_5541;
wire n_5568;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_5381;
wire n_2408;
wire n_5723;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_5696;
wire n_4486;
wire n_1816;
wire n_5848;
wire n_3024;
wire n_4612;
wire n_5673;
wire n_5443;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_5485;
wire n_5823;
wire n_2800;
wire n_3496;
wire n_5473;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_5537;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_3101;
wire n_1574;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_5630;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_5379;
wire n_5335;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_5424;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_5505;
wire n_5868;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_5018;
wire n_3896;
wire n_3815;
wire n_5274;
wire n_3274;
wire n_5401;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_5769;
wire n_4794;
wire n_722;
wire n_5613;
wire n_5612;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_5581;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_5375;
wire n_2451;
wire n_5370;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_5601;
wire n_5784;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_5248;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_5635;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_5528;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_873;
wire n_3946;
wire n_2989;
wire n_5778;
wire n_3395;
wire n_4474;
wire n_5665;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_5788;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_5317;
wire n_1094;
wire n_5430;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_5540;
wire n_3532;
wire n_5716;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_5762;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_808;
wire n_5519;
wire n_4047;
wire n_5753;
wire n_3413;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_4320;
wire n_3884;
wire n_5808;
wire n_5436;
wire n_5139;
wire n_757;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_5789;
wire n_2104;
wire n_3883;
wire n_5866;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5822;
wire n_5195;
wire n_3949;
wire n_5726;
wire n_2792;
wire n_5364;
wire n_3315;
wire n_5533;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_5718;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4526;
wire n_4277;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_5792;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_5554;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_5553;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_5711;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_5790;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_3917;
wire n_2347;
wire n_816;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_5404;
wire n_2916;
wire n_5739;
wire n_4292;
wire n_2467;
wire n_5549;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_3280;
wire n_5757;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_950;
wire n_3009;
wire n_5824;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_5488;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_5637;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_5728;
wire n_5471;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_5843;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_5484;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_5523;
wire n_1067;
wire n_3405;
wire n_5423;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_5204;
wire n_5333;
wire n_847;
wire n_851;
wire n_4991;
wire n_5594;
wire n_2554;
wire n_5422;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_5526;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_5551;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_5257;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4753;
wire n_4688;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_5631;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_5854;
wire n_2667;
wire n_5460;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_5686;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_2848;
wire n_1849;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5465;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_796;
wire n_1195;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_5721;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_5719;
wire n_1502;
wire n_5773;
wire n_1659;
wire n_5482;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_5793;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_5578;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5742;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_5676;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_5674;
wire n_3270;
wire n_5539;
wire n_2846;
wire n_5282;
wire n_970;
wire n_2488;
wire n_1980;
wire n_5464;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_5589;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_5475;
wire n_5807;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_4386;
wire n_2995;
wire n_5273;
wire n_1437;
wire n_4844;
wire n_4438;
wire n_4836;
wire n_5439;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_856;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_5706;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_5431;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_5627;
wire n_5774;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_5798;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_1508;
wire n_5621;
wire n_5608;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_5844;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_5867;
wire n_750;
wire n_5508;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_5597;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_5515;
wire n_1997;
wire n_5662;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_5862;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_5697;
wire n_3416;
wire n_3498;
wire n_5767;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_5462;
wire n_1497;
wire n_3672;
wire n_5318;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4192;
wire n_4109;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_5585;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_5348;
wire n_1332;
wire n_5480;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_936;
wire n_3045;
wire n_3821;
wire n_885;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_5461;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_5503;
wire n_5845;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_5600;
wire n_5755;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_5448;
wire n_2939;
wire n_5749;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_1650;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_5418;
wire n_4088;
wire n_3398;
wire n_5685;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_5459;
wire n_1019;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_5839;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_5514;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_5351;
wire n_4543;
wire n_740;
wire n_4157;
wire n_4229;
wire n_5293;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_5400;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_832;
wire n_3049;
wire n_5389;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_5623;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_5693;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_5663;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_5647;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_5203;
wire n_930;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_5426;
wire n_1656;
wire n_5803;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_5285;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_5365;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_5715;
wire n_4920;
wire n_870;
wire n_5395;
wire n_1253;
wire n_5709;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_5634;
wire n_5672;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_5799;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_5617;
wire n_1829;
wire n_5266;
wire n_5580;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_5390;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_5593;
wire n_4769;
wire n_5764;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_5385;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_5853;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5376;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_5561;
wire n_5410;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_5378;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_5691;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_5615;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_5468;
wire n_4730;
wire n_5399;
wire n_1234;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_1003;
wire n_5713;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_5550;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_5573;
wire n_1553;
wire n_5509;
wire n_5382;
wire n_5659;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_5863;
wire n_2645;
wire n_3904;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_5466;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_1056;
wire n_758;
wire n_5851;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_5796;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_5492;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_5829;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_5734;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_5770;
wire n_1333;
wire n_2496;
wire n_5705;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_5525;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_3943;
wire n_2300;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_5374;
wire n_5575;
wire n_1843;
wire n_5675;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_5297;
wire n_1309;
wire n_1123;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_5642;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_5302;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_5639;
wire n_5781;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_5543;
wire n_1251;
wire n_5361;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_1312;
wire n_5668;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_5463;
wire n_3022;
wire n_5489;
wire n_1165;
wire n_4773;
wire n_5654;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_5479;
wire n_3549;
wire n_5714;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_5510;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_5692;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_5555;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_825;
wire n_3785;
wire n_2963;
wire n_5366;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_5415;
wire n_5419;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_5732;
wire n_5372;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_5690;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_5801;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5347;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_5656;
wire n_1469;
wire n_5125;
wire n_5857;
wire n_2650;
wire n_5652;
wire n_987;
wire n_5499;
wire n_720;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_5507;
wire n_1809;
wire n_5569;
wire n_4280;
wire n_1181;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_5455;
wire n_5442;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_5511;
wire n_2898;
wire n_5295;
wire n_2368;
wire n_4175;
wire n_5490;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_5836;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_5834;
wire n_3191;
wire n_5584;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_1207;
wire n_5707;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_5497;
wire n_880;
wire n_3505;
wire n_3540;
wire n_3577;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_5481;
wire n_3590;
wire n_2435;
wire n_5344;
wire n_954;
wire n_4419;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_5794;
wire n_1382;
wire n_5408;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_5271;
wire n_2323;
wire n_2784;
wire n_5494;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_3755;
wire n_1125;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_5467;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5827;
wire n_5199;
wire n_3407;
wire n_5313;
wire n_3856;
wire n_1185;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_5513;
wire n_5614;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_3243;
wire n_2462;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_5835;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_5846;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_5592;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_5278;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_2993;
wire n_3016;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_5708;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_5474;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_5649;
wire n_1905;
wire n_3466;
wire n_762;
wire n_5704;
wire n_4983;
wire n_1778;
wire n_5287;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_5516;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_5698;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_5771;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_5538;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_5428;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_5677;
wire n_4124;
wire n_5570;
wire n_785;
wire n_5153;
wire n_4611;
wire n_5435;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_5566;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_5487;
wire n_5486;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_5391;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_5849;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_5574;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_5469;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_5804;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_5682;
wire n_5387;
wire n_5557;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_5681;
wire n_1271;
wire n_4901;
wire n_4145;
wire n_4821;
wire n_1545;
wire n_3121;
wire n_4040;
wire n_1640;
wire n_2406;
wire n_806;
wire n_2141;
wire n_5316;
wire n_5703;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_5564;
wire n_5620;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_5406;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_5724;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_5806;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_5738;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_5710;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_5517;
wire n_3207;
wire n_5605;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_5746;
wire n_2045;
wire n_817;
wire n_5451;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_5417;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_5864;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_5432;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_5453;
wire n_3658;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_5842;
wire n_5814;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_5699;
wire n_5531;
wire n_5765;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_5777;
wire n_4225;
wire n_747;
wire n_2565;
wire n_5495;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5655;
wire n_5064;
wire n_5610;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_5759;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_957;
wire n_1994;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_5559;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_5786;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_5737;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_5768;
wire n_3553;
wire n_2465;
wire n_2275;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_3494;
wire n_1721;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_5350;
wire n_5470;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_5858;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_5700;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_904;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_5588;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_5736;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_5478;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_5832;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_5812;
wire n_2540;
wire n_973;
wire n_5743;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_5368;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_5782;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_5563;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_5840;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_5717;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_5720;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_3626;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_5650;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_5567;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_5625;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_5022;
wire n_5670;
wire n_1280;
wire n_3296;
wire n_5276;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_5238;
wire n_5855;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_5429;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_5535;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_821;
wire n_4372;
wire n_1068;
wire n_982;
wire n_5640;
wire n_932;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_5560;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_5544;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_5744;
wire n_4013;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_5841;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_5611;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_5701;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_5502;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_5850;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_5521;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_5856;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_5837;
wire n_4675;
wire n_2663;
wire n_5825;
wire n_4018;
wire n_5491;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_5496;
wire n_5802;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_5547;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_5596;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_5604;
wire n_1756;
wire n_1128;
wire n_5411;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_5815;
wire n_4191;
wire n_5695;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_5331;
wire n_4330;
wire n_5311;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_5797;
wire n_4240;
wire n_3491;
wire n_5572;
wire n_1488;
wire n_2148;
wire n_4162;
wire n_5565;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_5520;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_5800;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_5669;
wire n_5772;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_5758;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_5603;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_5763;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_5751;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_1505;
wire n_5712;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_4871;
wire n_2403;
wire n_1070;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_5449;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1774;
wire n_1475;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_5398;
wire n_5860;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_5583;
wire n_4654;
wire n_3640;
wire n_1159;
wire n_995;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_5775;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2720;
wire n_2204;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_5483;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_5785;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_5780;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_994;
wire n_5735;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_5752;
wire n_1661;
wire n_5360;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_5632;
wire n_5582;
wire n_5425;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_5446;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_5678;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_3784;
wire n_5437;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_5454;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_5407;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_5810;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_5702;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_5590;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_5809;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_5349;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_5813;
wire n_790;
wire n_5833;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_5616;
wire n_5805;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_5816;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_5416;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_5167;
wire n_5661;
wire n_5830;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_5558;
wire n_1826;
wire n_5687;
wire n_5383;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5587;
wire n_5236;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_5651;
wire n_4630;
wire n_1217;
wire n_5645;
wire n_3990;
wire n_1628;
wire n_5766;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_5671;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_5412;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_5733;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_5791;
wire n_5727;
wire n_761;
wire n_2492;
wire n_3778;
wire n_5328;
wire n_5657;
wire n_1173;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_5602;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_5579;
wire n_1922;
wire n_5750;
wire n_4823;
wire n_5831;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_5666;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_5546;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_5626;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_5633;
wire n_5664;
wire n_1218;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_3764;
wire n_2360;
wire n_4784;
wire n_4075;
wire n_5340;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_5280;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_5369;
wire n_975;
wire n_5730;
wire n_5576;
wire n_3359;
wire n_5272;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_5646;
wire n_5624;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_2280;
wire n_1557;
wire n_3945;
wire n_730;
wire n_5817;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_5586;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_5861;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_5619;
wire n_3965;
wire n_5859;
wire n_5380;
wire n_4500;
wire n_5065;
wire n_862;
wire n_5776;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_5606;
wire n_5644;
wire n_2813;
wire n_1935;
wire n_5826;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_5683;
wire n_2677;
wire n_3182;
wire n_5756;
wire n_3283;
wire n_5527;
wire n_1742;
wire n_4030;

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_30),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_294),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_251),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_543),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_202),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_117),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_160),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_533),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_496),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_525),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_694),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_302),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_237),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_361),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_349),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_194),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_151),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_100),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_504),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_506),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_280),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_400),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_158),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_253),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_323),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_150),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_194),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_294),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_704),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_406),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_63),
.Y(n_738)
);

BUFx5_ASAP7_75t_L g739 ( 
.A(n_559),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_98),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_393),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_52),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_648),
.Y(n_743)
);

BUFx10_ASAP7_75t_L g744 ( 
.A(n_483),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_465),
.Y(n_745)
);

BUFx10_ASAP7_75t_L g746 ( 
.A(n_10),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_37),
.Y(n_747)
);

BUFx5_ASAP7_75t_L g748 ( 
.A(n_89),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_364),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_373),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_355),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_324),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_537),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_695),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_400),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_252),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_649),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_620),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_241),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_59),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_203),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_52),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_140),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_411),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_459),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_205),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_554),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_156),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_266),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_349),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_412),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_149),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_690),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_370),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_364),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_677),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_627),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_214),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_247),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_312),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_242),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_115),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_113),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_328),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_264),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_567),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_609),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_48),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_160),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_701),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_634),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_431),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_312),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_506),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_697),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_326),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_380),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_693),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_381),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_485),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_428),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_410),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_559),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_44),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_269),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_584),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_680),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_628),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_590),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_360),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_245),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_139),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_367),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_687),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_582),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_93),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_205),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_167),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_394),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_392),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_85),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_110),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_10),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_657),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_475),
.Y(n_825)
);

BUFx8_ASAP7_75t_SL g826 ( 
.A(n_137),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_503),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_605),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_180),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_206),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_33),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_570),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_566),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_614),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_157),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_100),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_245),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_109),
.Y(n_838)
);

CKINVDCx16_ASAP7_75t_R g839 ( 
.A(n_339),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_44),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_38),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_304),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_204),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_240),
.Y(n_844)
);

CKINVDCx14_ASAP7_75t_R g845 ( 
.A(n_115),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_78),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_480),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_149),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_566),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_686),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_522),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_407),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_351),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_551),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_564),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_666),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_169),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_707),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_110),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_227),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_629),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_514),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_589),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_624),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_111),
.Y(n_865)
);

INVxp33_ASAP7_75t_SL g866 ( 
.A(n_596),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_700),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_240),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_631),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_345),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_667),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_682),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_59),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_706),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_505),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_683),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_255),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_255),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_621),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_365),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_101),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_702),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_401),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_318),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_553),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_674),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_624),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_341),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_389),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_154),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_604),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_698),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_81),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_57),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_306),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_481),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_592),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_498),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_417),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_540),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_350),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_156),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_252),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_188),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_552),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_473),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_29),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_515),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_496),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_637),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_113),
.Y(n_911)
);

INVxp67_ASAP7_75t_SL g912 ( 
.A(n_270),
.Y(n_912)
);

BUFx10_ASAP7_75t_L g913 ( 
.A(n_143),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_601),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_47),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_572),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_65),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_696),
.Y(n_918)
);

BUFx5_ASAP7_75t_L g919 ( 
.A(n_336),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_134),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_625),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_560),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_397),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_22),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_514),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_324),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_705),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_327),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_106),
.Y(n_929)
);

BUFx5_ASAP7_75t_L g930 ( 
.A(n_375),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_237),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_509),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_225),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_304),
.Y(n_934)
);

BUFx10_ASAP7_75t_L g935 ( 
.A(n_441),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_105),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_703),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_128),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_597),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_626),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_444),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_456),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_492),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_466),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_176),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_287),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_617),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_550),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_654),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_169),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_27),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_158),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_502),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_644),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_38),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_27),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_675),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_293),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_383),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_132),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_286),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_204),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_551),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_154),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_585),
.Y(n_965)
);

BUFx8_ASAP7_75t_SL g966 ( 
.A(n_231),
.Y(n_966)
);

INVx1_ASAP7_75t_SL g967 ( 
.A(n_19),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_317),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_454),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_96),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_587),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_306),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_609),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_322),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_323),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_25),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_673),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_191),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_553),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_623),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_480),
.Y(n_981)
);

CKINVDCx16_ASAP7_75t_R g982 ( 
.A(n_218),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_103),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_182),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_587),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_254),
.Y(n_986)
);

CKINVDCx14_ASAP7_75t_R g987 ( 
.A(n_611),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_630),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_585),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_465),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_628),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_595),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_526),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_636),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_466),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_217),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_277),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_421),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_435),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_692),
.Y(n_1000)
);

BUFx10_ASAP7_75t_L g1001 ( 
.A(n_87),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_173),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_278),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_554),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_536),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_260),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_362),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_610),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_463),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_81),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_102),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_259),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_437),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_102),
.Y(n_1014)
);

BUFx10_ASAP7_75t_L g1015 ( 
.A(n_139),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_143),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_542),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_604),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_664),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_405),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_535),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_247),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_484),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_2),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_82),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_340),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_270),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_556),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_197),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_478),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_203),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_503),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_478),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_342),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_616),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_578),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_558),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_699),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_273),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_48),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_591),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_456),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_357),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_311),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_13),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_6),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_72),
.Y(n_1047)
);

CKINVDCx16_ASAP7_75t_R g1048 ( 
.A(n_217),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_225),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_334),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_429),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_534),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_632),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_122),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_123),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_577),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_661),
.Y(n_1057)
);

CKINVDCx12_ASAP7_75t_R g1058 ( 
.A(n_337),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_16),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_31),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_121),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_626),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_447),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_82),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_392),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_416),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_528),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_529),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_688),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_60),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_360),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_643),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_507),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_461),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_381),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_603),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_438),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_268),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_321),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_363),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_660),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_658),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_107),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_519),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_131),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_663),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_571),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_398),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_292),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_470),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_99),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_424),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_412),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_490),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_232),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_477),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_612),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_162),
.Y(n_1098)
);

CKINVDCx14_ASAP7_75t_R g1099 ( 
.A(n_406),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_384),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_33),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_403),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_475),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_535),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_219),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_233),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_414),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_170),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_399),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_647),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_596),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_74),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_284),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_541),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_200),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_219),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_65),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_620),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_277),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_574),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_579),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_358),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_348),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_571),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_355),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_128),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_386),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_689),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_460),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_366),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_483),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_328),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_569),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_290),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_157),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_415),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_417),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_564),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_9),
.Y(n_1139)
);

INVxp67_ASAP7_75t_L g1140 ( 
.A(n_62),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_133),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_182),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_619),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_653),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_91),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_326),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_607),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_691),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_505),
.Y(n_1149)
);

BUFx5_ASAP7_75t_L g1150 ( 
.A(n_299),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_479),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_501),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_420),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_303),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_301),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_130),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_185),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_633),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_433),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_216),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_380),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_548),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_592),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_408),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_69),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_409),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_191),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_685),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_404),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_565),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_34),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_250),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_455),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_537),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_534),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_226),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_538),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_530),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_283),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_432),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_78),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_568),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_147),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_168),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_230),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_335),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_276),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_488),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_242),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_446),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_290),
.Y(n_1191)
);

INVxp33_ASAP7_75t_R g1192 ( 
.A(n_179),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_315),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_253),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_679),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_85),
.Y(n_1196)
);

CKINVDCx16_ASAP7_75t_R g1197 ( 
.A(n_484),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_50),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_621),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_578),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_597),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_369),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_361),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_580),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_57),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_464),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_358),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_313),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_615),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_80),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_159),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_343),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_558),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_267),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_333),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_0),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_296),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_441),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_335),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_359),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_254),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_45),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_76),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_497),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_363),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_611),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_573),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_75),
.Y(n_1228)
);

CKINVDCx16_ASAP7_75t_R g1229 ( 
.A(n_16),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_159),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_271),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_288),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_652),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_166),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_606),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_487),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_195),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_569),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_739),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_882),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_739),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_882),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_826),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_739),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_739),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_739),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_739),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_739),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_966),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_739),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_739),
.Y(n_1251)
);

BUFx10_ASAP7_75t_L g1252 ( 
.A(n_716),
.Y(n_1252)
);

INVxp67_ASAP7_75t_L g1253 ( 
.A(n_724),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_748),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_748),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_748),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_748),
.Y(n_1257)
);

CKINVDCx14_ASAP7_75t_R g1258 ( 
.A(n_845),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_987),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_748),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_748),
.Y(n_1261)
);

INVxp33_ASAP7_75t_SL g1262 ( 
.A(n_779),
.Y(n_1262)
);

INVxp33_ASAP7_75t_L g1263 ( 
.A(n_830),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_748),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_748),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_715),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_919),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_919),
.Y(n_1268)
);

CKINVDCx16_ASAP7_75t_R g1269 ( 
.A(n_839),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_919),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_919),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_919),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_745),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1099),
.Y(n_1274)
);

CKINVDCx14_ASAP7_75t_R g1275 ( 
.A(n_718),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_724),
.B(n_775),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_737),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_743),
.B(n_1),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_919),
.Y(n_1279)
);

BUFx5_ASAP7_75t_L g1280 ( 
.A(n_776),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_919),
.Y(n_1281)
);

INVxp33_ASAP7_75t_SL g1282 ( 
.A(n_775),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_982),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_919),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1097),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_919),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_930),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_930),
.Y(n_1288)
);

BUFx2_ASAP7_75t_SL g1289 ( 
.A(n_798),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_930),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_930),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_930),
.Y(n_1292)
);

NOR2xp67_ASAP7_75t_L g1293 ( 
.A(n_730),
.B(n_0),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_858),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_930),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_930),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1097),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_930),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_930),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1150),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1150),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1150),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1048),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1150),
.Y(n_1304)
);

CKINVDCx16_ASAP7_75t_R g1305 ( 
.A(n_1197),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_761),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1150),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_730),
.Y(n_1308)
);

CKINVDCx16_ASAP7_75t_R g1309 ( 
.A(n_1229),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_776),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_708),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1222),
.Y(n_1312)
);

CKINVDCx16_ASAP7_75t_R g1313 ( 
.A(n_744),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1150),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1150),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1150),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1150),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_795),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_795),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_712),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_874),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_874),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_910),
.Y(n_1323)
);

INVxp33_ASAP7_75t_SL g1324 ( 
.A(n_1222),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_730),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_910),
.Y(n_1326)
);

INVxp33_ASAP7_75t_L g1327 ( 
.A(n_709),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_949),
.Y(n_1328)
);

CKINVDCx16_ASAP7_75t_R g1329 ( 
.A(n_744),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_949),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_871),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_977),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_977),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_994),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_994),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1000),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1000),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_709),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_717),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1081),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1081),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1128),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_793),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1128),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1144),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1144),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1148),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1148),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1233),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_719),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_793),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1233),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_785),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_793),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_871),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1119),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1119),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1119),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_781),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_781),
.Y(n_1360)
);

CKINVDCx14_ASAP7_75t_R g1361 ( 
.A(n_736),
.Y(n_1361)
);

INVxp33_ASAP7_75t_L g1362 ( 
.A(n_711),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_720),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_721),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_859),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_846),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_744),
.Y(n_1367)
);

INVxp33_ASAP7_75t_L g1368 ( 
.A(n_711),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_859),
.Y(n_1369)
);

INVxp33_ASAP7_75t_SL g1370 ( 
.A(n_722),
.Y(n_1370)
);

INVxp33_ASAP7_75t_L g1371 ( 
.A(n_713),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_847),
.Y(n_1372)
);

INVxp33_ASAP7_75t_SL g1373 ( 
.A(n_723),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_743),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_921),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_725),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_921),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_997),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_731),
.Y(n_1379)
);

INVxp33_ASAP7_75t_L g1380 ( 
.A(n_713),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_997),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1044),
.Y(n_1382)
);

INVxp67_ASAP7_75t_SL g1383 ( 
.A(n_850),
.Y(n_1383)
);

INVxp67_ASAP7_75t_SL g1384 ( 
.A(n_737),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_904),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_737),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_714),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1044),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1073),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_943),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1073),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1101),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_735),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1101),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_737),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_737),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_747),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_747),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_747),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_747),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_747),
.Y(n_1401)
);

INVxp67_ASAP7_75t_SL g1402 ( 
.A(n_819),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_819),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_754),
.B(n_1),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1058),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_819),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_819),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_819),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_855),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_855),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_855),
.Y(n_1411)
);

INVxp33_ASAP7_75t_SL g1412 ( 
.A(n_738),
.Y(n_1412)
);

INVxp33_ASAP7_75t_SL g1413 ( 
.A(n_740),
.Y(n_1413)
);

INVxp33_ASAP7_75t_SL g1414 ( 
.A(n_741),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_855),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_855),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_757),
.B(n_2),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_857),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_742),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_857),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_857),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_857),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_714),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_857),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_905),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_958),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_773),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_905),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_749),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_905),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_905),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_905),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_965),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_750),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_965),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_965),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_965),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_752),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_965),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_979),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_979),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_979),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_983),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_979),
.Y(n_1444)
);

INVxp33_ASAP7_75t_L g1445 ( 
.A(n_726),
.Y(n_1445)
);

INVxp67_ASAP7_75t_L g1446 ( 
.A(n_726),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_979),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1163),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1163),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1163),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1163),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1163),
.Y(n_1452)
);

INVxp33_ASAP7_75t_SL g1453 ( 
.A(n_753),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1178),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1178),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1178),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1178),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_984),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_763),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_764),
.Y(n_1460)
);

BUFx2_ASAP7_75t_SL g1461 ( 
.A(n_807),
.Y(n_1461)
);

INVxp67_ASAP7_75t_SL g1462 ( 
.A(n_1178),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1188),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1188),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1188),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1188),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1188),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1230),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1230),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1230),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_769),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1028),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1230),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1230),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1037),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_863),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_864),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_1046),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_728),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_869),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_873),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1102),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_770),
.Y(n_1483)
);

INVxp33_ASAP7_75t_SL g1484 ( 
.A(n_771),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1105),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1106),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1108),
.Y(n_1487)
);

INVxp67_ASAP7_75t_SL g1488 ( 
.A(n_1032),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_790),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1109),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_728),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_729),
.Y(n_1492)
);

INVxp33_ASAP7_75t_L g1493 ( 
.A(n_729),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_774),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_727),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_732),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_732),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_710),
.B(n_3),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_733),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_733),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_777),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_734),
.Y(n_1502)
);

INVxp33_ASAP7_75t_L g1503 ( 
.A(n_734),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_751),
.Y(n_1504)
);

INVxp33_ASAP7_75t_L g1505 ( 
.A(n_751),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_778),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_756),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_756),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_758),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_782),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_727),
.Y(n_1511)
);

CKINVDCx16_ASAP7_75t_R g1512 ( 
.A(n_744),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_783),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_758),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_759),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_759),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_791),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_762),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1078),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_786),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_762),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_755),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_1088),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_765),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_755),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_765),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_766),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_760),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_766),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_767),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_767),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_768),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_768),
.Y(n_1533)
);

INVxp33_ASAP7_75t_SL g1534 ( 
.A(n_788),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_772),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_772),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1058),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_760),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_784),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_784),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_814),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_787),
.Y(n_1542)
);

CKINVDCx16_ASAP7_75t_R g1543 ( 
.A(n_746),
.Y(n_1543)
);

INVxp67_ASAP7_75t_SL g1544 ( 
.A(n_1121),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_787),
.Y(n_1545)
);

CKINVDCx16_ASAP7_75t_R g1546 ( 
.A(n_746),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_789),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_780),
.Y(n_1548)
);

INVxp67_ASAP7_75t_SL g1549 ( 
.A(n_1140),
.Y(n_1549)
);

CKINVDCx20_ASAP7_75t_R g1550 ( 
.A(n_1098),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_789),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_804),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_804),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_805),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_792),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_805),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_808),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_808),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_810),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_810),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_815),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_815),
.Y(n_1562)
);

INVxp67_ASAP7_75t_SL g1563 ( 
.A(n_912),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_822),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_822),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_794),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_825),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_825),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_827),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_827),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_828),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_828),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_835),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_835),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_796),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_837),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_837),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_824),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_780),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_797),
.Y(n_1580)
);

INVxp33_ASAP7_75t_SL g1581 ( 
.A(n_799),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_840),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_840),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_841),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_841),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_849),
.Y(n_1586)
);

INVxp67_ASAP7_75t_SL g1587 ( 
.A(n_820),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_849),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_852),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_852),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_890),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_890),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_867),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_897),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_897),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_900),
.Y(n_1596)
);

CKINVDCx16_ASAP7_75t_R g1597 ( 
.A(n_746),
.Y(n_1597)
);

INVxp33_ASAP7_75t_L g1598 ( 
.A(n_900),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_820),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_834),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_901),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_901),
.Y(n_1602)
);

INVxp67_ASAP7_75t_SL g1603 ( 
.A(n_834),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_902),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_1132),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_902),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_907),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_907),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_911),
.Y(n_1609)
);

BUFx3_ASAP7_75t_L g1610 ( 
.A(n_872),
.Y(n_1610)
);

CKINVDCx14_ASAP7_75t_R g1611 ( 
.A(n_886),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_800),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_911),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_801),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_914),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_914),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_892),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_802),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_926),
.Y(n_1619)
);

CKINVDCx16_ASAP7_75t_R g1620 ( 
.A(n_746),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_926),
.Y(n_1621)
);

INVxp33_ASAP7_75t_L g1622 ( 
.A(n_940),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_940),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_941),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_941),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_942),
.Y(n_1626)
);

CKINVDCx16_ASAP7_75t_R g1627 ( 
.A(n_913),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_942),
.Y(n_1628)
);

INVxp33_ASAP7_75t_L g1629 ( 
.A(n_945),
.Y(n_1629)
);

INVxp33_ASAP7_75t_SL g1630 ( 
.A(n_803),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_927),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_945),
.Y(n_1632)
);

INVxp67_ASAP7_75t_SL g1633 ( 
.A(n_865),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1133),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_948),
.Y(n_1635)
);

INVxp33_ASAP7_75t_SL g1636 ( 
.A(n_806),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_809),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1146),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_865),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_948),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_960),
.Y(n_1641)
);

CKINVDCx16_ASAP7_75t_R g1642 ( 
.A(n_913),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_1149),
.Y(n_1643)
);

BUFx6f_ASAP7_75t_L g1644 ( 
.A(n_868),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_960),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_961),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_868),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_811),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_961),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_812),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_813),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_816),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_963),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_817),
.Y(n_1654)
);

CKINVDCx16_ASAP7_75t_R g1655 ( 
.A(n_913),
.Y(n_1655)
);

INVxp33_ASAP7_75t_SL g1656 ( 
.A(n_821),
.Y(n_1656)
);

CKINVDCx16_ASAP7_75t_R g1657 ( 
.A(n_913),
.Y(n_1657)
);

INVxp33_ASAP7_75t_L g1658 ( 
.A(n_963),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_969),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_1153),
.Y(n_1660)
);

CKINVDCx16_ASAP7_75t_R g1661 ( 
.A(n_935),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_969),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_975),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_975),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_985),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_985),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_823),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_829),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_908),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_991),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_991),
.Y(n_1671)
);

INVxp33_ASAP7_75t_SL g1672 ( 
.A(n_831),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_908),
.Y(n_1673)
);

BUFx2_ASAP7_75t_SL g1674 ( 
.A(n_876),
.Y(n_1674)
);

INVxp67_ASAP7_75t_SL g1675 ( 
.A(n_931),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_993),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_993),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_832),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_996),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1427),
.B(n_937),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1439),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1427),
.B(n_954),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1439),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1278),
.B(n_866),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1439),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1489),
.B(n_856),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1439),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_1440),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1440),
.Y(n_1689)
);

BUFx6f_ASAP7_75t_L g1690 ( 
.A(n_1440),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1258),
.B(n_935),
.Y(n_1691)
);

CKINVDCx20_ASAP7_75t_R g1692 ( 
.A(n_1266),
.Y(n_1692)
);

BUFx12f_ASAP7_75t_L g1693 ( 
.A(n_1243),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1455),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1258),
.B(n_935),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1489),
.B(n_957),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1294),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1517),
.B(n_918),
.Y(n_1698)
);

BUFx12f_ASAP7_75t_L g1699 ( 
.A(n_1243),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1429),
.B(n_935),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1294),
.Y(n_1701)
);

INVx4_ASAP7_75t_L g1702 ( 
.A(n_1517),
.Y(n_1702)
);

BUFx8_ASAP7_75t_L g1703 ( 
.A(n_1367),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1384),
.Y(n_1704)
);

BUFx8_ASAP7_75t_L g1705 ( 
.A(n_1367),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1383),
.B(n_710),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1525),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1285),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1262),
.B(n_1093),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1566),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1541),
.B(n_1057),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1525),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1402),
.Y(n_1713)
);

AND2x6_ASAP7_75t_L g1714 ( 
.A(n_1251),
.B(n_931),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1455),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1283),
.Y(n_1716)
);

BUFx12f_ASAP7_75t_L g1717 ( 
.A(n_1249),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1297),
.Y(n_1718)
);

INVx5_ASAP7_75t_L g1719 ( 
.A(n_1277),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1386),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1386),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1612),
.B(n_1001),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1541),
.B(n_1069),
.Y(n_1723)
);

BUFx8_ASAP7_75t_L g1724 ( 
.A(n_1276),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_1525),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1525),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1578),
.B(n_1093),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_L g1728 ( 
.A(n_1374),
.B(n_1228),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1578),
.B(n_1228),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1637),
.B(n_1001),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1289),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1667),
.B(n_1001),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1593),
.B(n_1072),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1593),
.B(n_938),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1293),
.B(n_1001),
.Y(n_1735)
);

BUFx12f_ASAP7_75t_L g1736 ( 
.A(n_1249),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1563),
.B(n_1015),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1528),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1610),
.B(n_938),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1276),
.B(n_1015),
.Y(n_1740)
);

INVx4_ASAP7_75t_L g1741 ( 
.A(n_1610),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1617),
.B(n_1082),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1461),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1308),
.B(n_1015),
.Y(n_1744)
);

BUFx12f_ASAP7_75t_L g1745 ( 
.A(n_1283),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1303),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1430),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1312),
.Y(n_1748)
);

AND2x6_ASAP7_75t_L g1749 ( 
.A(n_1251),
.B(n_959),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1396),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1617),
.B(n_959),
.Y(n_1751)
);

BUFx12f_ASAP7_75t_L g1752 ( 
.A(n_1303),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1631),
.B(n_1054),
.Y(n_1753)
);

BUFx12f_ASAP7_75t_L g1754 ( 
.A(n_1259),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1405),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1631),
.B(n_1086),
.Y(n_1756)
);

INVx5_ASAP7_75t_L g1757 ( 
.A(n_1277),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1528),
.Y(n_1758)
);

INVx5_ASAP7_75t_L g1759 ( 
.A(n_1277),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1311),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1240),
.B(n_1054),
.Y(n_1761)
);

BUFx2_ASAP7_75t_L g1762 ( 
.A(n_1311),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1240),
.B(n_1096),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1242),
.B(n_1096),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1351),
.B(n_1110),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1275),
.B(n_1158),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1528),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1262),
.B(n_833),
.Y(n_1768)
);

CKINVDCx6p67_ASAP7_75t_R g1769 ( 
.A(n_1269),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1275),
.B(n_1168),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1242),
.B(n_1180),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_L g1772 ( 
.A(n_1528),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1462),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1259),
.B(n_1015),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1396),
.Y(n_1775)
);

BUFx8_ASAP7_75t_L g1776 ( 
.A(n_1498),
.Y(n_1776)
);

AND2x6_ASAP7_75t_L g1777 ( 
.A(n_1257),
.B(n_1180),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1320),
.Y(n_1778)
);

BUFx12f_ASAP7_75t_L g1779 ( 
.A(n_1274),
.Y(n_1779)
);

INVx5_ASAP7_75t_L g1780 ( 
.A(n_1331),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1395),
.Y(n_1781)
);

BUFx6f_ASAP7_75t_L g1782 ( 
.A(n_1579),
.Y(n_1782)
);

INVx5_ASAP7_75t_L g1783 ( 
.A(n_1331),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1320),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1274),
.B(n_1226),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1488),
.B(n_1195),
.Y(n_1786)
);

BUFx12f_ASAP7_75t_L g1787 ( 
.A(n_1252),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_1579),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1370),
.B(n_1373),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1398),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1537),
.B(n_1190),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1370),
.B(n_836),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1397),
.Y(n_1793)
);

AND2x2_ASAP7_75t_R g1794 ( 
.A(n_1282),
.B(n_1192),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1361),
.B(n_838),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1361),
.B(n_842),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1305),
.B(n_1309),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_SL g1798 ( 
.A(n_1313),
.B(n_1019),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1404),
.B(n_1236),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1339),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1579),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1579),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1611),
.B(n_844),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1599),
.Y(n_1804)
);

BUFx6f_ASAP7_75t_L g1805 ( 
.A(n_1599),
.Y(n_1805)
);

INVx5_ASAP7_75t_L g1806 ( 
.A(n_1331),
.Y(n_1806)
);

BUFx6f_ASAP7_75t_L g1807 ( 
.A(n_1599),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1329),
.B(n_818),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1599),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1399),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1373),
.B(n_848),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1400),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1339),
.Y(n_1813)
);

BUFx2_ASAP7_75t_L g1814 ( 
.A(n_1350),
.Y(n_1814)
);

BUFx12f_ASAP7_75t_L g1815 ( 
.A(n_1350),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1639),
.Y(n_1816)
);

INVx3_ASAP7_75t_L g1817 ( 
.A(n_1639),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1417),
.B(n_1224),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1611),
.B(n_851),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1412),
.B(n_853),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1544),
.B(n_854),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1549),
.B(n_1190),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1374),
.B(n_860),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1363),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1363),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1374),
.B(n_861),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1253),
.B(n_1206),
.Y(n_1827)
);

BUFx8_ASAP7_75t_SL g1828 ( 
.A(n_1266),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1397),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1442),
.Y(n_1830)
);

INVx5_ASAP7_75t_L g1831 ( 
.A(n_1331),
.Y(n_1831)
);

BUFx12f_ASAP7_75t_L g1832 ( 
.A(n_1252),
.Y(n_1832)
);

NOR2x1_ASAP7_75t_L g1833 ( 
.A(n_1355),
.B(n_1038),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1374),
.B(n_862),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1412),
.B(n_870),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1359),
.B(n_1206),
.Y(n_1836)
);

BUFx3_ASAP7_75t_L g1837 ( 
.A(n_1360),
.Y(n_1837)
);

INVx5_ASAP7_75t_L g1838 ( 
.A(n_1639),
.Y(n_1838)
);

NAND2xp33_ASAP7_75t_L g1839 ( 
.A(n_1280),
.B(n_1223),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1413),
.B(n_1414),
.Y(n_1840)
);

BUFx6f_ASAP7_75t_L g1841 ( 
.A(n_1639),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1442),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1364),
.B(n_1376),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1364),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1365),
.B(n_875),
.Y(n_1845)
);

BUFx12f_ASAP7_75t_L g1846 ( 
.A(n_1376),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1369),
.B(n_1223),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1413),
.B(n_877),
.Y(n_1848)
);

INVx5_ASAP7_75t_L g1849 ( 
.A(n_1644),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1375),
.B(n_878),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1377),
.B(n_996),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1644),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1378),
.B(n_879),
.Y(n_1853)
);

AND2x6_ASAP7_75t_L g1854 ( 
.A(n_1257),
.B(n_998),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1379),
.B(n_880),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1381),
.B(n_881),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1644),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1382),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1401),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1467),
.Y(n_1860)
);

XOR2xp5_ASAP7_75t_L g1861 ( 
.A(n_1674),
.B(n_1166),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1644),
.Y(n_1862)
);

BUFx3_ASAP7_75t_L g1863 ( 
.A(n_1388),
.Y(n_1863)
);

BUFx3_ASAP7_75t_L g1864 ( 
.A(n_1389),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1379),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_SL g1866 ( 
.A(n_1512),
.B(n_843),
.Y(n_1866)
);

INVx4_ASAP7_75t_L g1867 ( 
.A(n_1393),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1393),
.B(n_883),
.Y(n_1868)
);

INVxp67_ASAP7_75t_L g1869 ( 
.A(n_1391),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1392),
.B(n_998),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1467),
.Y(n_1871)
);

BUFx3_ASAP7_75t_L g1872 ( 
.A(n_1394),
.Y(n_1872)
);

BUFx2_ASAP7_75t_L g1873 ( 
.A(n_1419),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1469),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1469),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1419),
.B(n_884),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1434),
.Y(n_1877)
);

BUFx6f_ASAP7_75t_L g1878 ( 
.A(n_1403),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1406),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1434),
.B(n_885),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1280),
.B(n_887),
.Y(n_1881)
);

AND2x4_ASAP7_75t_L g1882 ( 
.A(n_1310),
.B(n_1004),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1438),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1414),
.B(n_888),
.Y(n_1884)
);

INVx3_ASAP7_75t_L g1885 ( 
.A(n_1495),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1407),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1310),
.B(n_1341),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_1453),
.B(n_889),
.Y(n_1888)
);

XNOR2x2_ASAP7_75t_L g1889 ( 
.A(n_1353),
.B(n_915),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1408),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1438),
.Y(n_1891)
);

INVxp67_ASAP7_75t_L g1892 ( 
.A(n_1341),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1280),
.B(n_891),
.Y(n_1893)
);

INVx4_ASAP7_75t_L g1894 ( 
.A(n_1459),
.Y(n_1894)
);

INVx5_ASAP7_75t_L g1895 ( 
.A(n_1325),
.Y(n_1895)
);

BUFx12f_ASAP7_75t_L g1896 ( 
.A(n_1459),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1409),
.Y(n_1897)
);

INVx5_ASAP7_75t_L g1898 ( 
.A(n_1325),
.Y(n_1898)
);

BUFx2_ASAP7_75t_L g1899 ( 
.A(n_1460),
.Y(n_1899)
);

BUFx6f_ASAP7_75t_L g1900 ( 
.A(n_1410),
.Y(n_1900)
);

BUFx12f_ASAP7_75t_L g1901 ( 
.A(n_1460),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1471),
.B(n_893),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1280),
.B(n_894),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1471),
.B(n_895),
.Y(n_1904)
);

BUFx6f_ASAP7_75t_L g1905 ( 
.A(n_1411),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1483),
.Y(n_1906)
);

INVx3_ASAP7_75t_L g1907 ( 
.A(n_1495),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1483),
.B(n_896),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1280),
.B(n_898),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1415),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1416),
.Y(n_1911)
);

BUFx3_ASAP7_75t_L g1912 ( 
.A(n_1355),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_SL g1913 ( 
.A(n_1543),
.B(n_947),
.Y(n_1913)
);

BUFx8_ASAP7_75t_L g1914 ( 
.A(n_1318),
.Y(n_1914)
);

INVxp67_ASAP7_75t_L g1915 ( 
.A(n_1587),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1494),
.B(n_899),
.Y(n_1916)
);

BUFx8_ASAP7_75t_L g1917 ( 
.A(n_1319),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1280),
.B(n_903),
.Y(n_1918)
);

INVx4_ASAP7_75t_L g1919 ( 
.A(n_1494),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1280),
.B(n_906),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1501),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1354),
.B(n_1004),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1356),
.B(n_1006),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1418),
.Y(n_1924)
);

INVx5_ASAP7_75t_L g1925 ( 
.A(n_1343),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1420),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1453),
.B(n_909),
.Y(n_1927)
);

BUFx12f_ASAP7_75t_L g1928 ( 
.A(n_1252),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_SL g1929 ( 
.A(n_1546),
.B(n_967),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1421),
.B(n_916),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1422),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1424),
.B(n_917),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1358),
.B(n_1006),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1597),
.B(n_1009),
.Y(n_1934)
);

BUFx8_ASAP7_75t_SL g1935 ( 
.A(n_1273),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1484),
.B(n_920),
.Y(n_1936)
);

INVx5_ASAP7_75t_L g1937 ( 
.A(n_1343),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1425),
.Y(n_1938)
);

BUFx3_ASAP7_75t_L g1939 ( 
.A(n_1428),
.Y(n_1939)
);

INVx5_ASAP7_75t_L g1940 ( 
.A(n_1357),
.Y(n_1940)
);

INVx5_ASAP7_75t_L g1941 ( 
.A(n_1357),
.Y(n_1941)
);

INVx4_ASAP7_75t_L g1942 ( 
.A(n_1501),
.Y(n_1942)
);

INVx3_ASAP7_75t_L g1943 ( 
.A(n_1511),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1431),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1603),
.B(n_1010),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1432),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1484),
.B(n_922),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1506),
.Y(n_1948)
);

CKINVDCx6p67_ASAP7_75t_R g1949 ( 
.A(n_1620),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1633),
.B(n_1010),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1433),
.Y(n_1951)
);

BUFx2_ASAP7_75t_L g1952 ( 
.A(n_1506),
.Y(n_1952)
);

BUFx3_ASAP7_75t_L g1953 ( 
.A(n_1435),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1510),
.B(n_923),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1436),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1437),
.B(n_924),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1510),
.B(n_925),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1441),
.Y(n_1958)
);

BUFx6f_ASAP7_75t_L g1959 ( 
.A(n_1444),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1513),
.B(n_928),
.Y(n_1960)
);

BUFx12f_ASAP7_75t_L g1961 ( 
.A(n_1513),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1447),
.B(n_929),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1520),
.B(n_932),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_1520),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1448),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1449),
.B(n_933),
.Y(n_1966)
);

INVxp67_ASAP7_75t_L g1967 ( 
.A(n_1647),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1450),
.Y(n_1968)
);

XNOR2x1_ASAP7_75t_L g1969 ( 
.A(n_1390),
.B(n_934),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1555),
.B(n_936),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1555),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_SL g1972 ( 
.A(n_1282),
.B(n_1232),
.Y(n_1972)
);

NOR2x1_ASAP7_75t_L g1973 ( 
.A(n_1451),
.B(n_1020),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1452),
.B(n_939),
.Y(n_1974)
);

BUFx6f_ASAP7_75t_L g1975 ( 
.A(n_1454),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1324),
.B(n_1237),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1456),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1669),
.B(n_1020),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1575),
.Y(n_1979)
);

INVxp33_ASAP7_75t_SL g1980 ( 
.A(n_1575),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1457),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_1463),
.Y(n_1982)
);

AND2x6_ASAP7_75t_L g1983 ( 
.A(n_1279),
.B(n_1023),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1464),
.B(n_944),
.Y(n_1984)
);

BUFx6f_ASAP7_75t_L g1985 ( 
.A(n_1465),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1580),
.B(n_946),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1466),
.B(n_950),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1468),
.Y(n_1988)
);

BUFx6f_ASAP7_75t_L g1989 ( 
.A(n_1470),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1473),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1474),
.B(n_951),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1302),
.Y(n_1992)
);

BUFx6f_ASAP7_75t_L g1993 ( 
.A(n_1511),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1522),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1675),
.B(n_952),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1580),
.Y(n_1996)
);

BUFx8_ASAP7_75t_SL g1997 ( 
.A(n_1273),
.Y(n_1997)
);

HB1xp67_ASAP7_75t_L g1998 ( 
.A(n_1614),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1239),
.B(n_1247),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1614),
.B(n_953),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1534),
.B(n_955),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1302),
.Y(n_2002)
);

BUFx12f_ASAP7_75t_L g2003 ( 
.A(n_1618),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1522),
.Y(n_2004)
);

INVx3_ASAP7_75t_L g2005 ( 
.A(n_1538),
.Y(n_2005)
);

INVx5_ASAP7_75t_L g2006 ( 
.A(n_1538),
.Y(n_2006)
);

AND2x4_ASAP7_75t_L g2007 ( 
.A(n_1338),
.B(n_1023),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1241),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1244),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1245),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1246),
.B(n_956),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1618),
.B(n_962),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1648),
.B(n_964),
.Y(n_2013)
);

INVxp33_ASAP7_75t_SL g2014 ( 
.A(n_1648),
.Y(n_2014)
);

BUFx6f_ASAP7_75t_L g2015 ( 
.A(n_1548),
.Y(n_2015)
);

BUFx6f_ASAP7_75t_L g2016 ( 
.A(n_1548),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_L g2017 ( 
.A(n_1534),
.B(n_968),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1650),
.B(n_970),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1248),
.B(n_971),
.Y(n_2019)
);

BUFx6f_ASAP7_75t_L g2020 ( 
.A(n_1600),
.Y(n_2020)
);

INVx4_ASAP7_75t_L g2021 ( 
.A(n_1650),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1581),
.B(n_972),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1321),
.Y(n_2023)
);

BUFx6f_ASAP7_75t_L g2024 ( 
.A(n_1600),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1581),
.B(n_973),
.Y(n_2025)
);

AND2x6_ASAP7_75t_L g2026 ( 
.A(n_1250),
.B(n_1026),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1322),
.Y(n_2027)
);

BUFx6f_ASAP7_75t_L g2028 ( 
.A(n_1673),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1323),
.Y(n_2029)
);

INVx5_ASAP7_75t_L g2030 ( 
.A(n_1673),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1254),
.B(n_974),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1255),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1256),
.B(n_976),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1651),
.B(n_978),
.Y(n_2034)
);

BUFx6f_ASAP7_75t_L g2035 ( 
.A(n_1260),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1261),
.B(n_980),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1326),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1651),
.B(n_981),
.Y(n_2038)
);

AND3x2_ASAP7_75t_L g2039 ( 
.A(n_1684),
.B(n_1913),
.C(n_1866),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2023),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1720),
.Y(n_2041)
);

INVx3_ASAP7_75t_L g2042 ( 
.A(n_1725),
.Y(n_2042)
);

BUFx6f_ASAP7_75t_L g2043 ( 
.A(n_1725),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2027),
.Y(n_2044)
);

OA21x2_ASAP7_75t_L g2045 ( 
.A1(n_1881),
.A2(n_1903),
.B(n_1893),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2029),
.Y(n_2046)
);

HB1xp67_ASAP7_75t_L g2047 ( 
.A(n_1708),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2037),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1939),
.Y(n_2049)
);

OA21x2_ASAP7_75t_L g2050 ( 
.A1(n_1909),
.A2(n_1265),
.B(n_1264),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1708),
.B(n_1652),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1720),
.Y(n_2052)
);

BUFx3_ASAP7_75t_L g2053 ( 
.A(n_1912),
.Y(n_2053)
);

OA21x2_ASAP7_75t_L g2054 ( 
.A1(n_1918),
.A2(n_1268),
.B(n_1267),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1939),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_1725),
.Y(n_2056)
);

OR2x6_ASAP7_75t_L g2057 ( 
.A(n_1718),
.B(n_1387),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1944),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1944),
.Y(n_2059)
);

BUFx6f_ASAP7_75t_L g2060 ( 
.A(n_1725),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1704),
.B(n_1270),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1713),
.B(n_1271),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_1718),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1953),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1953),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1747),
.B(n_1272),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1982),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1773),
.B(n_1281),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1721),
.Y(n_2069)
);

AOI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_1684),
.A2(n_1768),
.B1(n_1811),
.B2(n_1792),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1765),
.B(n_1284),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1726),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1721),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1982),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_1748),
.B(n_1519),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1707),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1748),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1707),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1712),
.Y(n_2079)
);

OAI22xp5_ASAP7_75t_SL g2080 ( 
.A1(n_1861),
.A2(n_1193),
.B1(n_1366),
.B2(n_1306),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1712),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1758),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_1726),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1740),
.B(n_1652),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_L g2085 ( 
.A(n_1915),
.B(n_1672),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1726),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1758),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1915),
.B(n_1286),
.Y(n_2088)
);

INVxp33_ASAP7_75t_SL g2089 ( 
.A(n_1798),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1686),
.B(n_1654),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_1912),
.B(n_1476),
.Y(n_2091)
);

AOI22xp5_ASAP7_75t_SL g2092 ( 
.A1(n_1789),
.A2(n_1306),
.B1(n_1372),
.B2(n_1366),
.Y(n_2092)
);

BUFx3_ASAP7_75t_L g2093 ( 
.A(n_1697),
.Y(n_2093)
);

INVx3_ASAP7_75t_L g2094 ( 
.A(n_1726),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1817),
.Y(n_2095)
);

BUFx6f_ASAP7_75t_L g2096 ( 
.A(n_1738),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1967),
.B(n_1287),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1817),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1750),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_1738),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1837),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_L g2102 ( 
.A(n_1738),
.Y(n_2102)
);

INVx3_ASAP7_75t_L g2103 ( 
.A(n_1738),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1967),
.B(n_1920),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1750),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1837),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1858),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1858),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1686),
.B(n_1654),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_1767),
.Y(n_2110)
);

NOR2x1_ASAP7_75t_L g2111 ( 
.A(n_1867),
.B(n_1328),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1786),
.B(n_1288),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1863),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1775),
.Y(n_2114)
);

AOI22xp5_ASAP7_75t_L g2115 ( 
.A1(n_1768),
.A2(n_1636),
.B1(n_1656),
.B2(n_1630),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1892),
.B(n_1668),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1863),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1864),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1864),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1872),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1872),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_1698),
.B(n_1668),
.Y(n_2122)
);

INVx4_ASAP7_75t_L g2123 ( 
.A(n_1702),
.Y(n_2123)
);

BUFx3_ASAP7_75t_L g2124 ( 
.A(n_1697),
.Y(n_2124)
);

INVx3_ASAP7_75t_L g2125 ( 
.A(n_1767),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2008),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2008),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1775),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1793),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1892),
.B(n_1887),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1793),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1829),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2009),
.Y(n_2133)
);

INVxp67_ASAP7_75t_L g2134 ( 
.A(n_1709),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_1792),
.A2(n_1636),
.B1(n_1656),
.B2(n_1630),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2009),
.Y(n_2136)
);

BUFx6f_ASAP7_75t_L g2137 ( 
.A(n_1767),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_1698),
.B(n_1678),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_SL g2139 ( 
.A(n_1887),
.B(n_1678),
.Y(n_2139)
);

BUFx3_ASAP7_75t_L g2140 ( 
.A(n_1701),
.Y(n_2140)
);

INVx5_ASAP7_75t_L g2141 ( 
.A(n_1714),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2026),
.B(n_2011),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2010),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1829),
.Y(n_2144)
);

BUFx2_ASAP7_75t_L g2145 ( 
.A(n_1724),
.Y(n_2145)
);

BUFx6f_ASAP7_75t_L g2146 ( 
.A(n_1767),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2026),
.B(n_1290),
.Y(n_2147)
);

HB1xp67_ASAP7_75t_L g2148 ( 
.A(n_1761),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1830),
.Y(n_2149)
);

BUFx8_ASAP7_75t_L g2150 ( 
.A(n_1779),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2010),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_1772),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2032),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1821),
.B(n_1627),
.Y(n_2154)
);

NOR2xp33_ASAP7_75t_L g2155 ( 
.A(n_1995),
.B(n_1672),
.Y(n_2155)
);

HB1xp67_ASAP7_75t_L g2156 ( 
.A(n_1761),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2032),
.Y(n_2157)
);

NOR2xp33_ASAP7_75t_L g2158 ( 
.A(n_2019),
.B(n_1324),
.Y(n_2158)
);

AND2x4_ASAP7_75t_SL g2159 ( 
.A(n_1769),
.B(n_1372),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_1701),
.B(n_1477),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_2031),
.B(n_1263),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2035),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1830),
.Y(n_2163)
);

HB1xp67_ASAP7_75t_L g2164 ( 
.A(n_1763),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1842),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1842),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2035),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2026),
.B(n_1291),
.Y(n_2168)
);

INVxp67_ASAP7_75t_L g2169 ( 
.A(n_1709),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_1734),
.B(n_1480),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1860),
.Y(n_2171)
);

OA21x2_ASAP7_75t_L g2172 ( 
.A1(n_1999),
.A2(n_1295),
.B(n_1292),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_1700),
.B(n_1642),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1860),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2026),
.B(n_1296),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1871),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_1772),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_1772),
.Y(n_2178)
);

AND2x6_ASAP7_75t_L g2179 ( 
.A(n_1691),
.B(n_1298),
.Y(n_2179)
);

INVx3_ASAP7_75t_L g2180 ( 
.A(n_1772),
.Y(n_2180)
);

BUFx2_ASAP7_75t_L g2181 ( 
.A(n_1724),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2035),
.Y(n_2182)
);

CKINVDCx8_ASAP7_75t_R g2183 ( 
.A(n_1731),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2035),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1781),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1871),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_SL g2187 ( 
.A(n_1980),
.B(n_1655),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_1722),
.B(n_1657),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1790),
.Y(n_2189)
);

INVx3_ASAP7_75t_L g2190 ( 
.A(n_1782),
.Y(n_2190)
);

AND2x4_ASAP7_75t_L g2191 ( 
.A(n_1734),
.B(n_1481),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1810),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1782),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1812),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_2033),
.B(n_1263),
.Y(n_2195)
);

INVxp67_ASAP7_75t_L g2196 ( 
.A(n_1808),
.Y(n_2196)
);

AND2x2_ASAP7_75t_SL g2197 ( 
.A(n_1839),
.B(n_1026),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1859),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1911),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1992),
.Y(n_2200)
);

INVx1_ASAP7_75t_SL g2201 ( 
.A(n_1828),
.Y(n_2201)
);

AND2x6_ASAP7_75t_L g2202 ( 
.A(n_1695),
.B(n_1299),
.Y(n_2202)
);

INVx3_ASAP7_75t_L g2203 ( 
.A(n_1782),
.Y(n_2203)
);

BUFx6f_ASAP7_75t_L g2204 ( 
.A(n_1782),
.Y(n_2204)
);

INVx3_ASAP7_75t_L g2205 ( 
.A(n_1788),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_1739),
.B(n_1482),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2026),
.B(n_1300),
.Y(n_2207)
);

AND2x4_ASAP7_75t_L g2208 ( 
.A(n_1739),
.B(n_1485),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1938),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1955),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_1730),
.B(n_1661),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1958),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_1788),
.Y(n_2213)
);

BUFx6f_ASAP7_75t_L g2214 ( 
.A(n_1788),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1965),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1992),
.Y(n_2216)
);

OA21x2_ASAP7_75t_L g2217 ( 
.A1(n_2036),
.A2(n_1304),
.B(n_1301),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_1732),
.B(n_1327),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1968),
.Y(n_2219)
);

BUFx8_ASAP7_75t_L g2220 ( 
.A(n_1779),
.Y(n_2220)
);

BUFx6f_ASAP7_75t_L g2221 ( 
.A(n_1788),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1680),
.B(n_1307),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1682),
.B(n_1314),
.Y(n_2223)
);

INVx3_ASAP7_75t_L g2224 ( 
.A(n_1801),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1977),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1801),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1833),
.B(n_1327),
.Y(n_2227)
);

INVxp67_ASAP7_75t_L g2228 ( 
.A(n_1934),
.Y(n_2228)
);

NOR2xp33_ASAP7_75t_L g2229 ( 
.A(n_1755),
.B(n_1362),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1801),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_1801),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_1737),
.B(n_1362),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_SL g2233 ( 
.A(n_1751),
.B(n_1315),
.Y(n_2233)
);

AND2x2_ASAP7_75t_SL g2234 ( 
.A(n_1839),
.B(n_1041),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1802),
.Y(n_2235)
);

AOI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_1811),
.A2(n_1638),
.B1(n_1634),
.B2(n_1165),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1802),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1802),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2002),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1802),
.Y(n_2240)
);

BUFx3_ASAP7_75t_L g2241 ( 
.A(n_1751),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_1710),
.B(n_1368),
.Y(n_2242)
);

HB1xp67_ASAP7_75t_L g2243 ( 
.A(n_1763),
.Y(n_2243)
);

OAI22xp5_ASAP7_75t_SL g2244 ( 
.A1(n_1692),
.A2(n_1385),
.B1(n_1443),
.B2(n_1426),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_1696),
.B(n_1711),
.Y(n_2245)
);

BUFx8_ASAP7_75t_L g2246 ( 
.A(n_1754),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1804),
.Y(n_2247)
);

XNOR2x2_ASAP7_75t_R g2248 ( 
.A(n_1794),
.B(n_1385),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2002),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_1723),
.B(n_1733),
.Y(n_2250)
);

OA21x2_ASAP7_75t_L g2251 ( 
.A1(n_1930),
.A2(n_1317),
.B(n_1316),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_1742),
.B(n_1330),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1804),
.Y(n_2253)
);

AND2x4_ASAP7_75t_L g2254 ( 
.A(n_1753),
.B(n_1486),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_L g2255 ( 
.A(n_1755),
.B(n_1368),
.Y(n_2255)
);

BUFx6f_ASAP7_75t_L g2256 ( 
.A(n_1804),
.Y(n_2256)
);

INVx6_ASAP7_75t_L g2257 ( 
.A(n_1702),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1804),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1879),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1805),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1805),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_1753),
.B(n_1332),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1805),
.Y(n_2263)
);

INVx5_ASAP7_75t_L g2264 ( 
.A(n_1714),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1805),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1807),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_1741),
.B(n_1371),
.Y(n_2267)
);

AND2x4_ASAP7_75t_L g2268 ( 
.A(n_1945),
.B(n_1487),
.Y(n_2268)
);

BUFx6f_ASAP7_75t_L g2269 ( 
.A(n_1807),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1807),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1756),
.B(n_1333),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1807),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1809),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_1727),
.B(n_1334),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1809),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1727),
.B(n_1335),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1879),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1809),
.Y(n_2278)
);

BUFx6f_ASAP7_75t_L g2279 ( 
.A(n_1809),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1816),
.Y(n_2280)
);

INVx6_ASAP7_75t_L g2281 ( 
.A(n_1741),
.Y(n_2281)
);

INVx3_ASAP7_75t_L g2282 ( 
.A(n_1816),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1816),
.Y(n_2283)
);

CKINVDCx5p33_ASAP7_75t_R g2284 ( 
.A(n_1828),
.Y(n_2284)
);

INVx5_ASAP7_75t_L g2285 ( 
.A(n_1714),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1816),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1841),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_1886),
.Y(n_2288)
);

BUFx6f_ASAP7_75t_L g2289 ( 
.A(n_1841),
.Y(n_2289)
);

OR2x6_ASAP7_75t_L g2290 ( 
.A(n_1745),
.B(n_1423),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1841),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1841),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1852),
.Y(n_2293)
);

OA21x2_ASAP7_75t_L g2294 ( 
.A1(n_1932),
.A2(n_1337),
.B(n_1336),
.Y(n_2294)
);

BUFx6f_ASAP7_75t_L g2295 ( 
.A(n_1852),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1886),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1890),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_1890),
.Y(n_2298)
);

BUFx3_ASAP7_75t_L g2299 ( 
.A(n_1852),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_1852),
.Y(n_2300)
);

CKINVDCx5p33_ASAP7_75t_R g2301 ( 
.A(n_1935),
.Y(n_2301)
);

CKINVDCx6p67_ASAP7_75t_R g2302 ( 
.A(n_1949),
.Y(n_2302)
);

INVx3_ASAP7_75t_L g2303 ( 
.A(n_1857),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_1945),
.B(n_1490),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_1897),
.Y(n_2305)
);

INVx3_ASAP7_75t_L g2306 ( 
.A(n_1857),
.Y(n_2306)
);

OR2x6_ASAP7_75t_L g2307 ( 
.A(n_1752),
.B(n_1693),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1897),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1857),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1729),
.B(n_1340),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1857),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_L g2312 ( 
.A(n_1710),
.B(n_1371),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_1910),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_1862),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1862),
.Y(n_2315)
);

INVx3_ASAP7_75t_L g2316 ( 
.A(n_1862),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_1729),
.B(n_1342),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1862),
.Y(n_2318)
);

BUFx6f_ASAP7_75t_L g2319 ( 
.A(n_1681),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_1744),
.B(n_1344),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_1843),
.B(n_1380),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_1910),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1683),
.B(n_1345),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_1924),
.Y(n_2324)
);

OAI21x1_ASAP7_75t_L g2325 ( 
.A1(n_1956),
.A2(n_1347),
.B(n_1346),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1878),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_1924),
.Y(n_2327)
);

BUFx6f_ASAP7_75t_L g2328 ( 
.A(n_1681),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1878),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_1855),
.B(n_1380),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_L g2331 ( 
.A(n_1820),
.B(n_1445),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_1681),
.Y(n_2332)
);

BUFx6f_ASAP7_75t_L g2333 ( 
.A(n_1681),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1878),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1878),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1900),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_1900),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1900),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_1926),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_1683),
.B(n_1348),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_1900),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1905),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_1685),
.B(n_1349),
.Y(n_2343)
);

AND2x4_ASAP7_75t_L g2344 ( 
.A(n_1950),
.B(n_1491),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_1926),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_1935),
.Y(n_2346)
);

BUFx6f_ASAP7_75t_L g2347 ( 
.A(n_1687),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1905),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1905),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1685),
.B(n_1352),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_1905),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_SL g2352 ( 
.A(n_1868),
.B(n_986),
.Y(n_2352)
);

HB1xp67_ASAP7_75t_L g2353 ( 
.A(n_1764),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_1931),
.Y(n_2354)
);

INVx3_ASAP7_75t_L g2355 ( 
.A(n_1687),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1931),
.Y(n_2356)
);

AND2x4_ASAP7_75t_L g2357 ( 
.A(n_1950),
.B(n_1492),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1931),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1931),
.Y(n_2359)
);

INVx3_ASAP7_75t_L g2360 ( 
.A(n_1687),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_1946),
.Y(n_2361)
);

AND2x6_ASAP7_75t_L g2362 ( 
.A(n_1774),
.B(n_1041),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_1990),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_1946),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_1946),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_SL g2366 ( 
.A(n_2014),
.B(n_1033),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_1823),
.B(n_1496),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_1946),
.Y(n_2368)
);

HB1xp67_ASAP7_75t_L g2369 ( 
.A(n_1764),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1951),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1951),
.Y(n_2371)
);

BUFx6f_ASAP7_75t_L g2372 ( 
.A(n_1687),
.Y(n_2372)
);

INVxp67_ASAP7_75t_L g2373 ( 
.A(n_1706),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1951),
.Y(n_2374)
);

BUFx6f_ASAP7_75t_L g2375 ( 
.A(n_1688),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1951),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_SL g2377 ( 
.A(n_1876),
.B(n_988),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_1959),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_1688),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_1990),
.Y(n_2380)
);

AND3x2_ASAP7_75t_L g2381 ( 
.A(n_1929),
.B(n_1045),
.C(n_1043),
.Y(n_2381)
);

BUFx2_ASAP7_75t_L g2382 ( 
.A(n_1969),
.Y(n_2382)
);

BUFx2_ASAP7_75t_L g2383 ( 
.A(n_1716),
.Y(n_2383)
);

AND2x4_ASAP7_75t_L g2384 ( 
.A(n_1978),
.B(n_1497),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_1826),
.B(n_1499),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_1834),
.B(n_1500),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_1978),
.B(n_1502),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1959),
.Y(n_2388)
);

HB1xp67_ASAP7_75t_L g2389 ( 
.A(n_1771),
.Y(n_2389)
);

INVxp67_ASAP7_75t_L g2390 ( 
.A(n_1706),
.Y(n_2390)
);

BUFx6f_ASAP7_75t_L g2391 ( 
.A(n_1688),
.Y(n_2391)
);

HB1xp67_ASAP7_75t_L g2392 ( 
.A(n_1771),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_1993),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1959),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1959),
.Y(n_2395)
);

AND2x4_ASAP7_75t_L g2396 ( 
.A(n_1882),
.B(n_1504),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_L g2397 ( 
.A(n_1688),
.Y(n_2397)
);

INVx3_ASAP7_75t_L g2398 ( 
.A(n_1689),
.Y(n_2398)
);

INVx3_ASAP7_75t_L g2399 ( 
.A(n_1689),
.Y(n_2399)
);

BUFx6f_ASAP7_75t_L g2400 ( 
.A(n_1689),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_1993),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_1993),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_1993),
.Y(n_2403)
);

AND2x6_ASAP7_75t_L g2404 ( 
.A(n_1880),
.B(n_1043),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_1994),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_1994),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_1994),
.Y(n_2407)
);

INVx3_ASAP7_75t_L g2408 ( 
.A(n_1689),
.Y(n_2408)
);

XOR2xp5_ASAP7_75t_L g2409 ( 
.A(n_1692),
.B(n_1426),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_1994),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_1975),
.Y(n_2411)
);

BUFx6f_ASAP7_75t_L g2412 ( 
.A(n_1690),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2015),
.Y(n_2413)
);

BUFx2_ASAP7_75t_L g2414 ( 
.A(n_1746),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_1975),
.Y(n_2415)
);

AND3x1_ASAP7_75t_L g2416 ( 
.A(n_1820),
.B(n_1055),
.C(n_1045),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2015),
.Y(n_2417)
);

AND2x4_ASAP7_75t_L g2418 ( 
.A(n_1882),
.B(n_1507),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_1791),
.B(n_1851),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1975),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_1975),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2015),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_1981),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2015),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2016),
.Y(n_2425)
);

INVx5_ASAP7_75t_L g2426 ( 
.A(n_1714),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_1981),
.Y(n_2427)
);

CKINVDCx20_ASAP7_75t_R g2428 ( 
.A(n_1997),
.Y(n_2428)
);

AND2x4_ASAP7_75t_L g2429 ( 
.A(n_1791),
.B(n_1508),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2016),
.B(n_1509),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_1981),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_1981),
.Y(n_2432)
);

BUFx6f_ASAP7_75t_L g2433 ( 
.A(n_1690),
.Y(n_2433)
);

NOR2xp33_ASAP7_75t_L g2434 ( 
.A(n_1835),
.B(n_1445),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_SL g2435 ( 
.A(n_1902),
.B(n_1904),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2016),
.B(n_1514),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_1985),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2016),
.Y(n_2438)
);

NOR2xp33_ASAP7_75t_L g2439 ( 
.A(n_1835),
.B(n_1493),
.Y(n_2439)
);

INVx3_ASAP7_75t_L g2440 ( 
.A(n_1690),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_1985),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_1848),
.B(n_1493),
.Y(n_2442)
);

BUFx6f_ASAP7_75t_L g2443 ( 
.A(n_1690),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_1985),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_1985),
.Y(n_2445)
);

INVxp67_ASAP7_75t_L g2446 ( 
.A(n_1848),
.Y(n_2446)
);

HB1xp67_ASAP7_75t_L g2447 ( 
.A(n_1827),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_1988),
.Y(n_2448)
);

INVx5_ASAP7_75t_L g2449 ( 
.A(n_1714),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2020),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_1988),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2020),
.Y(n_2452)
);

NOR2xp33_ASAP7_75t_L g2453 ( 
.A(n_1884),
.B(n_1503),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2020),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2259),
.Y(n_2455)
);

OR2x6_ASAP7_75t_L g2456 ( 
.A(n_2307),
.B(n_1815),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2148),
.Y(n_2457)
);

BUFx2_ASAP7_75t_L g2458 ( 
.A(n_2047),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2200),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2200),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2232),
.B(n_1822),
.Y(n_2461)
);

INVx5_ASAP7_75t_L g2462 ( 
.A(n_2141),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2216),
.Y(n_2463)
);

INVx3_ASAP7_75t_L g2464 ( 
.A(n_2216),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2239),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2239),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2249),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2218),
.B(n_1822),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2259),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2330),
.B(n_1869),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2277),
.Y(n_2471)
);

BUFx2_ASAP7_75t_L g2472 ( 
.A(n_2047),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2277),
.Y(n_2473)
);

AOI22x1_ASAP7_75t_L g2474 ( 
.A1(n_2373),
.A2(n_1916),
.B1(n_1954),
.B2(n_1908),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2288),
.Y(n_2475)
);

INVx3_ASAP7_75t_L g2476 ( 
.A(n_2249),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2321),
.B(n_1869),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2104),
.B(n_1884),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_L g2479 ( 
.A(n_2197),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2041),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2245),
.B(n_1888),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2041),
.Y(n_2482)
);

INVx2_ASAP7_75t_SL g2483 ( 
.A(n_2241),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2250),
.B(n_1888),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2148),
.Y(n_2485)
);

INVx3_ASAP7_75t_L g2486 ( 
.A(n_2052),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2052),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2197),
.B(n_1927),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2156),
.Y(n_2489)
);

OR2x2_ASAP7_75t_L g2490 ( 
.A(n_2075),
.B(n_1797),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_SL g2491 ( 
.A(n_2070),
.B(n_1743),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2156),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2164),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2164),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2243),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2243),
.Y(n_2496)
);

AND2x4_ASAP7_75t_L g2497 ( 
.A(n_2241),
.B(n_1922),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2234),
.B(n_1927),
.Y(n_2498)
);

NAND2xp33_ASAP7_75t_L g2499 ( 
.A(n_2404),
.B(n_1749),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2288),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_2227),
.B(n_2021),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2353),
.Y(n_2502)
);

AND2x2_ASAP7_75t_SL g2503 ( 
.A(n_2234),
.B(n_1789),
.Y(n_2503)
);

BUFx6f_ASAP7_75t_L g2504 ( 
.A(n_2043),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_SL g2505 ( 
.A(n_2331),
.B(n_2021),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_SL g2506 ( 
.A(n_2331),
.B(n_1867),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2242),
.B(n_1957),
.Y(n_2507)
);

AND3x1_ASAP7_75t_L g2508 ( 
.A(n_2366),
.B(n_1947),
.C(n_1936),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_L g2509 ( 
.A(n_2446),
.B(n_1971),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2069),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2069),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2353),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2369),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2073),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2369),
.Y(n_2515)
);

INVx5_ASAP7_75t_L g2516 ( 
.A(n_2141),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2073),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2389),
.Y(n_2518)
);

CKINVDCx5p33_ASAP7_75t_R g2519 ( 
.A(n_2284),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2389),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2099),
.Y(n_2521)
);

INVx4_ASAP7_75t_L g2522 ( 
.A(n_2141),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2392),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2222),
.B(n_1936),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2099),
.Y(n_2525)
);

BUFx2_ASAP7_75t_L g2526 ( 
.A(n_2063),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2105),
.Y(n_2527)
);

AO21x2_ASAP7_75t_L g2528 ( 
.A1(n_2142),
.A2(n_1818),
.B(n_1799),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2105),
.Y(n_2529)
);

BUFx10_ASAP7_75t_L g2530 ( 
.A(n_2434),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2114),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2114),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2128),
.Y(n_2533)
);

BUFx3_ASAP7_75t_L g2534 ( 
.A(n_2053),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2296),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_L g2536 ( 
.A(n_2446),
.B(n_1996),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2128),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2129),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2129),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2296),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2297),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2131),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2131),
.Y(n_2543)
);

BUFx2_ASAP7_75t_L g2544 ( 
.A(n_2063),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_SL g2545 ( 
.A(n_2434),
.B(n_1894),
.Y(n_2545)
);

NOR2xp33_ASAP7_75t_L g2546 ( 
.A(n_2134),
.B(n_1894),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2132),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2132),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_L g2549 ( 
.A(n_2134),
.B(n_1919),
.Y(n_2549)
);

INVxp67_ASAP7_75t_SL g2550 ( 
.A(n_2043),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_SL g2551 ( 
.A(n_2439),
.B(n_1919),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2144),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2223),
.B(n_1947),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2439),
.B(n_2001),
.Y(n_2554)
);

AND3x2_ASAP7_75t_L g2555 ( 
.A(n_2145),
.B(n_1762),
.C(n_1760),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2442),
.B(n_2001),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2297),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2298),
.Y(n_2558)
);

AND2x6_ASAP7_75t_L g2559 ( 
.A(n_2084),
.B(n_1960),
.Y(n_2559)
);

BUFx6f_ASAP7_75t_SL g2560 ( 
.A(n_2307),
.Y(n_2560)
);

AO21x2_ASAP7_75t_L g2561 ( 
.A1(n_2325),
.A2(n_2168),
.B(n_2147),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_SL g2562 ( 
.A(n_2442),
.B(n_1942),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2453),
.B(n_2071),
.Y(n_2563)
);

INVx2_ASAP7_75t_SL g2564 ( 
.A(n_2130),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_SL g2565 ( 
.A(n_2453),
.B(n_2155),
.Y(n_2565)
);

NAND2xp33_ASAP7_75t_SL g2566 ( 
.A(n_2435),
.B(n_1799),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2392),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_2155),
.B(n_2267),
.Y(n_2568)
);

INVx3_ASAP7_75t_L g2569 ( 
.A(n_2144),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2373),
.B(n_1963),
.Y(n_2570)
);

INVx5_ASAP7_75t_L g2571 ( 
.A(n_2141),
.Y(n_2571)
);

INVx3_ASAP7_75t_L g2572 ( 
.A(n_2149),
.Y(n_2572)
);

INVx3_ASAP7_75t_L g2573 ( 
.A(n_2149),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2252),
.B(n_2017),
.Y(n_2574)
);

BUFx6f_ASAP7_75t_L g2575 ( 
.A(n_2043),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2040),
.Y(n_2576)
);

OR2x6_ASAP7_75t_L g2577 ( 
.A(n_2307),
.B(n_1815),
.Y(n_2577)
);

INVx3_ASAP7_75t_L g2578 ( 
.A(n_2163),
.Y(n_2578)
);

INVx3_ASAP7_75t_L g2579 ( 
.A(n_2163),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2044),
.Y(n_2580)
);

BUFx4f_ASAP7_75t_L g2581 ( 
.A(n_2404),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2046),
.Y(n_2582)
);

INVx4_ASAP7_75t_L g2583 ( 
.A(n_2264),
.Y(n_2583)
);

HB1xp67_ASAP7_75t_L g2584 ( 
.A(n_2077),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2271),
.B(n_2112),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2165),
.Y(n_2586)
);

NAND2xp33_ASAP7_75t_SL g2587 ( 
.A(n_2435),
.B(n_1818),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2165),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_SL g2589 ( 
.A(n_2267),
.B(n_1942),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2166),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2048),
.Y(n_2591)
);

INVx8_ASAP7_75t_L g2592 ( 
.A(n_2179),
.Y(n_2592)
);

BUFx6f_ASAP7_75t_L g2593 ( 
.A(n_2043),
.Y(n_2593)
);

CKINVDCx11_ASAP7_75t_R g2594 ( 
.A(n_2428),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2091),
.Y(n_2595)
);

BUFx6f_ASAP7_75t_L g2596 ( 
.A(n_2060),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2166),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2171),
.Y(n_2598)
);

NOR3xp33_ASAP7_75t_L g2599 ( 
.A(n_2090),
.B(n_1840),
.C(n_1972),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2171),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_SL g2601 ( 
.A(n_2085),
.B(n_1891),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2174),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2091),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2161),
.B(n_2195),
.Y(n_2604)
);

BUFx10_ASAP7_75t_L g2605 ( 
.A(n_2312),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_SL g2606 ( 
.A(n_2085),
.B(n_1840),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2174),
.Y(n_2607)
);

INVx3_ASAP7_75t_L g2608 ( 
.A(n_2176),
.Y(n_2608)
);

INVx2_ASAP7_75t_SL g2609 ( 
.A(n_2077),
.Y(n_2609)
);

INVx4_ASAP7_75t_L g2610 ( 
.A(n_2264),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2049),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2055),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2176),
.Y(n_2613)
);

AND2x4_ASAP7_75t_L g2614 ( 
.A(n_2053),
.B(n_1922),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2058),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2186),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_L g2617 ( 
.A(n_2169),
.B(n_2017),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2390),
.B(n_1970),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2186),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2059),
.Y(n_2620)
);

INVx1_ASAP7_75t_SL g2621 ( 
.A(n_2051),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2298),
.Y(n_2622)
);

INVx1_ASAP7_75t_SL g2623 ( 
.A(n_2383),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2305),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_SL g2625 ( 
.A(n_2158),
.B(n_1703),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2390),
.B(n_2312),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2161),
.B(n_2022),
.Y(n_2627)
);

BUFx6f_ASAP7_75t_L g2628 ( 
.A(n_2060),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2305),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2308),
.Y(n_2630)
);

INVxp67_ASAP7_75t_SL g2631 ( 
.A(n_2060),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2308),
.Y(n_2632)
);

BUFx10_ASAP7_75t_L g2633 ( 
.A(n_2229),
.Y(n_2633)
);

AOI21x1_ASAP7_75t_L g2634 ( 
.A1(n_2126),
.A2(n_1966),
.B(n_1962),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2195),
.B(n_2022),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2088),
.B(n_2025),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2313),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2313),
.Y(n_2638)
);

NOR2xp33_ASAP7_75t_L g2639 ( 
.A(n_2169),
.B(n_2025),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_SL g2640 ( 
.A(n_2158),
.B(n_1703),
.Y(n_2640)
);

INVx2_ASAP7_75t_SL g2641 ( 
.A(n_2160),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2064),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2322),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2322),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2065),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2324),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_SL g2647 ( 
.A(n_2116),
.B(n_2154),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2067),
.Y(n_2648)
);

NAND3xp33_ASAP7_75t_L g2649 ( 
.A(n_2229),
.B(n_2255),
.C(n_2447),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2324),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2327),
.Y(n_2651)
);

BUFx3_ASAP7_75t_L g2652 ( 
.A(n_2093),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_SL g2653 ( 
.A(n_2255),
.B(n_1705),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_2301),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2074),
.Y(n_2655)
);

INVx3_ASAP7_75t_L g2656 ( 
.A(n_2172),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2323),
.Y(n_2657)
);

CKINVDCx6p67_ASAP7_75t_R g2658 ( 
.A(n_2302),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_SL g2659 ( 
.A(n_2344),
.B(n_2357),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2340),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2327),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2343),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2339),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2339),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2345),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2345),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2097),
.B(n_2038),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2363),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2363),
.Y(n_2669)
);

INVx3_ASAP7_75t_L g2670 ( 
.A(n_2172),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2380),
.Y(n_2671)
);

INVx4_ASAP7_75t_L g2672 ( 
.A(n_2264),
.Y(n_2672)
);

INVx2_ASAP7_75t_SL g2673 ( 
.A(n_2160),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2380),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2127),
.Y(n_2675)
);

INVx3_ASAP7_75t_L g2676 ( 
.A(n_2172),
.Y(n_2676)
);

BUFx6f_ASAP7_75t_L g2677 ( 
.A(n_2060),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2133),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2136),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2143),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_SL g2681 ( 
.A(n_2344),
.B(n_1705),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_L g2682 ( 
.A(n_2090),
.B(n_1824),
.Y(n_2682)
);

AND2x4_ASAP7_75t_L g2683 ( 
.A(n_2093),
.B(n_1923),
.Y(n_2683)
);

AND2x6_ASAP7_75t_L g2684 ( 
.A(n_2111),
.B(n_1986),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2151),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2153),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2157),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2393),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2061),
.B(n_2000),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_SL g2690 ( 
.A(n_2357),
.B(n_1778),
.Y(n_2690)
);

BUFx6f_ASAP7_75t_L g2691 ( 
.A(n_2072),
.Y(n_2691)
);

INVx3_ASAP7_75t_L g2692 ( 
.A(n_2393),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_2346),
.Y(n_2693)
);

HB1xp67_ASAP7_75t_L g2694 ( 
.A(n_2057),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2350),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2401),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2430),
.Y(n_2697)
);

INVx2_ASAP7_75t_SL g2698 ( 
.A(n_2294),
.Y(n_2698)
);

NOR2x1p5_ASAP7_75t_L g2699 ( 
.A(n_2173),
.B(n_1787),
.Y(n_2699)
);

INVxp33_ASAP7_75t_L g2700 ( 
.A(n_2244),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2185),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2401),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2062),
.B(n_2066),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2402),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_SL g2705 ( 
.A(n_2384),
.B(n_1784),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2402),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2403),
.Y(n_2707)
);

INVx8_ASAP7_75t_L g2708 ( 
.A(n_2179),
.Y(n_2708)
);

INVxp33_ASAP7_75t_L g2709 ( 
.A(n_2447),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2068),
.B(n_2012),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2320),
.B(n_2013),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2189),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_SL g2713 ( 
.A(n_2384),
.B(n_1800),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2192),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2194),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2403),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2198),
.Y(n_2717)
);

INVx4_ASAP7_75t_L g2718 ( 
.A(n_2264),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_SL g2719 ( 
.A(n_2387),
.B(n_1813),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2367),
.B(n_2018),
.Y(n_2720)
);

INVx8_ASAP7_75t_L g2721 ( 
.A(n_2179),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2385),
.B(n_2034),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2199),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2405),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2209),
.Y(n_2725)
);

OR2x6_ASAP7_75t_L g2726 ( 
.A(n_2123),
.B(n_1846),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2210),
.Y(n_2727)
);

INVx4_ASAP7_75t_L g2728 ( 
.A(n_2285),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2405),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2436),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2406),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2406),
.Y(n_2732)
);

INVx2_ASAP7_75t_SL g2733 ( 
.A(n_2294),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2212),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2215),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2219),
.Y(n_2736)
);

OR2x2_ASAP7_75t_L g2737 ( 
.A(n_2057),
.B(n_1972),
.Y(n_2737)
);

INVx3_ASAP7_75t_L g2738 ( 
.A(n_2407),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2225),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_SL g2740 ( 
.A(n_2387),
.B(n_1814),
.Y(n_2740)
);

INVx8_ASAP7_75t_L g2741 ( 
.A(n_2179),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2268),
.B(n_2007),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2407),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2410),
.Y(n_2744)
);

AND2x2_ASAP7_75t_L g2745 ( 
.A(n_2268),
.B(n_2007),
.Y(n_2745)
);

AOI21x1_ASAP7_75t_L g2746 ( 
.A1(n_2175),
.A2(n_1984),
.B(n_1974),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2386),
.B(n_1854),
.Y(n_2747)
);

INVx3_ASAP7_75t_L g2748 ( 
.A(n_2410),
.Y(n_2748)
);

AND3x2_ASAP7_75t_L g2749 ( 
.A(n_2181),
.B(n_1899),
.C(n_1873),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2404),
.B(n_1854),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_SL g2751 ( 
.A(n_2419),
.B(n_1952),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2101),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2106),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2413),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2107),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2413),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2108),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2417),
.Y(n_2758)
);

AOI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2404),
.A2(n_2362),
.B1(n_2122),
.B2(n_2138),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_SL g2760 ( 
.A(n_2419),
.B(n_1883),
.Y(n_2760)
);

INVxp67_ASAP7_75t_SL g2761 ( 
.A(n_2072),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2417),
.Y(n_2762)
);

OR2x6_ASAP7_75t_L g2763 ( 
.A(n_2123),
.B(n_1846),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2113),
.Y(n_2764)
);

AND2x2_ASAP7_75t_L g2765 ( 
.A(n_2304),
.B(n_1923),
.Y(n_2765)
);

BUFx2_ASAP7_75t_L g2766 ( 
.A(n_2057),
.Y(n_2766)
);

INVx2_ASAP7_75t_SL g2767 ( 
.A(n_2294),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2422),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2422),
.Y(n_2769)
);

BUFx6f_ASAP7_75t_L g2770 ( 
.A(n_2072),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2117),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2118),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2424),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2424),
.Y(n_2774)
);

INVxp33_ASAP7_75t_SL g2775 ( 
.A(n_2187),
.Y(n_2775)
);

BUFx2_ASAP7_75t_L g2776 ( 
.A(n_2414),
.Y(n_2776)
);

INVx3_ASAP7_75t_L g2777 ( 
.A(n_2425),
.Y(n_2777)
);

NOR2xp33_ASAP7_75t_L g2778 ( 
.A(n_2109),
.B(n_1824),
.Y(n_2778)
);

INVx2_ASAP7_75t_SL g2779 ( 
.A(n_2257),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2425),
.Y(n_2780)
);

INVx2_ASAP7_75t_SL g2781 ( 
.A(n_2257),
.Y(n_2781)
);

NOR2xp33_ASAP7_75t_L g2782 ( 
.A(n_2109),
.B(n_1825),
.Y(n_2782)
);

BUFx16f_ASAP7_75t_R g2783 ( 
.A(n_2150),
.Y(n_2783)
);

OR2x2_ASAP7_75t_L g2784 ( 
.A(n_2196),
.B(n_1976),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2119),
.Y(n_2785)
);

INVx3_ASAP7_75t_L g2786 ( 
.A(n_2438),
.Y(n_2786)
);

INVx3_ASAP7_75t_L g2787 ( 
.A(n_2438),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2120),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2404),
.B(n_2362),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2450),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2450),
.Y(n_2791)
);

INVxp67_ASAP7_75t_SL g2792 ( 
.A(n_2072),
.Y(n_2792)
);

INVx3_ASAP7_75t_L g2793 ( 
.A(n_2452),
.Y(n_2793)
);

INVx3_ASAP7_75t_L g2794 ( 
.A(n_2452),
.Y(n_2794)
);

NAND2xp33_ASAP7_75t_L g2795 ( 
.A(n_2179),
.B(n_1749),
.Y(n_2795)
);

NOR2x1p5_ASAP7_75t_L g2796 ( 
.A(n_2188),
.B(n_1832),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_SL g2797 ( 
.A(n_2304),
.B(n_1865),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2454),
.Y(n_2798)
);

INVx8_ASAP7_75t_L g2799 ( 
.A(n_2202),
.Y(n_2799)
);

BUFx6f_ASAP7_75t_SL g2800 ( 
.A(n_2290),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2454),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2217),
.Y(n_2802)
);

BUFx10_ASAP7_75t_L g2803 ( 
.A(n_2039),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2217),
.Y(n_2804)
);

BUFx6f_ASAP7_75t_SL g2805 ( 
.A(n_2290),
.Y(n_2805)
);

INVxp33_ASAP7_75t_SL g2806 ( 
.A(n_2092),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2217),
.Y(n_2807)
);

CKINVDCx5p33_ASAP7_75t_R g2808 ( 
.A(n_2428),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2050),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2122),
.B(n_1825),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_2150),
.Y(n_2811)
);

INVxp67_ASAP7_75t_SL g2812 ( 
.A(n_2083),
.Y(n_2812)
);

INVx2_ASAP7_75t_SL g2813 ( 
.A(n_2257),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2050),
.Y(n_2814)
);

NOR2xp33_ASAP7_75t_L g2815 ( 
.A(n_2138),
.B(n_1844),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_L g2816 ( 
.A(n_2196),
.B(n_1844),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2050),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_SL g2818 ( 
.A(n_2135),
.B(n_1964),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_L g2819 ( 
.A(n_2228),
.B(n_1865),
.Y(n_2819)
);

INVx5_ASAP7_75t_L g2820 ( 
.A(n_2285),
.Y(n_2820)
);

INVx2_ASAP7_75t_SL g2821 ( 
.A(n_2281),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2054),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2054),
.Y(n_2823)
);

INVxp33_ASAP7_75t_SL g2824 ( 
.A(n_2080),
.Y(n_2824)
);

BUFx6f_ASAP7_75t_SL g2825 ( 
.A(n_2290),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2076),
.Y(n_2826)
);

INVxp33_ASAP7_75t_L g2827 ( 
.A(n_2409),
.Y(n_2827)
);

INVx3_ASAP7_75t_L g2828 ( 
.A(n_2251),
.Y(n_2828)
);

INVx2_ASAP7_75t_SL g2829 ( 
.A(n_2281),
.Y(n_2829)
);

INVx3_ASAP7_75t_L g2830 ( 
.A(n_2251),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2362),
.B(n_1854),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_SL g2832 ( 
.A(n_2115),
.B(n_1877),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2362),
.B(n_1854),
.Y(n_2833)
);

NAND2xp33_ASAP7_75t_L g2834 ( 
.A(n_2202),
.B(n_1749),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2054),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2251),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2121),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2078),
.Y(n_2838)
);

CKINVDCx5p33_ASAP7_75t_R g2839 ( 
.A(n_2220),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2396),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2396),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2079),
.Y(n_2842)
);

INVx3_ASAP7_75t_L g2843 ( 
.A(n_2042),
.Y(n_2843)
);

NAND3xp33_ASAP7_75t_L g2844 ( 
.A(n_2416),
.B(n_1976),
.C(n_1785),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2081),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2082),
.Y(n_2846)
);

AO21x2_ASAP7_75t_L g2847 ( 
.A1(n_2207),
.A2(n_1785),
.B(n_1987),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2362),
.B(n_2202),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2087),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2202),
.B(n_1854),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2095),
.Y(n_2851)
);

NAND2xp33_ASAP7_75t_L g2852 ( 
.A(n_2202),
.B(n_1749),
.Y(n_2852)
);

NAND2xp33_ASAP7_75t_SL g2853 ( 
.A(n_2211),
.B(n_1735),
.Y(n_2853)
);

CKINVDCx5p33_ASAP7_75t_R g2854 ( 
.A(n_2220),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2098),
.Y(n_2855)
);

NOR2xp33_ASAP7_75t_L g2856 ( 
.A(n_2228),
.B(n_1877),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2042),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2233),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2233),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_SL g2860 ( 
.A(n_2236),
.B(n_1883),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2056),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2056),
.Y(n_2862)
);

OAI22xp33_ASAP7_75t_L g2863 ( 
.A1(n_2274),
.A2(n_1921),
.B1(n_1948),
.B2(n_1906),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2162),
.B(n_1983),
.Y(n_2864)
);

AND3x1_ASAP7_75t_L g2865 ( 
.A(n_2276),
.B(n_1921),
.C(n_1906),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2094),
.Y(n_2866)
);

NAND2xp33_ASAP7_75t_L g2867 ( 
.A(n_2285),
.B(n_1749),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2094),
.Y(n_2868)
);

NOR2xp33_ASAP7_75t_L g2869 ( 
.A(n_2352),
.B(n_1948),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2418),
.Y(n_2870)
);

BUFx6f_ASAP7_75t_SL g2871 ( 
.A(n_2124),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2167),
.B(n_1983),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2418),
.Y(n_2873)
);

NOR2xp33_ASAP7_75t_L g2874 ( 
.A(n_2352),
.B(n_1964),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2170),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2103),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2182),
.B(n_1983),
.Y(n_2877)
);

INVx3_ASAP7_75t_L g2878 ( 
.A(n_2103),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2110),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2170),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2184),
.Y(n_2881)
);

BUFx6f_ASAP7_75t_SL g2882 ( 
.A(n_2124),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_SL g2883 ( 
.A(n_2429),
.B(n_1998),
.Y(n_2883)
);

BUFx6f_ASAP7_75t_L g2884 ( 
.A(n_2534),
.Y(n_2884)
);

AND2x2_ASAP7_75t_L g2885 ( 
.A(n_2604),
.B(n_1979),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2455),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2455),
.Y(n_2887)
);

INVx2_ASAP7_75t_SL g2888 ( 
.A(n_2609),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2469),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2469),
.Y(n_2890)
);

BUFx3_ASAP7_75t_L g2891 ( 
.A(n_2776),
.Y(n_2891)
);

AND2x2_ASAP7_75t_SL g2892 ( 
.A(n_2503),
.B(n_2382),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2563),
.B(n_2045),
.Y(n_2893)
);

NOR2xp33_ASAP7_75t_L g2894 ( 
.A(n_2565),
.B(n_2089),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2471),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_L g2896 ( 
.A(n_2554),
.B(n_2039),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2471),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2459),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2473),
.Y(n_2899)
);

AND2x4_ASAP7_75t_L g2900 ( 
.A(n_2534),
.B(n_2140),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2473),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2475),
.Y(n_2902)
);

OR2x2_ASAP7_75t_L g2903 ( 
.A(n_2556),
.B(n_1979),
.Y(n_2903)
);

CKINVDCx20_ASAP7_75t_R g2904 ( 
.A(n_2594),
.Y(n_2904)
);

CKINVDCx20_ASAP7_75t_R g2905 ( 
.A(n_2594),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2475),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2500),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2500),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2535),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2535),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2540),
.Y(n_2911)
);

NOR2xp33_ASAP7_75t_L g2912 ( 
.A(n_2627),
.B(n_1998),
.Y(n_2912)
);

BUFx6f_ASAP7_75t_L g2913 ( 
.A(n_2652),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2585),
.B(n_2045),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2540),
.Y(n_2915)
);

NAND2x1p5_ASAP7_75t_L g2916 ( 
.A(n_2479),
.B(n_2449),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2541),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2541),
.Y(n_2918)
);

BUFx8_ASAP7_75t_L g2919 ( 
.A(n_2560),
.Y(n_2919)
);

BUFx6f_ASAP7_75t_SL g2920 ( 
.A(n_2456),
.Y(n_2920)
);

AND2x2_ASAP7_75t_L g2921 ( 
.A(n_2477),
.B(n_2429),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2459),
.Y(n_2922)
);

NAND2xp33_ASAP7_75t_R g2923 ( 
.A(n_2806),
.B(n_2381),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2557),
.Y(n_2924)
);

NOR2xp33_ASAP7_75t_L g2925 ( 
.A(n_2635),
.B(n_2139),
.Y(n_2925)
);

NOR2xp33_ASAP7_75t_L g2926 ( 
.A(n_2617),
.B(n_2639),
.Y(n_2926)
);

CKINVDCx20_ASAP7_75t_R g2927 ( 
.A(n_2658),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2557),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2558),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2558),
.Y(n_2930)
);

BUFx6f_ASAP7_75t_L g2931 ( 
.A(n_2652),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2629),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2481),
.B(n_2045),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2477),
.B(n_2191),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2629),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2630),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2630),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2666),
.Y(n_2938)
);

NAND2xp33_ASAP7_75t_R g2939 ( 
.A(n_2806),
.B(n_2381),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2666),
.Y(n_2940)
);

AND2x2_ASAP7_75t_L g2941 ( 
.A(n_2470),
.B(n_2191),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2668),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2668),
.Y(n_2943)
);

CKINVDCx5p33_ASAP7_75t_R g2944 ( 
.A(n_2519),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2669),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2460),
.Y(n_2946)
);

NOR2xp33_ASAP7_75t_L g2947 ( 
.A(n_2484),
.B(n_2139),
.Y(n_2947)
);

XOR2xp5_ASAP7_75t_L g2948 ( 
.A(n_2519),
.B(n_2654),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2669),
.Y(n_2949)
);

XOR2xp5_ASAP7_75t_L g2950 ( 
.A(n_2654),
.B(n_1443),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2671),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2671),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2622),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2460),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_SL g2955 ( 
.A(n_2478),
.B(n_2183),
.Y(n_2955)
);

BUFx3_ASAP7_75t_L g2956 ( 
.A(n_2776),
.Y(n_2956)
);

CKINVDCx20_ASAP7_75t_R g2957 ( 
.A(n_2658),
.Y(n_2957)
);

XOR2xp5_ASAP7_75t_L g2958 ( 
.A(n_2693),
.B(n_1458),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2622),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2624),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2624),
.Y(n_2961)
);

XNOR2x2_ASAP7_75t_L g2962 ( 
.A(n_2606),
.B(n_1889),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2632),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2470),
.B(n_2206),
.Y(n_2964)
);

INVx2_ASAP7_75t_SL g2965 ( 
.A(n_2609),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2632),
.Y(n_2966)
);

INVx1_ASAP7_75t_SL g2967 ( 
.A(n_2458),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2524),
.B(n_2310),
.Y(n_2968)
);

NOR2xp33_ASAP7_75t_L g2969 ( 
.A(n_2568),
.B(n_2377),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2637),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2637),
.Y(n_2971)
);

NOR2xp67_ASAP7_75t_L g2972 ( 
.A(n_2649),
.B(n_1961),
.Y(n_2972)
);

INVx2_ASAP7_75t_SL g2973 ( 
.A(n_2458),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2638),
.Y(n_2974)
);

INVx2_ASAP7_75t_SL g2975 ( 
.A(n_2472),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2638),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2643),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2643),
.Y(n_2978)
);

AND2x6_ASAP7_75t_L g2979 ( 
.A(n_2809),
.B(n_2140),
.Y(n_2979)
);

NOR2xp33_ASAP7_75t_L g2980 ( 
.A(n_2626),
.B(n_2377),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_2626),
.B(n_2317),
.Y(n_2981)
);

XOR2xp5_ASAP7_75t_L g2982 ( 
.A(n_2693),
.B(n_2827),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2463),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_SL g2984 ( 
.A(n_2636),
.B(n_2206),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2644),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2644),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2621),
.B(n_2208),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2646),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2646),
.Y(n_2989)
);

OR2x2_ASAP7_75t_L g2990 ( 
.A(n_2490),
.B(n_1795),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2463),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2650),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2650),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2465),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2553),
.B(n_2208),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2651),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2651),
.Y(n_2997)
);

NOR2xp33_ASAP7_75t_L g2998 ( 
.A(n_2488),
.B(n_2498),
.Y(n_2998)
);

NOR2xp33_ASAP7_75t_L g2999 ( 
.A(n_2574),
.B(n_2530),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2661),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_L g3001 ( 
.A(n_2530),
.B(n_1796),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2661),
.Y(n_3002)
);

NAND2x1p5_ASAP7_75t_L g3003 ( 
.A(n_2479),
.B(n_2449),
.Y(n_3003)
);

BUFx3_ASAP7_75t_L g3004 ( 
.A(n_2472),
.Y(n_3004)
);

NOR2xp33_ASAP7_75t_L g3005 ( 
.A(n_2530),
.B(n_1803),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2663),
.Y(n_3006)
);

XNOR2xp5_ASAP7_75t_L g3007 ( 
.A(n_2827),
.B(n_2159),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2663),
.Y(n_3008)
);

XOR2xp5_ASAP7_75t_L g3009 ( 
.A(n_2808),
.B(n_1458),
.Y(n_3009)
);

AND2x4_ASAP7_75t_L g3010 ( 
.A(n_2614),
.B(n_2254),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2664),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2664),
.Y(n_3012)
);

NOR2xp33_ASAP7_75t_SL g3013 ( 
.A(n_2503),
.B(n_1896),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2465),
.Y(n_3014)
);

AND2x2_ASAP7_75t_L g3015 ( 
.A(n_2468),
.B(n_2254),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2665),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2665),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2674),
.Y(n_3018)
);

BUFx6f_ASAP7_75t_L g3019 ( 
.A(n_2504),
.Y(n_3019)
);

AND2x2_ASAP7_75t_L g3020 ( 
.A(n_2468),
.B(n_2461),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2703),
.B(n_2262),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2697),
.B(n_2262),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2674),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2675),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2675),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2678),
.Y(n_3026)
);

OR2x2_ASAP7_75t_SL g3027 ( 
.A(n_2844),
.B(n_2248),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2678),
.Y(n_3028)
);

NOR2xp33_ASAP7_75t_L g3029 ( 
.A(n_2509),
.B(n_1819),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2679),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2679),
.Y(n_3031)
);

XOR2xp5_ASAP7_75t_L g3032 ( 
.A(n_2808),
.B(n_1472),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2680),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2680),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2685),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2697),
.B(n_1983),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2685),
.Y(n_3037)
);

XNOR2x2_ASAP7_75t_L g3038 ( 
.A(n_2682),
.B(n_1735),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2686),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2730),
.B(n_1983),
.Y(n_3040)
);

AOI21xp5_ASAP7_75t_L g3041 ( 
.A1(n_2747),
.A2(n_2426),
.B(n_2285),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_2461),
.B(n_1827),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2686),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2730),
.B(n_2281),
.Y(n_3044)
);

OR2x2_ASAP7_75t_L g3045 ( 
.A(n_2490),
.B(n_2201),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2687),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2687),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2466),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_SL g3049 ( 
.A(n_2720),
.B(n_1896),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2466),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2570),
.B(n_2159),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2467),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2467),
.Y(n_3053)
);

INVxp67_ASAP7_75t_SL g3054 ( 
.A(n_2504),
.Y(n_3054)
);

OAI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2809),
.A2(n_2329),
.B(n_2326),
.Y(n_3055)
);

CKINVDCx20_ASAP7_75t_R g3056 ( 
.A(n_2811),
.Y(n_3056)
);

INVxp33_ASAP7_75t_L g3057 ( 
.A(n_2584),
.Y(n_3057)
);

BUFx6f_ASAP7_75t_SL g3058 ( 
.A(n_2456),
.Y(n_3058)
);

INVx1_ASAP7_75t_SL g3059 ( 
.A(n_2526),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2667),
.B(n_2334),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2480),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2480),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2482),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2482),
.Y(n_3064)
);

BUFx3_ASAP7_75t_L g3065 ( 
.A(n_2526),
.Y(n_3065)
);

AOI21xp5_ASAP7_75t_L g3066 ( 
.A1(n_2802),
.A2(n_2449),
.B(n_2426),
.Y(n_3066)
);

BUFx6f_ASAP7_75t_SL g3067 ( 
.A(n_2456),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2487),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2487),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2510),
.Y(n_3070)
);

CKINVDCx20_ASAP7_75t_R g3071 ( 
.A(n_2811),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2510),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2511),
.Y(n_3073)
);

XNOR2xp5_ASAP7_75t_L g3074 ( 
.A(n_2699),
.B(n_1472),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2695),
.B(n_2335),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2511),
.Y(n_3076)
);

INVx4_ASAP7_75t_SL g3077 ( 
.A(n_2559),
.Y(n_3077)
);

XOR2xp5_ASAP7_75t_L g3078 ( 
.A(n_2839),
.B(n_1475),
.Y(n_3078)
);

XNOR2x2_ASAP7_75t_L g3079 ( 
.A(n_2778),
.B(n_1055),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2514),
.Y(n_3080)
);

NOR2xp33_ASAP7_75t_L g3081 ( 
.A(n_2536),
.B(n_1766),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2514),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2517),
.Y(n_3083)
);

CKINVDCx20_ASAP7_75t_R g3084 ( 
.A(n_2839),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_SL g3085 ( 
.A(n_2722),
.B(n_1901),
.Y(n_3085)
);

NOR2xp33_ASAP7_75t_L g3086 ( 
.A(n_2570),
.B(n_1770),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2517),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2521),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2521),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2695),
.B(n_2336),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2525),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2525),
.Y(n_3092)
);

INVx2_ASAP7_75t_L g3093 ( 
.A(n_2527),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2479),
.B(n_2337),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2527),
.Y(n_3095)
);

AND2x4_ASAP7_75t_L g3096 ( 
.A(n_2614),
.B(n_1851),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2529),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2529),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2531),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2531),
.Y(n_3100)
);

OR2x2_ASAP7_75t_L g3101 ( 
.A(n_2544),
.B(n_1845),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_2532),
.Y(n_3102)
);

AOI21x1_ASAP7_75t_L g3103 ( 
.A1(n_2634),
.A2(n_2341),
.B(n_2338),
.Y(n_3103)
);

XOR2xp5_ASAP7_75t_L g3104 ( 
.A(n_2854),
.B(n_1475),
.Y(n_3104)
);

BUFx3_ASAP7_75t_L g3105 ( 
.A(n_2544),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2532),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2533),
.Y(n_3107)
);

CKINVDCx5p33_ASAP7_75t_R g3108 ( 
.A(n_2871),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2533),
.Y(n_3109)
);

INVx2_ASAP7_75t_SL g3110 ( 
.A(n_2623),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2537),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2537),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2538),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2538),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2539),
.Y(n_3115)
);

AND2x2_ASAP7_75t_L g3116 ( 
.A(n_2618),
.B(n_1901),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2539),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2542),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2542),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_L g3120 ( 
.A(n_2618),
.B(n_2003),
.Y(n_3120)
);

INVx1_ASAP7_75t_SL g3121 ( 
.A(n_2507),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_2507),
.B(n_2003),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2543),
.Y(n_3123)
);

AND2x2_ASAP7_75t_L g3124 ( 
.A(n_2709),
.B(n_2816),
.Y(n_3124)
);

CKINVDCx16_ASAP7_75t_R g3125 ( 
.A(n_2871),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2543),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2547),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_2547),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2548),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2479),
.B(n_2342),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_2709),
.B(n_1503),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2548),
.Y(n_3132)
);

XNOR2x2_ASAP7_75t_L g3133 ( 
.A(n_2782),
.B(n_1056),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2552),
.Y(n_3134)
);

XNOR2x2_ASAP7_75t_L g3135 ( 
.A(n_2810),
.B(n_1056),
.Y(n_3135)
);

NAND2xp33_ASAP7_75t_SL g3136 ( 
.A(n_2871),
.B(n_1850),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2552),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2586),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2586),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2588),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2588),
.Y(n_3141)
);

XOR2xp5_ASAP7_75t_L g3142 ( 
.A(n_2854),
.B(n_1478),
.Y(n_3142)
);

AND2x2_ASAP7_75t_L g3143 ( 
.A(n_2819),
.B(n_1505),
.Y(n_3143)
);

CKINVDCx5p33_ASAP7_75t_R g3144 ( 
.A(n_2882),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2590),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_2856),
.B(n_1505),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2590),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2597),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2597),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2598),
.Y(n_3150)
);

NOR2xp67_ASAP7_75t_L g3151 ( 
.A(n_2869),
.B(n_1699),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2598),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2479),
.B(n_2348),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_SL g3154 ( 
.A(n_2711),
.B(n_2426),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2600),
.Y(n_3155)
);

NAND2xp33_ASAP7_75t_R g3156 ( 
.A(n_2824),
.B(n_1870),
.Y(n_3156)
);

NOR2xp33_ASAP7_75t_L g3157 ( 
.A(n_2784),
.B(n_1776),
.Y(n_3157)
);

CKINVDCx16_ASAP7_75t_R g3158 ( 
.A(n_2882),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_2600),
.Y(n_3159)
);

NAND2x1p5_ASAP7_75t_L g3160 ( 
.A(n_2581),
.B(n_2449),
.Y(n_3160)
);

AND2x4_ASAP7_75t_L g3161 ( 
.A(n_2614),
.B(n_1870),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2602),
.Y(n_3162)
);

INVxp33_ASAP7_75t_L g3163 ( 
.A(n_2815),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2602),
.Y(n_3164)
);

AND2x2_ASAP7_75t_L g3165 ( 
.A(n_2742),
.B(n_2745),
.Y(n_3165)
);

XNOR2xp5_ASAP7_75t_L g3166 ( 
.A(n_2796),
.B(n_1478),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2607),
.Y(n_3167)
);

INVx4_ASAP7_75t_SL g3168 ( 
.A(n_2559),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2607),
.Y(n_3169)
);

XNOR2xp5_ASAP7_75t_L g3170 ( 
.A(n_2508),
.B(n_1523),
.Y(n_3170)
);

NOR2xp33_ASAP7_75t_L g3171 ( 
.A(n_2784),
.B(n_1776),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_2689),
.B(n_2349),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2613),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2613),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2616),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2616),
.Y(n_3176)
);

INVxp67_ASAP7_75t_SL g3177 ( 
.A(n_2504),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2619),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2619),
.Y(n_3179)
);

INVxp67_ASAP7_75t_SL g3180 ( 
.A(n_2504),
.Y(n_3180)
);

XOR2xp5_ASAP7_75t_L g3181 ( 
.A(n_2775),
.B(n_1523),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2881),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2881),
.Y(n_3183)
);

NOR2xp33_ASAP7_75t_L g3184 ( 
.A(n_2633),
.B(n_1853),
.Y(n_3184)
);

INVxp33_ASAP7_75t_L g3185 ( 
.A(n_2874),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2576),
.Y(n_3186)
);

XOR2xp5_ASAP7_75t_L g3187 ( 
.A(n_2775),
.B(n_1550),
.Y(n_3187)
);

NOR2xp33_ASAP7_75t_L g3188 ( 
.A(n_2633),
.B(n_1856),
.Y(n_3188)
);

CKINVDCx20_ASAP7_75t_R g3189 ( 
.A(n_2491),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2580),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2582),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2591),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2701),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2712),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2714),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2464),
.Y(n_3196)
);

BUFx6f_ASAP7_75t_L g3197 ( 
.A(n_2504),
.Y(n_3197)
);

XNOR2xp5_ASAP7_75t_L g3198 ( 
.A(n_2555),
.B(n_1550),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_2464),
.Y(n_3199)
);

XOR2xp5_ASAP7_75t_L g3200 ( 
.A(n_2824),
.B(n_1605),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2715),
.Y(n_3201)
);

NOR2xp33_ASAP7_75t_L g3202 ( 
.A(n_2633),
.B(n_1991),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2710),
.B(n_2351),
.Y(n_3203)
);

XOR2xp5_ASAP7_75t_L g3204 ( 
.A(n_2474),
.B(n_1605),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2717),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_2464),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2723),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2725),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2727),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2657),
.B(n_2354),
.Y(n_3210)
);

XNOR2xp5_ASAP7_75t_SL g3211 ( 
.A(n_2749),
.B(n_1997),
.Y(n_3211)
);

INVxp67_ASAP7_75t_SL g3212 ( 
.A(n_2575),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2734),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2735),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2736),
.Y(n_3215)
);

XOR2xp5_ASAP7_75t_L g3216 ( 
.A(n_2474),
.B(n_1643),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2739),
.Y(n_3217)
);

OR2x2_ASAP7_75t_L g3218 ( 
.A(n_2647),
.B(n_1446),
.Y(n_3218)
);

OR2x2_ASAP7_75t_L g3219 ( 
.A(n_2457),
.B(n_1479),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_2742),
.B(n_1598),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2485),
.Y(n_3221)
);

XOR2xp5_ASAP7_75t_L g3222 ( 
.A(n_2759),
.B(n_1643),
.Y(n_3222)
);

OR2x6_ASAP7_75t_L g3223 ( 
.A(n_2456),
.B(n_2577),
.Y(n_3223)
);

NOR2xp33_ASAP7_75t_L g3224 ( 
.A(n_2605),
.B(n_1660),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2489),
.Y(n_3225)
);

BUFx6f_ASAP7_75t_L g3226 ( 
.A(n_2575),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_2492),
.Y(n_3227)
);

INVxp33_ASAP7_75t_SL g3228 ( 
.A(n_2546),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2493),
.Y(n_3229)
);

AND2x2_ASAP7_75t_L g3230 ( 
.A(n_2745),
.B(n_1598),
.Y(n_3230)
);

XOR2xp5_ASAP7_75t_L g3231 ( 
.A(n_2700),
.B(n_1660),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2494),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_2495),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2496),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2502),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2476),
.Y(n_3236)
);

NOR2xp33_ASAP7_75t_SL g3237 ( 
.A(n_2803),
.B(n_1717),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2512),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2476),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2476),
.Y(n_3240)
);

INVx8_ASAP7_75t_L g3241 ( 
.A(n_2882),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_2513),
.B(n_1622),
.Y(n_3242)
);

CKINVDCx20_ASAP7_75t_R g3243 ( 
.A(n_2803),
.Y(n_3243)
);

INVx2_ASAP7_75t_SL g3244 ( 
.A(n_2883),
.Y(n_3244)
);

AND2x2_ASAP7_75t_L g3245 ( 
.A(n_2515),
.B(n_1622),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_2518),
.Y(n_3246)
);

INVxp67_ASAP7_75t_SL g3247 ( 
.A(n_2575),
.Y(n_3247)
);

INVx3_ASAP7_75t_R g3248 ( 
.A(n_2766),
.Y(n_3248)
);

CKINVDCx20_ASAP7_75t_R g3249 ( 
.A(n_2803),
.Y(n_3249)
);

AND2x4_ASAP7_75t_L g3250 ( 
.A(n_2683),
.B(n_1933),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_L g3251 ( 
.A(n_2605),
.B(n_1629),
.Y(n_3251)
);

INVxp33_ASAP7_75t_L g3252 ( 
.A(n_2694),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_2520),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2523),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2567),
.Y(n_3255)
);

NOR2xp33_ASAP7_75t_L g3256 ( 
.A(n_2605),
.B(n_1629),
.Y(n_3256)
);

XNOR2x2_ASAP7_75t_L g3257 ( 
.A(n_2818),
.B(n_1062),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2798),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2798),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_2826),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2826),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2611),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_2612),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2615),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2620),
.Y(n_3265)
);

INVxp33_ASAP7_75t_L g3266 ( 
.A(n_2797),
.Y(n_3266)
);

INVx3_ASAP7_75t_L g3267 ( 
.A(n_2692),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_2564),
.B(n_2549),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2642),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2645),
.Y(n_3270)
);

BUFx3_ASAP7_75t_L g3271 ( 
.A(n_2766),
.Y(n_3271)
);

CKINVDCx20_ASAP7_75t_R g3272 ( 
.A(n_2853),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2648),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_2655),
.Y(n_3274)
);

AND2x2_ASAP7_75t_L g3275 ( 
.A(n_2564),
.B(n_2765),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_2660),
.B(n_2356),
.Y(n_3276)
);

CKINVDCx20_ASAP7_75t_R g3277 ( 
.A(n_2853),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_2765),
.B(n_1658),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_2486),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_2486),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2752),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2753),
.Y(n_3282)
);

AND2x2_ASAP7_75t_L g3283 ( 
.A(n_2641),
.B(n_1658),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2755),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2757),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_2764),
.Y(n_3286)
);

CKINVDCx5p33_ASAP7_75t_R g3287 ( 
.A(n_2726),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_2486),
.Y(n_3288)
);

NOR2xp33_ASAP7_75t_L g3289 ( 
.A(n_2505),
.B(n_2365),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_2771),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2772),
.Y(n_3291)
);

NOR2xp33_ASAP7_75t_L g3292 ( 
.A(n_2506),
.B(n_2368),
.Y(n_3292)
);

HB1xp67_ASAP7_75t_L g3293 ( 
.A(n_2858),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_2785),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_2788),
.Y(n_3295)
);

AND2x2_ASAP7_75t_SL g3296 ( 
.A(n_2581),
.B(n_1062),
.Y(n_3296)
);

OR2x6_ASAP7_75t_L g3297 ( 
.A(n_2577),
.B(n_1736),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2837),
.Y(n_3298)
);

NOR2xp33_ASAP7_75t_L g3299 ( 
.A(n_2545),
.B(n_2394),
.Y(n_3299)
);

CKINVDCx20_ASAP7_75t_R g3300 ( 
.A(n_2566),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2569),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_2569),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2569),
.Y(n_3303)
);

INVxp33_ASAP7_75t_L g3304 ( 
.A(n_2690),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2572),
.Y(n_3305)
);

XOR2xp5_ASAP7_75t_L g3306 ( 
.A(n_2700),
.B(n_2246),
.Y(n_3306)
);

INVx2_ASAP7_75t_SL g3307 ( 
.A(n_2737),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_SL g3308 ( 
.A(n_2599),
.B(n_2551),
.Y(n_3308)
);

NOR2xp33_ASAP7_75t_L g3309 ( 
.A(n_2562),
.B(n_2395),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_2572),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_2572),
.Y(n_3311)
);

AOI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_2802),
.A2(n_2426),
.B(n_2359),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2573),
.Y(n_3313)
);

INVxp67_ASAP7_75t_L g3314 ( 
.A(n_2566),
.Y(n_3314)
);

AND2x2_ASAP7_75t_L g3315 ( 
.A(n_2885),
.B(n_2737),
.Y(n_3315)
);

BUFx2_ASAP7_75t_L g3316 ( 
.A(n_2891),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_SL g3317 ( 
.A(n_2947),
.B(n_2641),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_2898),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_2998),
.B(n_2662),
.Y(n_3319)
);

AOI21xp5_ASAP7_75t_L g3320 ( 
.A1(n_2914),
.A2(n_2581),
.B(n_2592),
.Y(n_3320)
);

NOR2xp33_ASAP7_75t_L g3321 ( 
.A(n_2926),
.B(n_2601),
.Y(n_3321)
);

AOI22xp33_ASAP7_75t_L g3322 ( 
.A1(n_2926),
.A2(n_2587),
.B1(n_2559),
.B2(n_2858),
.Y(n_3322)
);

NOR2xp33_ASAP7_75t_L g3323 ( 
.A(n_3185),
.B(n_2832),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3143),
.B(n_3146),
.Y(n_3324)
);

NOR2xp67_ASAP7_75t_SL g3325 ( 
.A(n_3125),
.B(n_2789),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_2886),
.Y(n_3326)
);

OAI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_2933),
.A2(n_2733),
.B(n_2698),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_2998),
.B(n_2859),
.Y(n_3328)
);

OR2x2_ASAP7_75t_L g3329 ( 
.A(n_2903),
.B(n_2860),
.Y(n_3329)
);

INVx2_ASAP7_75t_SL g3330 ( 
.A(n_2956),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2968),
.B(n_2925),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_2887),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2968),
.B(n_2859),
.Y(n_3333)
);

NAND3xp33_ASAP7_75t_L g3334 ( 
.A(n_2912),
.B(n_2587),
.C(n_2705),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_SL g3335 ( 
.A(n_2947),
.B(n_2673),
.Y(n_3335)
);

OAI22xp33_ASAP7_75t_L g3336 ( 
.A1(n_3163),
.A2(n_2673),
.B1(n_2841),
.B2(n_2840),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_2925),
.B(n_2528),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_2981),
.B(n_2528),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_2981),
.B(n_2528),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_L g3340 ( 
.A(n_3228),
.B(n_2999),
.Y(n_3340)
);

NOR2xp33_ASAP7_75t_L g3341 ( 
.A(n_2999),
.B(n_2863),
.Y(n_3341)
);

OR2x2_ASAP7_75t_L g3342 ( 
.A(n_3121),
.B(n_2713),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_2922),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3021),
.B(n_2559),
.Y(n_3344)
);

AND2x6_ASAP7_75t_L g3345 ( 
.A(n_2914),
.B(n_2814),
.Y(n_3345)
);

INVx3_ASAP7_75t_L g3346 ( 
.A(n_3019),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3021),
.B(n_2559),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3314),
.B(n_2559),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3314),
.B(n_2698),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_SL g3350 ( 
.A(n_2894),
.B(n_2483),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2896),
.B(n_2733),
.Y(n_3351)
);

INVxp67_ASAP7_75t_L g3352 ( 
.A(n_3110),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_SL g3353 ( 
.A(n_2894),
.B(n_2483),
.Y(n_3353)
);

NOR2xp33_ASAP7_75t_L g3354 ( 
.A(n_2912),
.B(n_2501),
.Y(n_3354)
);

AND2x2_ASAP7_75t_L g3355 ( 
.A(n_3220),
.B(n_2719),
.Y(n_3355)
);

AOI22xp33_ASAP7_75t_L g3356 ( 
.A1(n_2896),
.A2(n_2684),
.B1(n_2497),
.B2(n_2847),
.Y(n_3356)
);

NOR2xp33_ASAP7_75t_L g3357 ( 
.A(n_3029),
.B(n_2589),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_2980),
.B(n_2767),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_2980),
.B(n_2767),
.Y(n_3359)
);

NOR2xp33_ASAP7_75t_L g3360 ( 
.A(n_3029),
.B(n_2740),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_2889),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_2890),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_SL g3363 ( 
.A(n_2995),
.B(n_2683),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3081),
.B(n_2684),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2895),
.Y(n_3365)
);

O2A1O1Ixp5_ASAP7_75t_L g3366 ( 
.A1(n_3308),
.A2(n_2634),
.B(n_2640),
.C(n_2625),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_SL g3367 ( 
.A(n_2995),
.B(n_2683),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3081),
.B(n_2684),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_3086),
.B(n_2760),
.Y(n_3369)
);

INVx2_ASAP7_75t_SL g3370 ( 
.A(n_3004),
.Y(n_3370)
);

INVx2_ASAP7_75t_SL g3371 ( 
.A(n_3065),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3086),
.B(n_2684),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_2946),
.Y(n_3373)
);

INVx2_ASAP7_75t_SL g3374 ( 
.A(n_3105),
.Y(n_3374)
);

BUFx3_ASAP7_75t_L g3375 ( 
.A(n_3271),
.Y(n_3375)
);

NOR2xp33_ASAP7_75t_L g3376 ( 
.A(n_3121),
.B(n_3251),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_2897),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_3251),
.B(n_2751),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3268),
.B(n_2684),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_3020),
.B(n_2684),
.Y(n_3380)
);

AOI22xp33_ASAP7_75t_L g3381 ( 
.A1(n_2969),
.A2(n_2497),
.B1(n_2847),
.B2(n_2870),
.Y(n_3381)
);

A2O1A1Ixp33_ASAP7_75t_L g3382 ( 
.A1(n_2969),
.A2(n_2848),
.B(n_2603),
.C(n_2595),
.Y(n_3382)
);

INVx2_ASAP7_75t_SL g3383 ( 
.A(n_2973),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_2899),
.Y(n_3384)
);

AND2x2_ASAP7_75t_L g3385 ( 
.A(n_3230),
.B(n_2497),
.Y(n_3385)
);

INVxp67_ASAP7_75t_L g3386 ( 
.A(n_2967),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3293),
.B(n_2779),
.Y(n_3387)
);

NOR2xp67_ASAP7_75t_L g3388 ( 
.A(n_2944),
.B(n_2681),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3293),
.B(n_2779),
.Y(n_3389)
);

AND2x2_ASAP7_75t_L g3390 ( 
.A(n_3278),
.B(n_2873),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3060),
.B(n_2781),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3060),
.B(n_2781),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_2901),
.Y(n_3393)
);

NOR2x1p5_ASAP7_75t_L g3394 ( 
.A(n_3108),
.B(n_1928),
.Y(n_3394)
);

AOI221xp5_ASAP7_75t_L g3395 ( 
.A1(n_3222),
.A2(n_2865),
.B1(n_1641),
.B2(n_1559),
.C(n_2653),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_SL g3396 ( 
.A(n_2921),
.B(n_2659),
.Y(n_3396)
);

NOR2xp33_ASAP7_75t_L g3397 ( 
.A(n_3256),
.B(n_2875),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3172),
.B(n_3203),
.Y(n_3398)
);

NOR2x1p5_ASAP7_75t_L g3399 ( 
.A(n_3144),
.B(n_2880),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_SL g3400 ( 
.A(n_3001),
.B(n_2813),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_SL g3401 ( 
.A(n_3001),
.B(n_2813),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3172),
.B(n_2821),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_2902),
.Y(n_3403)
);

NOR2xp33_ASAP7_75t_L g3404 ( 
.A(n_3256),
.B(n_2726),
.Y(n_3404)
);

INVxp67_ASAP7_75t_L g3405 ( 
.A(n_2967),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_2954),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3203),
.B(n_3022),
.Y(n_3407)
);

NAND2x1_ASAP7_75t_L g3408 ( 
.A(n_3267),
.B(n_2843),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3022),
.B(n_2821),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2906),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_SL g3411 ( 
.A(n_3005),
.B(n_2829),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_L g3412 ( 
.A(n_2955),
.B(n_2726),
.Y(n_3412)
);

INVx3_ASAP7_75t_L g3413 ( 
.A(n_3019),
.Y(n_3413)
);

AOI22xp5_ASAP7_75t_L g3414 ( 
.A1(n_3300),
.A2(n_2847),
.B1(n_2838),
.B2(n_2845),
.Y(n_3414)
);

INVx4_ASAP7_75t_L g3415 ( 
.A(n_2884),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3202),
.B(n_2829),
.Y(n_3416)
);

INVxp33_ASAP7_75t_SL g3417 ( 
.A(n_2948),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_2933),
.B(n_2656),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3202),
.B(n_2656),
.Y(n_3419)
);

INVxp33_ASAP7_75t_L g3420 ( 
.A(n_3057),
.Y(n_3420)
);

INVx2_ASAP7_75t_SL g3421 ( 
.A(n_2975),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_2907),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3042),
.B(n_2656),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_SL g3424 ( 
.A(n_3005),
.B(n_2838),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3184),
.B(n_2670),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3184),
.B(n_2670),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_2983),
.Y(n_3427)
);

OR2x6_ASAP7_75t_L g3428 ( 
.A(n_3241),
.B(n_2726),
.Y(n_3428)
);

NOR2xp33_ASAP7_75t_L g3429 ( 
.A(n_3059),
.B(n_2763),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_SL g3430 ( 
.A(n_2934),
.B(n_2842),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_SL g3431 ( 
.A(n_2941),
.B(n_2842),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_SL g3432 ( 
.A(n_2964),
.B(n_2845),
.Y(n_3432)
);

NOR2x2_ASAP7_75t_L g3433 ( 
.A(n_3223),
.B(n_2577),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_L g3434 ( 
.A(n_3059),
.B(n_2763),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_3131),
.B(n_2763),
.Y(n_3435)
);

NOR2xp67_ASAP7_75t_L g3436 ( 
.A(n_3120),
.B(n_2846),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_SL g3437 ( 
.A(n_2892),
.B(n_2846),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3188),
.B(n_2984),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_3188),
.B(n_3124),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_2908),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_2991),
.Y(n_3441)
);

AND2x4_ASAP7_75t_L g3442 ( 
.A(n_2900),
.B(n_2763),
.Y(n_3442)
);

NOR2xp33_ASAP7_75t_L g3443 ( 
.A(n_2990),
.B(n_2849),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3075),
.B(n_2670),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3075),
.B(n_2676),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3090),
.B(n_3024),
.Y(n_3446)
);

INVx3_ASAP7_75t_L g3447 ( 
.A(n_3019),
.Y(n_3447)
);

HB1xp67_ASAP7_75t_L g3448 ( 
.A(n_2888),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_2994),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_2909),
.Y(n_3450)
);

AND2x2_ASAP7_75t_L g3451 ( 
.A(n_3283),
.B(n_1933),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_2910),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_SL g3453 ( 
.A(n_2892),
.B(n_2849),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_2911),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3014),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_3093),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3090),
.B(n_2676),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_SL g3458 ( 
.A(n_2965),
.B(n_2851),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_2915),
.Y(n_3459)
);

BUFx6f_ASAP7_75t_L g3460 ( 
.A(n_3197),
.Y(n_3460)
);

INVx8_ASAP7_75t_L g3461 ( 
.A(n_3241),
.Y(n_3461)
);

OAI22xp5_ASAP7_75t_L g3462 ( 
.A1(n_2893),
.A2(n_2807),
.B1(n_2836),
.B2(n_2804),
.Y(n_3462)
);

NOR2xp33_ASAP7_75t_L g3463 ( 
.A(n_3266),
.B(n_2851),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3025),
.B(n_3026),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_SL g3465 ( 
.A(n_3015),
.B(n_2855),
.Y(n_3465)
);

NOR2xp67_ASAP7_75t_L g3466 ( 
.A(n_3120),
.B(n_2855),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_2893),
.B(n_2676),
.Y(n_3467)
);

AOI22xp5_ASAP7_75t_L g3468 ( 
.A1(n_3272),
.A2(n_2499),
.B1(n_2834),
.B2(n_2795),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3210),
.B(n_2814),
.Y(n_3469)
);

AND2x2_ASAP7_75t_L g3470 ( 
.A(n_3242),
.B(n_1836),
.Y(n_3470)
);

INVx2_ASAP7_75t_L g3471 ( 
.A(n_3102),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3210),
.B(n_2817),
.Y(n_3472)
);

OAI21xp5_ASAP7_75t_L g3473 ( 
.A1(n_3055),
.A2(n_2807),
.B(n_2804),
.Y(n_3473)
);

INVxp67_ASAP7_75t_L g3474 ( 
.A(n_3219),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_SL g3475 ( 
.A(n_2884),
.B(n_2575),
.Y(n_3475)
);

AO221x1_ASAP7_75t_L g3476 ( 
.A1(n_3079),
.A2(n_2748),
.B1(n_2777),
.B2(n_2738),
.C(n_2692),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3276),
.B(n_2817),
.Y(n_3477)
);

AOI22xp5_ASAP7_75t_L g3478 ( 
.A1(n_3277),
.A2(n_2499),
.B1(n_2834),
.B2(n_2795),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_SL g3479 ( 
.A(n_2884),
.B(n_2575),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_SL g3480 ( 
.A(n_2913),
.B(n_2931),
.Y(n_3480)
);

OR2x2_ASAP7_75t_L g3481 ( 
.A(n_3045),
.B(n_2688),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3276),
.B(n_2822),
.Y(n_3482)
);

AOI21xp5_ASAP7_75t_L g3483 ( 
.A1(n_3044),
.A2(n_2708),
.B(n_2592),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3106),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_2917),
.Y(n_3485)
);

AOI22xp5_ASAP7_75t_L g3486 ( 
.A1(n_3165),
.A2(n_2852),
.B1(n_2750),
.B2(n_2561),
.Y(n_3486)
);

O2A1O1Ixp33_ASAP7_75t_L g3487 ( 
.A1(n_3049),
.A2(n_1728),
.B(n_2852),
.C(n_1064),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_2918),
.Y(n_3488)
);

NOR3xp33_ASAP7_75t_L g3489 ( 
.A(n_3157),
.B(n_2833),
.C(n_2831),
.Y(n_3489)
);

INVx8_ASAP7_75t_L g3490 ( 
.A(n_3241),
.Y(n_3490)
);

OAI22xp33_ASAP7_75t_L g3491 ( 
.A1(n_3013),
.A2(n_2577),
.B1(n_2708),
.B2(n_2592),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_2924),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3107),
.Y(n_3493)
);

INVx2_ASAP7_75t_L g3494 ( 
.A(n_3117),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3028),
.B(n_3030),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_3128),
.Y(n_3496)
);

INVx2_ASAP7_75t_L g3497 ( 
.A(n_3159),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3031),
.B(n_2822),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_SL g3499 ( 
.A(n_2913),
.B(n_2593),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3260),
.B(n_2823),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_SL g3501 ( 
.A(n_2913),
.B(n_2593),
.Y(n_3501)
);

NOR2xp33_ASAP7_75t_L g3502 ( 
.A(n_3304),
.B(n_2800),
.Y(n_3502)
);

INVx8_ASAP7_75t_L g3503 ( 
.A(n_2979),
.Y(n_3503)
);

NOR2xp33_ASAP7_75t_L g3504 ( 
.A(n_3307),
.B(n_2800),
.Y(n_3504)
);

NOR2xp33_ASAP7_75t_L g3505 ( 
.A(n_3101),
.B(n_2800),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3261),
.B(n_2823),
.Y(n_3506)
);

INVx8_ASAP7_75t_L g3507 ( 
.A(n_2979),
.Y(n_3507)
);

INVx2_ASAP7_75t_L g3508 ( 
.A(n_3167),
.Y(n_3508)
);

CKINVDCx20_ASAP7_75t_R g3509 ( 
.A(n_2904),
.Y(n_3509)
);

BUFx3_ASAP7_75t_L g3510 ( 
.A(n_2931),
.Y(n_3510)
);

BUFx3_ASAP7_75t_L g3511 ( 
.A(n_2931),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3245),
.B(n_1836),
.Y(n_3512)
);

INVx2_ASAP7_75t_SL g3513 ( 
.A(n_2987),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3094),
.B(n_2835),
.Y(n_3514)
);

CKINVDCx11_ASAP7_75t_R g3515 ( 
.A(n_2905),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_SL g3516 ( 
.A(n_3275),
.B(n_2593),
.Y(n_3516)
);

BUFx6f_ASAP7_75t_SL g3517 ( 
.A(n_3297),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_2928),
.Y(n_3518)
);

AND2x6_ASAP7_75t_SL g3519 ( 
.A(n_3297),
.B(n_2783),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_2953),
.Y(n_3520)
);

CKINVDCx5p33_ASAP7_75t_R g3521 ( 
.A(n_3056),
.Y(n_3521)
);

NOR2xp33_ASAP7_75t_L g3522 ( 
.A(n_3157),
.B(n_2805),
.Y(n_3522)
);

NOR2xp33_ASAP7_75t_L g3523 ( 
.A(n_3171),
.B(n_2805),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_SL g3524 ( 
.A(n_3010),
.B(n_2593),
.Y(n_3524)
);

INVxp67_ASAP7_75t_L g3525 ( 
.A(n_3051),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_2929),
.Y(n_3526)
);

BUFx6f_ASAP7_75t_L g3527 ( 
.A(n_3197),
.Y(n_3527)
);

NOR2xp33_ASAP7_75t_L g3528 ( 
.A(n_3171),
.B(n_2805),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3094),
.B(n_2835),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3186),
.B(n_2828),
.Y(n_3530)
);

AND2x4_ASAP7_75t_L g3531 ( 
.A(n_2900),
.B(n_2688),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_2959),
.Y(n_3532)
);

AOI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_3189),
.A2(n_2561),
.B1(n_2872),
.B2(n_2864),
.Y(n_3533)
);

HB1xp67_ASAP7_75t_L g3534 ( 
.A(n_3221),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3190),
.B(n_2828),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_SL g3536 ( 
.A(n_3010),
.B(n_2593),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3130),
.B(n_2836),
.Y(n_3537)
);

AOI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_3156),
.A2(n_2561),
.B1(n_2877),
.B2(n_2850),
.Y(n_3538)
);

OR2x6_ASAP7_75t_L g3539 ( 
.A(n_3223),
.B(n_2592),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_SL g3540 ( 
.A(n_3116),
.B(n_2596),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3191),
.B(n_2830),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_2960),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3130),
.B(n_2828),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3192),
.B(n_2830),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_SL g3545 ( 
.A(n_3013),
.B(n_2596),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3193),
.B(n_2830),
.Y(n_3546)
);

INVx2_ASAP7_75t_L g3547 ( 
.A(n_2961),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_SL g3548 ( 
.A(n_3244),
.B(n_2596),
.Y(n_3548)
);

AOI22xp5_ASAP7_75t_L g3549 ( 
.A1(n_3156),
.A2(n_2825),
.B1(n_2721),
.B2(n_2741),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_2930),
.Y(n_3550)
);

INVx2_ASAP7_75t_SL g3551 ( 
.A(n_3225),
.Y(n_3551)
);

OAI22xp5_ASAP7_75t_L g3552 ( 
.A1(n_3296),
.A2(n_3183),
.B1(n_3182),
.B2(n_3194),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3195),
.B(n_2573),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3201),
.B(n_2573),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3205),
.B(n_2578),
.Y(n_3555)
);

AND2x6_ASAP7_75t_L g3556 ( 
.A(n_3153),
.B(n_2696),
.Y(n_3556)
);

OR2x6_ASAP7_75t_L g3557 ( 
.A(n_3223),
.B(n_2708),
.Y(n_3557)
);

INVx2_ASAP7_75t_L g3558 ( 
.A(n_2963),
.Y(n_3558)
);

NOR2xp33_ASAP7_75t_L g3559 ( 
.A(n_3224),
.B(n_2825),
.Y(n_3559)
);

NOR2xp33_ASAP7_75t_L g3560 ( 
.A(n_3224),
.B(n_2825),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_2966),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_2970),
.Y(n_3562)
);

INVx2_ASAP7_75t_L g3563 ( 
.A(n_2971),
.Y(n_3563)
);

OAI22xp5_ASAP7_75t_L g3564 ( 
.A1(n_3296),
.A2(n_2708),
.B1(n_2741),
.B2(n_2721),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3207),
.B(n_2578),
.Y(n_3565)
);

NOR2xp33_ASAP7_75t_SL g3566 ( 
.A(n_3071),
.B(n_2246),
.Y(n_3566)
);

OAI22xp33_ASAP7_75t_L g3567 ( 
.A1(n_2923),
.A2(n_2741),
.B1(n_2799),
.B2(n_2721),
.Y(n_3567)
);

NOR2xp33_ASAP7_75t_L g3568 ( 
.A(n_3181),
.B(n_2746),
.Y(n_3568)
);

AOI21xp5_ASAP7_75t_L g3569 ( 
.A1(n_3044),
.A2(n_2741),
.B(n_2721),
.Y(n_3569)
);

OAI22xp5_ASAP7_75t_SL g3570 ( 
.A1(n_3231),
.A2(n_1017),
.B1(n_1030),
.B2(n_1005),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3208),
.B(n_2578),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_2974),
.Y(n_3572)
);

OR2x2_ASAP7_75t_L g3573 ( 
.A(n_3218),
.B(n_3187),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3209),
.B(n_2579),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_2932),
.Y(n_3575)
);

BUFx3_ASAP7_75t_L g3576 ( 
.A(n_2919),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_2976),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3153),
.B(n_2579),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_2935),
.Y(n_3579)
);

NOR2xp33_ASAP7_75t_L g3580 ( 
.A(n_3170),
.B(n_2746),
.Y(n_3580)
);

INVxp67_ASAP7_75t_L g3581 ( 
.A(n_3227),
.Y(n_3581)
);

OR2x2_ASAP7_75t_L g3582 ( 
.A(n_3229),
.B(n_2696),
.Y(n_3582)
);

OR2x2_ASAP7_75t_L g3583 ( 
.A(n_3232),
.B(n_2702),
.Y(n_3583)
);

NOR3x1_ASAP7_75t_L g3584 ( 
.A(n_3085),
.B(n_3234),
.C(n_3233),
.Y(n_3584)
);

AOI22xp5_ASAP7_75t_L g3585 ( 
.A1(n_2923),
.A2(n_2799),
.B1(n_2861),
.B2(n_2857),
.Y(n_3585)
);

BUFx2_ASAP7_75t_L g3586 ( 
.A(n_3243),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_2936),
.B(n_2579),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_2937),
.B(n_2608),
.Y(n_3588)
);

NAND3xp33_ASAP7_75t_L g3589 ( 
.A(n_3235),
.B(n_3246),
.C(n_3238),
.Y(n_3589)
);

BUFx6f_ASAP7_75t_L g3590 ( 
.A(n_3197),
.Y(n_3590)
);

NOR2xp33_ASAP7_75t_L g3591 ( 
.A(n_2962),
.B(n_2692),
.Y(n_3591)
);

AOI22xp33_ASAP7_75t_L g3592 ( 
.A1(n_3038),
.A2(n_2702),
.B1(n_2706),
.B2(n_2704),
.Y(n_3592)
);

INVx2_ASAP7_75t_L g3593 ( 
.A(n_2977),
.Y(n_3593)
);

BUFx8_ASAP7_75t_L g3594 ( 
.A(n_2920),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_SL g3595 ( 
.A(n_3151),
.B(n_2596),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_2978),
.Y(n_3596)
);

O2A1O1Ixp33_ASAP7_75t_L g3597 ( 
.A1(n_3213),
.A2(n_1728),
.B(n_1064),
.C(n_1065),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3214),
.B(n_3215),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_2938),
.Y(n_3599)
);

AOI22xp33_ASAP7_75t_L g3600 ( 
.A1(n_3133),
.A2(n_3135),
.B1(n_3217),
.B2(n_3257),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_2940),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3262),
.B(n_2608),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3263),
.B(n_2608),
.Y(n_3603)
);

NAND2xp33_ASAP7_75t_L g3604 ( 
.A(n_2979),
.B(n_2799),
.Y(n_3604)
);

INVx4_ASAP7_75t_L g3605 ( 
.A(n_3226),
.Y(n_3605)
);

INVxp67_ASAP7_75t_L g3606 ( 
.A(n_3253),
.Y(n_3606)
);

NOR2xp33_ASAP7_75t_L g3607 ( 
.A(n_3204),
.B(n_3216),
.Y(n_3607)
);

NOR2xp33_ASAP7_75t_SL g3608 ( 
.A(n_3084),
.B(n_2560),
.Y(n_3608)
);

INVx2_ASAP7_75t_L g3609 ( 
.A(n_2985),
.Y(n_3609)
);

NOR2xp67_ASAP7_75t_L g3610 ( 
.A(n_3007),
.B(n_2704),
.Y(n_3610)
);

AOI22xp33_ASAP7_75t_L g3611 ( 
.A1(n_3264),
.A2(n_2706),
.B1(n_2716),
.B2(n_2707),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_2986),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_SL g3613 ( 
.A(n_3122),
.B(n_2596),
.Y(n_3613)
);

CKINVDCx5p33_ASAP7_75t_R g3614 ( 
.A(n_2927),
.Y(n_3614)
);

INVx5_ASAP7_75t_L g3615 ( 
.A(n_2979),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_L g3616 ( 
.A(n_3265),
.B(n_2707),
.Y(n_3616)
);

OR2x2_ASAP7_75t_L g3617 ( 
.A(n_3254),
.B(n_2716),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3269),
.B(n_2724),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3270),
.B(n_2724),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_2988),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3273),
.B(n_2729),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3274),
.B(n_2729),
.Y(n_3622)
);

INVxp67_ASAP7_75t_L g3623 ( 
.A(n_3255),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_2942),
.Y(n_3624)
);

NOR2xp33_ASAP7_75t_L g3625 ( 
.A(n_3252),
.B(n_2738),
.Y(n_3625)
);

NAND3xp33_ASAP7_75t_L g3626 ( 
.A(n_2939),
.B(n_1917),
.C(n_1914),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_2943),
.Y(n_3627)
);

NOR2xp33_ASAP7_75t_L g3628 ( 
.A(n_3009),
.B(n_2738),
.Y(n_3628)
);

BUFx6f_ASAP7_75t_L g3629 ( 
.A(n_3226),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3281),
.B(n_2731),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_2945),
.Y(n_3631)
);

INVxp67_ASAP7_75t_SL g3632 ( 
.A(n_3054),
.Y(n_3632)
);

HB1xp67_ASAP7_75t_SL g3633 ( 
.A(n_2919),
.Y(n_3633)
);

OR2x2_ASAP7_75t_SL g3634 ( 
.A(n_3158),
.B(n_1063),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_2949),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_2951),
.Y(n_3636)
);

OR2x2_ASAP7_75t_L g3637 ( 
.A(n_3032),
.B(n_2731),
.Y(n_3637)
);

NOR3xp33_ASAP7_75t_L g3638 ( 
.A(n_2972),
.B(n_1973),
.C(n_990),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_SL g3639 ( 
.A(n_3250),
.B(n_2628),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_2952),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_3282),
.B(n_3284),
.Y(n_3641)
);

AOI221xp5_ASAP7_75t_L g3642 ( 
.A1(n_3285),
.A2(n_995),
.B1(n_999),
.B2(n_992),
.C(n_989),
.Y(n_3642)
);

AND2x2_ASAP7_75t_L g3643 ( 
.A(n_3250),
.B(n_1847),
.Y(n_3643)
);

NOR2xp33_ASAP7_75t_L g3644 ( 
.A(n_2950),
.B(n_2748),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3286),
.B(n_2732),
.Y(n_3645)
);

AND2x4_ASAP7_75t_L g3646 ( 
.A(n_3096),
.B(n_2732),
.Y(n_3646)
);

AOI22xp5_ASAP7_75t_L g3647 ( 
.A1(n_2939),
.A2(n_2799),
.B1(n_2861),
.B2(n_2857),
.Y(n_3647)
);

INVx2_ASAP7_75t_SL g3648 ( 
.A(n_3096),
.Y(n_3648)
);

NOR2xp33_ASAP7_75t_L g3649 ( 
.A(n_2958),
.B(n_2748),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_SL g3650 ( 
.A(n_3161),
.B(n_2628),
.Y(n_3650)
);

OR2x2_ASAP7_75t_L g3651 ( 
.A(n_3290),
.B(n_2743),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3258),
.Y(n_3652)
);

NOR2xp33_ASAP7_75t_R g3653 ( 
.A(n_3249),
.B(n_2560),
.Y(n_3653)
);

NOR3xp33_ASAP7_75t_L g3654 ( 
.A(n_3136),
.B(n_1003),
.C(n_1002),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_3291),
.B(n_2743),
.Y(n_3655)
);

NOR2xp33_ASAP7_75t_L g3656 ( 
.A(n_3200),
.B(n_2777),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3259),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3294),
.B(n_2744),
.Y(n_3658)
);

AOI22xp33_ASAP7_75t_L g3659 ( 
.A1(n_3295),
.A2(n_2744),
.B1(n_2756),
.B2(n_2754),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_2989),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_2992),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_2993),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3298),
.B(n_2754),
.Y(n_3663)
);

AOI22xp33_ASAP7_75t_L g3664 ( 
.A1(n_3033),
.A2(n_2756),
.B1(n_2762),
.B2(n_2758),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3034),
.B(n_2801),
.Y(n_3665)
);

BUFx4f_ASAP7_75t_L g3666 ( 
.A(n_3297),
.Y(n_3666)
);

INVx4_ASAP7_75t_L g3667 ( 
.A(n_3226),
.Y(n_3667)
);

BUFx3_ASAP7_75t_L g3668 ( 
.A(n_2957),
.Y(n_3668)
);

NOR2xp33_ASAP7_75t_L g3669 ( 
.A(n_2982),
.B(n_2777),
.Y(n_3669)
);

AO22x1_ASAP7_75t_L g3670 ( 
.A1(n_3287),
.A2(n_1917),
.B1(n_1914),
.B2(n_1008),
.Y(n_3670)
);

AOI22xp33_ASAP7_75t_L g3671 ( 
.A1(n_3035),
.A2(n_2758),
.B1(n_2768),
.B2(n_2762),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_2996),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3037),
.B(n_2768),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_SL g3674 ( 
.A(n_3161),
.B(n_2628),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3039),
.B(n_2769),
.Y(n_3675)
);

INVx2_ASAP7_75t_SL g3676 ( 
.A(n_3198),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_2997),
.Y(n_3677)
);

A2O1A1Ixp33_ASAP7_75t_L g3678 ( 
.A1(n_3289),
.A2(n_2773),
.B(n_2774),
.C(n_2769),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3043),
.B(n_3046),
.Y(n_3679)
);

AOI22xp33_ASAP7_75t_L g3680 ( 
.A1(n_3047),
.A2(n_2773),
.B1(n_2780),
.B2(n_2774),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3000),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3054),
.B(n_2780),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_SL g3683 ( 
.A(n_3237),
.B(n_2628),
.Y(n_3683)
);

A2O1A1Ixp33_ASAP7_75t_L g3684 ( 
.A1(n_3289),
.A2(n_2791),
.B(n_2801),
.C(n_2790),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_SL g3685 ( 
.A(n_3237),
.B(n_2628),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_SL g3686 ( 
.A(n_3292),
.B(n_2677),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3002),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_SL g3688 ( 
.A(n_3292),
.B(n_2677),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3177),
.B(n_3180),
.Y(n_3689)
);

NAND2xp33_ASAP7_75t_L g3690 ( 
.A(n_2979),
.B(n_2677),
.Y(n_3690)
);

INVx3_ASAP7_75t_L g3691 ( 
.A(n_3267),
.Y(n_3691)
);

NOR2xp33_ASAP7_75t_L g3692 ( 
.A(n_3078),
.B(n_2786),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3006),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_SL g3694 ( 
.A(n_3299),
.B(n_2677),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3177),
.B(n_2790),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_L g3696 ( 
.A(n_3180),
.B(n_2791),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3008),
.Y(n_3697)
);

INVx2_ASAP7_75t_SL g3698 ( 
.A(n_3104),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3212),
.B(n_2786),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3011),
.Y(n_3700)
);

NOR2xp33_ASAP7_75t_L g3701 ( 
.A(n_3142),
.B(n_2786),
.Y(n_3701)
);

NOR2xp33_ASAP7_75t_L g3702 ( 
.A(n_3248),
.B(n_2787),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3212),
.B(n_2787),
.Y(n_3703)
);

AND2x2_ASAP7_75t_L g3704 ( 
.A(n_3074),
.B(n_1847),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3012),
.Y(n_3705)
);

AND2x4_ASAP7_75t_L g3706 ( 
.A(n_3077),
.B(n_2793),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3016),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3247),
.B(n_2787),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3247),
.B(n_2793),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3017),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3299),
.B(n_2793),
.Y(n_3711)
);

NAND2xp33_ASAP7_75t_SL g3712 ( 
.A(n_2920),
.B(n_2677),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3018),
.Y(n_3713)
);

CKINVDCx5p33_ASAP7_75t_R g3714 ( 
.A(n_3058),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_SL g3715 ( 
.A(n_3309),
.B(n_3077),
.Y(n_3715)
);

NOR2xp33_ASAP7_75t_L g3716 ( 
.A(n_3027),
.B(n_2794),
.Y(n_3716)
);

AOI21xp5_ASAP7_75t_L g3717 ( 
.A1(n_3398),
.A2(n_3055),
.B(n_3154),
.Y(n_3717)
);

AOI21xp5_ASAP7_75t_L g3718 ( 
.A1(n_3407),
.A2(n_3690),
.B(n_3320),
.Y(n_3718)
);

NOR2xp33_ASAP7_75t_L g3719 ( 
.A(n_3321),
.B(n_3166),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3331),
.A2(n_3160),
.B(n_3309),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3331),
.B(n_3023),
.Y(n_3721)
);

BUFx6f_ASAP7_75t_L g3722 ( 
.A(n_3461),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3319),
.B(n_3048),
.Y(n_3723)
);

AOI21xp5_ASAP7_75t_L g3724 ( 
.A1(n_3604),
.A2(n_3160),
.B(n_2583),
.Y(n_3724)
);

INVx6_ASAP7_75t_L g3725 ( 
.A(n_3594),
.Y(n_3725)
);

O2A1O1Ixp33_ASAP7_75t_L g3726 ( 
.A1(n_3341),
.A2(n_3040),
.B(n_3036),
.C(n_1065),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3319),
.B(n_3050),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_SL g3728 ( 
.A(n_3360),
.B(n_3369),
.Y(n_3728)
);

AND2x2_ASAP7_75t_SL g3729 ( 
.A(n_3666),
.B(n_3211),
.Y(n_3729)
);

INVxp67_ASAP7_75t_L g3730 ( 
.A(n_3316),
.Y(n_3730)
);

AO21x1_ASAP7_75t_L g3731 ( 
.A1(n_3357),
.A2(n_3040),
.B(n_3036),
.Y(n_3731)
);

AOI21xp5_ASAP7_75t_L g3732 ( 
.A1(n_3469),
.A2(n_2583),
.B(n_2522),
.Y(n_3732)
);

INVx3_ASAP7_75t_L g3733 ( 
.A(n_3706),
.Y(n_3733)
);

AOI22xp5_ASAP7_75t_L g3734 ( 
.A1(n_3568),
.A2(n_3067),
.B1(n_3058),
.B2(n_3052),
.Y(n_3734)
);

AOI21xp5_ASAP7_75t_L g3735 ( 
.A1(n_3469),
.A2(n_2583),
.B(n_2522),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_SL g3736 ( 
.A(n_3378),
.B(n_3077),
.Y(n_3736)
);

BUFx6f_ASAP7_75t_L g3737 ( 
.A(n_3461),
.Y(n_3737)
);

AOI21xp5_ASAP7_75t_L g3738 ( 
.A1(n_3472),
.A2(n_2610),
.B(n_2522),
.Y(n_3738)
);

AND2x2_ASAP7_75t_L g3739 ( 
.A(n_3324),
.B(n_3315),
.Y(n_3739)
);

O2A1O1Ixp33_ASAP7_75t_L g3740 ( 
.A1(n_3354),
.A2(n_1066),
.B(n_1091),
.C(n_1063),
.Y(n_3740)
);

NOR3xp33_ASAP7_75t_L g3741 ( 
.A(n_3334),
.B(n_1091),
.C(n_1066),
.Y(n_3741)
);

A2O1A1Ixp33_ASAP7_75t_L g3742 ( 
.A1(n_3580),
.A2(n_3312),
.B(n_3053),
.C(n_3062),
.Y(n_3742)
);

A2O1A1Ixp33_ASAP7_75t_L g3743 ( 
.A1(n_3438),
.A2(n_3312),
.B(n_3061),
.C(n_3064),
.Y(n_3743)
);

INVxp67_ASAP7_75t_SL g3744 ( 
.A(n_3689),
.Y(n_3744)
);

NOR2xp33_ASAP7_75t_L g3745 ( 
.A(n_3439),
.B(n_3306),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_SL g3746 ( 
.A(n_3323),
.B(n_3168),
.Y(n_3746)
);

AOI21xp5_ASAP7_75t_L g3747 ( 
.A1(n_3472),
.A2(n_2672),
.B(n_2610),
.Y(n_3747)
);

AOI21xp5_ASAP7_75t_L g3748 ( 
.A1(n_3477),
.A2(n_2672),
.B(n_2610),
.Y(n_3748)
);

NOR2x1_ASAP7_75t_L g3749 ( 
.A(n_3415),
.B(n_3301),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3326),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3332),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_SL g3752 ( 
.A(n_3340),
.B(n_3168),
.Y(n_3752)
);

BUFx6f_ASAP7_75t_L g3753 ( 
.A(n_3461),
.Y(n_3753)
);

INVx2_ASAP7_75t_SL g3754 ( 
.A(n_3375),
.Y(n_3754)
);

CKINVDCx6p67_ASAP7_75t_R g3755 ( 
.A(n_3515),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3333),
.B(n_3063),
.Y(n_3756)
);

OAI21x1_ASAP7_75t_L g3757 ( 
.A1(n_3483),
.A2(n_3103),
.B(n_3066),
.Y(n_3757)
);

BUFx6f_ASAP7_75t_L g3758 ( 
.A(n_3490),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3361),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3333),
.B(n_3068),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3362),
.Y(n_3761)
);

A2O1A1Ixp33_ASAP7_75t_L g3762 ( 
.A1(n_3322),
.A2(n_3069),
.B(n_3072),
.C(n_3070),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_3355),
.B(n_3073),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_3376),
.B(n_3076),
.Y(n_3764)
);

INVx2_ASAP7_75t_L g3765 ( 
.A(n_3582),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_3470),
.B(n_3080),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3443),
.B(n_3082),
.Y(n_3767)
);

AOI21xp5_ASAP7_75t_L g3768 ( 
.A1(n_3477),
.A2(n_2718),
.B(n_2672),
.Y(n_3768)
);

AOI22xp33_ASAP7_75t_L g3769 ( 
.A1(n_3607),
.A2(n_3067),
.B1(n_3236),
.B2(n_3199),
.Y(n_3769)
);

AOI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_3482),
.A2(n_2728),
.B(n_2718),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3583),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3365),
.Y(n_3772)
);

OAI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3364),
.A2(n_3368),
.B(n_3372),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3328),
.B(n_3083),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3328),
.B(n_3087),
.Y(n_3775)
);

AOI21xp5_ASAP7_75t_L g3776 ( 
.A1(n_3482),
.A2(n_3347),
.B(n_3344),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3397),
.B(n_3088),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3377),
.Y(n_3778)
);

NAND3xp33_ASAP7_75t_L g3779 ( 
.A(n_3395),
.B(n_1011),
.C(n_1007),
.Y(n_3779)
);

NOR3xp33_ASAP7_75t_L g3780 ( 
.A(n_3626),
.B(n_1113),
.C(n_1112),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3446),
.B(n_3089),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3344),
.A2(n_2728),
.B(n_2718),
.Y(n_3782)
);

NAND2x1_ASAP7_75t_L g3783 ( 
.A(n_3706),
.B(n_2691),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3385),
.B(n_3091),
.Y(n_3784)
);

AOI21xp5_ASAP7_75t_L g3785 ( 
.A1(n_3347),
.A2(n_3473),
.B(n_3445),
.Y(n_3785)
);

BUFx6f_ASAP7_75t_L g3786 ( 
.A(n_3490),
.Y(n_3786)
);

INVx3_ASAP7_75t_L g3787 ( 
.A(n_3539),
.Y(n_3787)
);

AOI21xp5_ASAP7_75t_L g3788 ( 
.A1(n_3473),
.A2(n_2728),
.B(n_2691),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3384),
.Y(n_3789)
);

AND2x4_ASAP7_75t_L g3790 ( 
.A(n_3442),
.B(n_3168),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3390),
.B(n_3092),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3451),
.B(n_3095),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3416),
.B(n_3097),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3393),
.Y(n_3794)
);

AOI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3444),
.A2(n_2770),
.B(n_2691),
.Y(n_3795)
);

BUFx2_ASAP7_75t_L g3796 ( 
.A(n_3386),
.Y(n_3796)
);

AND2x4_ASAP7_75t_L g3797 ( 
.A(n_3442),
.B(n_3196),
.Y(n_3797)
);

AOI21xp5_ASAP7_75t_L g3798 ( 
.A1(n_3457),
.A2(n_2770),
.B(n_2691),
.Y(n_3798)
);

OAI321xp33_ASAP7_75t_L g3799 ( 
.A1(n_3600),
.A2(n_1123),
.A3(n_1113),
.B1(n_1124),
.B2(n_1117),
.C(n_1112),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_SL g3800 ( 
.A(n_3405),
.B(n_3206),
.Y(n_3800)
);

INVx2_ASAP7_75t_SL g3801 ( 
.A(n_3330),
.Y(n_3801)
);

NOR2xp33_ASAP7_75t_SL g3802 ( 
.A(n_3521),
.B(n_3417),
.Y(n_3802)
);

AOI21xp5_ASAP7_75t_L g3803 ( 
.A1(n_3689),
.A2(n_2770),
.B(n_2691),
.Y(n_3803)
);

HB1xp67_ASAP7_75t_L g3804 ( 
.A(n_3352),
.Y(n_3804)
);

NOR2xp33_ASAP7_75t_L g3805 ( 
.A(n_3420),
.B(n_3098),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3409),
.B(n_3099),
.Y(n_3806)
);

OAI21xp5_ASAP7_75t_L g3807 ( 
.A1(n_3337),
.A2(n_3109),
.B(n_3100),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3350),
.B(n_3111),
.Y(n_3808)
);

NOR2xp33_ASAP7_75t_L g3809 ( 
.A(n_3573),
.B(n_3112),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3353),
.B(n_3113),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_SL g3811 ( 
.A(n_3329),
.B(n_3239),
.Y(n_3811)
);

HB1xp67_ASAP7_75t_L g3812 ( 
.A(n_3383),
.Y(n_3812)
);

AOI21xp5_ASAP7_75t_L g3813 ( 
.A1(n_3391),
.A2(n_2770),
.B(n_2516),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_SL g3814 ( 
.A(n_3513),
.B(n_3240),
.Y(n_3814)
);

BUFx3_ASAP7_75t_L g3815 ( 
.A(n_3370),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_3617),
.Y(n_3816)
);

NOR2xp33_ASAP7_75t_L g3817 ( 
.A(n_3637),
.B(n_3525),
.Y(n_3817)
);

INVx3_ASAP7_75t_L g3818 ( 
.A(n_3539),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3392),
.B(n_3402),
.Y(n_3819)
);

O2A1O1Ixp33_ASAP7_75t_L g3820 ( 
.A1(n_3437),
.A2(n_1123),
.B(n_1124),
.C(n_1117),
.Y(n_3820)
);

NOR3xp33_ASAP7_75t_L g3821 ( 
.A(n_3404),
.B(n_1129),
.C(n_1126),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_3569),
.A2(n_2770),
.B(n_2516),
.Y(n_3822)
);

O2A1O1Ixp33_ASAP7_75t_L g3823 ( 
.A1(n_3453),
.A2(n_1129),
.B(n_1130),
.C(n_1126),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3436),
.B(n_3114),
.Y(n_3824)
);

INVx2_ASAP7_75t_L g3825 ( 
.A(n_3651),
.Y(n_3825)
);

NOR2x1p5_ASAP7_75t_L g3826 ( 
.A(n_3668),
.B(n_3115),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_SL g3827 ( 
.A(n_3466),
.B(n_3279),
.Y(n_3827)
);

OAI21x1_ASAP7_75t_L g3828 ( 
.A1(n_3462),
.A2(n_3066),
.B(n_3041),
.Y(n_3828)
);

NAND2x1_ASAP7_75t_L g3829 ( 
.A(n_3605),
.B(n_3280),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3520),
.Y(n_3830)
);

INVx2_ASAP7_75t_L g3831 ( 
.A(n_3532),
.Y(n_3831)
);

NOR2xp33_ASAP7_75t_SL g3832 ( 
.A(n_3614),
.B(n_3288),
.Y(n_3832)
);

AND2x4_ASAP7_75t_L g3833 ( 
.A(n_3539),
.B(n_3302),
.Y(n_3833)
);

AND2x2_ASAP7_75t_SL g3834 ( 
.A(n_3666),
.B(n_1130),
.Y(n_3834)
);

OAI21xp5_ASAP7_75t_L g3835 ( 
.A1(n_3337),
.A2(n_3414),
.B(n_3339),
.Y(n_3835)
);

HB1xp67_ASAP7_75t_L g3836 ( 
.A(n_3421),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_3512),
.B(n_3118),
.Y(n_3837)
);

INVx4_ASAP7_75t_L g3838 ( 
.A(n_3490),
.Y(n_3838)
);

INVx1_ASAP7_75t_SL g3839 ( 
.A(n_3371),
.Y(n_3839)
);

OAI22xp5_ASAP7_75t_L g3840 ( 
.A1(n_3632),
.A2(n_3478),
.B1(n_3468),
.B2(n_3356),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3351),
.B(n_3119),
.Y(n_3841)
);

NOR2xp33_ASAP7_75t_L g3842 ( 
.A(n_3628),
.B(n_3123),
.Y(n_3842)
);

AOI22xp5_ASAP7_75t_L g3843 ( 
.A1(n_3552),
.A2(n_3126),
.B1(n_3129),
.B2(n_3127),
.Y(n_3843)
);

NOR2x1p5_ASAP7_75t_L g3844 ( 
.A(n_3576),
.B(n_3132),
.Y(n_3844)
);

AOI21xp5_ASAP7_75t_L g3845 ( 
.A1(n_3327),
.A2(n_2516),
.B(n_2462),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_3351),
.B(n_3134),
.Y(n_3846)
);

HB1xp67_ASAP7_75t_L g3847 ( 
.A(n_3374),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_SL g3848 ( 
.A(n_3342),
.B(n_3303),
.Y(n_3848)
);

AND2x4_ASAP7_75t_L g3849 ( 
.A(n_3557),
.B(n_3137),
.Y(n_3849)
);

BUFx6f_ASAP7_75t_L g3850 ( 
.A(n_3460),
.Y(n_3850)
);

AND2x4_ASAP7_75t_L g3851 ( 
.A(n_3557),
.B(n_3138),
.Y(n_3851)
);

AOI21xp5_ASAP7_75t_L g3852 ( 
.A1(n_3327),
.A2(n_3529),
.B(n_3514),
.Y(n_3852)
);

INVx3_ASAP7_75t_L g3853 ( 
.A(n_3557),
.Y(n_3853)
);

AOI21xp5_ASAP7_75t_L g3854 ( 
.A1(n_3514),
.A2(n_2516),
.B(n_2462),
.Y(n_3854)
);

AOI21xp5_ASAP7_75t_L g3855 ( 
.A1(n_3529),
.A2(n_2516),
.B(n_2462),
.Y(n_3855)
);

O2A1O1Ixp33_ASAP7_75t_L g3856 ( 
.A1(n_3336),
.A2(n_1134),
.B(n_1135),
.C(n_1131),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3463),
.B(n_3495),
.Y(n_3857)
);

AOI21xp5_ASAP7_75t_L g3858 ( 
.A1(n_3537),
.A2(n_2571),
.B(n_2462),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3495),
.B(n_3139),
.Y(n_3859)
);

O2A1O1Ixp33_ASAP7_75t_L g3860 ( 
.A1(n_3366),
.A2(n_1134),
.B(n_1135),
.C(n_1131),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3598),
.B(n_3140),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3403),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3410),
.Y(n_3863)
);

AOI21xp5_ASAP7_75t_L g3864 ( 
.A1(n_3537),
.A2(n_2571),
.B(n_2462),
.Y(n_3864)
);

CKINVDCx5p33_ASAP7_75t_R g3865 ( 
.A(n_3509),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3641),
.B(n_3141),
.Y(n_3866)
);

NOR2x1_ASAP7_75t_L g3867 ( 
.A(n_3415),
.B(n_3510),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_3358),
.B(n_3145),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3358),
.B(n_3147),
.Y(n_3869)
);

NOR2xp33_ASAP7_75t_L g3870 ( 
.A(n_3474),
.B(n_3148),
.Y(n_3870)
);

AOI21xp5_ASAP7_75t_L g3871 ( 
.A1(n_3359),
.A2(n_2820),
.B(n_2571),
.Y(n_3871)
);

AOI21xp33_ASAP7_75t_L g3872 ( 
.A1(n_3591),
.A2(n_3367),
.B(n_3363),
.Y(n_3872)
);

AOI21xp5_ASAP7_75t_L g3873 ( 
.A1(n_3359),
.A2(n_2820),
.B(n_2571),
.Y(n_3873)
);

OAI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_3338),
.A2(n_3339),
.B(n_3381),
.Y(n_3874)
);

O2A1O1Ixp5_ASAP7_75t_L g3875 ( 
.A1(n_3545),
.A2(n_3683),
.B(n_3685),
.C(n_3595),
.Y(n_3875)
);

AND2x2_ASAP7_75t_L g3876 ( 
.A(n_3704),
.B(n_3149),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3542),
.Y(n_3877)
);

AOI21xp5_ASAP7_75t_L g3878 ( 
.A1(n_3338),
.A2(n_3564),
.B(n_3467),
.Y(n_3878)
);

AOI21xp5_ASAP7_75t_L g3879 ( 
.A1(n_3564),
.A2(n_2820),
.B(n_2571),
.Y(n_3879)
);

INVx6_ASAP7_75t_L g3880 ( 
.A(n_3594),
.Y(n_3880)
);

AOI21x1_ASAP7_75t_L g3881 ( 
.A1(n_3419),
.A2(n_3041),
.B(n_2235),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3422),
.Y(n_3882)
);

AOI21xp5_ASAP7_75t_L g3883 ( 
.A1(n_3467),
.A2(n_2820),
.B(n_2867),
.Y(n_3883)
);

AOI22xp33_ASAP7_75t_L g3884 ( 
.A1(n_3656),
.A2(n_3152),
.B1(n_3155),
.B2(n_3150),
.Y(n_3884)
);

BUFx6f_ASAP7_75t_L g3885 ( 
.A(n_3460),
.Y(n_3885)
);

NAND2xp33_ASAP7_75t_L g3886 ( 
.A(n_3489),
.B(n_2916),
.Y(n_3886)
);

O2A1O1Ixp5_ASAP7_75t_L g3887 ( 
.A1(n_3400),
.A2(n_3162),
.B(n_3169),
.C(n_3164),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3440),
.Y(n_3888)
);

NOR2x1p5_ASAP7_75t_L g3889 ( 
.A(n_3714),
.B(n_3173),
.Y(n_3889)
);

INVx2_ASAP7_75t_L g3890 ( 
.A(n_3547),
.Y(n_3890)
);

OAI321xp33_ASAP7_75t_L g3891 ( 
.A1(n_3570),
.A2(n_1143),
.A3(n_1139),
.B1(n_1151),
.B2(n_1141),
.C(n_1138),
.Y(n_3891)
);

AOI22xp5_ASAP7_75t_L g3892 ( 
.A1(n_3552),
.A2(n_3174),
.B1(n_3176),
.B2(n_3175),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_SL g3893 ( 
.A(n_3610),
.B(n_3305),
.Y(n_3893)
);

AOI21xp33_ASAP7_75t_L g3894 ( 
.A1(n_3396),
.A2(n_3179),
.B(n_3178),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3450),
.Y(n_3895)
);

NOR2xp33_ASAP7_75t_L g3896 ( 
.A(n_3644),
.B(n_3310),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_3464),
.B(n_3311),
.Y(n_3897)
);

AND2x4_ASAP7_75t_L g3898 ( 
.A(n_3511),
.B(n_3313),
.Y(n_3898)
);

HB1xp67_ASAP7_75t_L g3899 ( 
.A(n_3448),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_SL g3900 ( 
.A(n_3649),
.B(n_2916),
.Y(n_3900)
);

INVx3_ASAP7_75t_L g3901 ( 
.A(n_3503),
.Y(n_3901)
);

AOI21xp33_ASAP7_75t_L g3902 ( 
.A1(n_3380),
.A2(n_2866),
.B(n_2862),
.Y(n_3902)
);

BUFx12f_ASAP7_75t_L g3903 ( 
.A(n_3519),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3317),
.B(n_2794),
.Y(n_3904)
);

AOI21xp5_ASAP7_75t_L g3905 ( 
.A1(n_3418),
.A2(n_2820),
.B(n_2867),
.Y(n_3905)
);

AOI22xp5_ASAP7_75t_L g3906 ( 
.A1(n_3335),
.A2(n_1777),
.B1(n_1013),
.B2(n_1014),
.Y(n_3906)
);

OAI22xp5_ASAP7_75t_L g3907 ( 
.A1(n_3549),
.A2(n_3003),
.B1(n_2550),
.B2(n_2761),
.Y(n_3907)
);

INVx1_ASAP7_75t_SL g3908 ( 
.A(n_3481),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3452),
.Y(n_3909)
);

O2A1O1Ixp5_ASAP7_75t_L g3910 ( 
.A1(n_3401),
.A2(n_2794),
.B(n_2792),
.C(n_2631),
.Y(n_3910)
);

AOI21xp5_ASAP7_75t_L g3911 ( 
.A1(n_3418),
.A2(n_2812),
.B(n_3003),
.Y(n_3911)
);

AOI21xp5_ASAP7_75t_L g3912 ( 
.A1(n_3711),
.A2(n_1783),
.B(n_1780),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_SL g3913 ( 
.A(n_3388),
.B(n_2843),
.Y(n_3913)
);

INVx3_ASAP7_75t_L g3914 ( 
.A(n_3503),
.Y(n_3914)
);

NOR2xp33_ASAP7_75t_L g3915 ( 
.A(n_3692),
.B(n_2862),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3454),
.Y(n_3916)
);

OAI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3425),
.A2(n_2868),
.B(n_2866),
.Y(n_3917)
);

BUFx2_ASAP7_75t_L g3918 ( 
.A(n_3435),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3581),
.B(n_2868),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3459),
.Y(n_3920)
);

OAI21xp5_ASAP7_75t_L g3921 ( 
.A1(n_3426),
.A2(n_2879),
.B(n_2876),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_SL g3922 ( 
.A(n_3669),
.B(n_2843),
.Y(n_3922)
);

HB1xp67_ASAP7_75t_L g3923 ( 
.A(n_3534),
.Y(n_3923)
);

BUFx4f_ASAP7_75t_L g3924 ( 
.A(n_3428),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_SL g3925 ( 
.A(n_3551),
.B(n_2878),
.Y(n_3925)
);

AOI21xp5_ASAP7_75t_L g3926 ( 
.A1(n_3615),
.A2(n_1783),
.B(n_1780),
.Y(n_3926)
);

BUFx12f_ASAP7_75t_L g3927 ( 
.A(n_3399),
.Y(n_3927)
);

AOI22xp5_ASAP7_75t_L g3928 ( 
.A1(n_3716),
.A2(n_1777),
.B1(n_1016),
.B2(n_1018),
.Y(n_3928)
);

AND2x2_ASAP7_75t_SL g3929 ( 
.A(n_3608),
.B(n_1138),
.Y(n_3929)
);

AND2x2_ASAP7_75t_L g3930 ( 
.A(n_3701),
.B(n_1515),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3606),
.B(n_2876),
.Y(n_3931)
);

BUFx6f_ASAP7_75t_L g3932 ( 
.A(n_3460),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3623),
.B(n_2879),
.Y(n_3933)
);

AOI21xp5_ASAP7_75t_L g3934 ( 
.A1(n_3615),
.A2(n_1783),
.B(n_1780),
.Y(n_3934)
);

AOI21xp5_ASAP7_75t_L g3935 ( 
.A1(n_3615),
.A2(n_1783),
.B(n_1780),
.Y(n_3935)
);

AOI21x1_ASAP7_75t_L g3936 ( 
.A1(n_3348),
.A2(n_2237),
.B(n_2230),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3485),
.Y(n_3937)
);

OAI21xp33_ASAP7_75t_L g3938 ( 
.A1(n_3642),
.A2(n_1021),
.B(n_1012),
.Y(n_3938)
);

INVx4_ASAP7_75t_L g3939 ( 
.A(n_3527),
.Y(n_3939)
);

INVx3_ASAP7_75t_L g3940 ( 
.A(n_3503),
.Y(n_3940)
);

AOI21xp5_ASAP7_75t_L g3941 ( 
.A1(n_3615),
.A2(n_1831),
.B(n_1806),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3488),
.Y(n_3942)
);

AOI21xp5_ASAP7_75t_L g3943 ( 
.A1(n_3543),
.A2(n_1831),
.B(n_1806),
.Y(n_3943)
);

BUFx3_ASAP7_75t_L g3944 ( 
.A(n_3586),
.Y(n_3944)
);

AOI21xp5_ASAP7_75t_L g3945 ( 
.A1(n_3543),
.A2(n_1831),
.B(n_1806),
.Y(n_3945)
);

OAI21xp5_ASAP7_75t_L g3946 ( 
.A1(n_3533),
.A2(n_2878),
.B(n_2240),
.Y(n_3946)
);

AND2x2_ASAP7_75t_L g3947 ( 
.A(n_3643),
.B(n_1516),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3387),
.B(n_2878),
.Y(n_3948)
);

AO21x1_ASAP7_75t_L g3949 ( 
.A1(n_3379),
.A2(n_2247),
.B(n_2238),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3389),
.B(n_1885),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_SL g3951 ( 
.A(n_3505),
.B(n_1022),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_SL g3952 ( 
.A(n_3531),
.B(n_1024),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3492),
.B(n_1885),
.Y(n_3953)
);

AOI22xp5_ASAP7_75t_L g3954 ( 
.A1(n_3412),
.A2(n_1777),
.B1(n_1027),
.B2(n_1029),
.Y(n_3954)
);

INVx2_ASAP7_75t_L g3955 ( 
.A(n_3558),
.Y(n_3955)
);

AOI21xp5_ASAP7_75t_L g3956 ( 
.A1(n_3462),
.A2(n_1806),
.B(n_1831),
.Y(n_3956)
);

INVx3_ASAP7_75t_L g3957 ( 
.A(n_3507),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3518),
.B(n_1907),
.Y(n_3958)
);

OAI22xp5_ASAP7_75t_L g3959 ( 
.A1(n_3585),
.A2(n_3647),
.B1(n_3589),
.B2(n_3526),
.Y(n_3959)
);

OAI22xp5_ASAP7_75t_L g3960 ( 
.A1(n_3550),
.A2(n_2299),
.B1(n_2125),
.B2(n_2152),
.Y(n_3960)
);

INVx1_ASAP7_75t_SL g3961 ( 
.A(n_3653),
.Y(n_3961)
);

AOI21xp5_ASAP7_75t_L g3962 ( 
.A1(n_3578),
.A2(n_2086),
.B(n_2083),
.Y(n_3962)
);

BUFx2_ASAP7_75t_L g3963 ( 
.A(n_3531),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3575),
.B(n_1907),
.Y(n_3964)
);

A2O1A1Ixp33_ASAP7_75t_L g3965 ( 
.A1(n_3382),
.A2(n_1141),
.B(n_1143),
.C(n_1139),
.Y(n_3965)
);

AOI21xp5_ASAP7_75t_L g3966 ( 
.A1(n_3578),
.A2(n_2086),
.B(n_2083),
.Y(n_3966)
);

AOI21xp5_ASAP7_75t_L g3967 ( 
.A1(n_3686),
.A2(n_2086),
.B(n_2083),
.Y(n_3967)
);

AOI21xp5_ASAP7_75t_L g3968 ( 
.A1(n_3688),
.A2(n_3694),
.B(n_3715),
.Y(n_3968)
);

AOI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3423),
.A2(n_3699),
.B(n_3703),
.Y(n_3969)
);

BUFx6f_ASAP7_75t_L g3970 ( 
.A(n_3527),
.Y(n_3970)
);

BUFx2_ASAP7_75t_L g3971 ( 
.A(n_3527),
.Y(n_3971)
);

OAI21xp5_ASAP7_75t_L g3972 ( 
.A1(n_3538),
.A2(n_3486),
.B(n_3348),
.Y(n_3972)
);

AOI21xp5_ASAP7_75t_L g3973 ( 
.A1(n_3699),
.A2(n_2096),
.B(n_2086),
.Y(n_3973)
);

AOI22xp33_ASAP7_75t_L g3974 ( 
.A1(n_3654),
.A2(n_1157),
.B1(n_1159),
.B2(n_1151),
.Y(n_3974)
);

AOI22xp5_ASAP7_75t_L g3975 ( 
.A1(n_3559),
.A2(n_1777),
.B1(n_1031),
.B2(n_1034),
.Y(n_3975)
);

O2A1O1Ixp33_ASAP7_75t_L g3976 ( 
.A1(n_3613),
.A2(n_1159),
.B(n_1162),
.C(n_1157),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3579),
.B(n_1943),
.Y(n_3977)
);

BUFx6f_ASAP7_75t_L g3978 ( 
.A(n_3590),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3599),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3601),
.Y(n_3980)
);

OAI22xp5_ASAP7_75t_L g3981 ( 
.A1(n_3624),
.A2(n_2299),
.B1(n_2125),
.B2(n_2152),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3627),
.Y(n_3982)
);

OAI21x1_ASAP7_75t_L g3983 ( 
.A1(n_3665),
.A2(n_2180),
.B(n_2110),
.Y(n_3983)
);

NOR2xp33_ASAP7_75t_SL g3984 ( 
.A(n_3566),
.B(n_1025),
.Y(n_3984)
);

AOI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3703),
.A2(n_2100),
.B(n_2096),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3631),
.B(n_1943),
.Y(n_3986)
);

CKINVDCx5p33_ASAP7_75t_R g3987 ( 
.A(n_3633),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3708),
.A2(n_2100),
.B(n_2096),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3635),
.B(n_2004),
.Y(n_3989)
);

INVx2_ASAP7_75t_L g3990 ( 
.A(n_3561),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_3636),
.B(n_2004),
.Y(n_3991)
);

AOI21xp5_ASAP7_75t_L g3992 ( 
.A1(n_3708),
.A2(n_2100),
.B(n_2096),
.Y(n_3992)
);

INVx3_ASAP7_75t_L g3993 ( 
.A(n_3507),
.Y(n_3993)
);

AOI21xp5_ASAP7_75t_L g3994 ( 
.A1(n_3567),
.A2(n_3695),
.B(n_3682),
.Y(n_3994)
);

AOI21x1_ASAP7_75t_L g3995 ( 
.A1(n_3424),
.A2(n_2258),
.B(n_2253),
.Y(n_3995)
);

AOI21xp5_ASAP7_75t_L g3996 ( 
.A1(n_3682),
.A2(n_2102),
.B(n_2100),
.Y(n_3996)
);

NOR3xp33_ASAP7_75t_L g3997 ( 
.A(n_3522),
.B(n_1172),
.C(n_1162),
.Y(n_3997)
);

AOI21xp5_ASAP7_75t_L g3998 ( 
.A1(n_3695),
.A2(n_2137),
.B(n_2102),
.Y(n_3998)
);

BUFx2_ASAP7_75t_L g3999 ( 
.A(n_3590),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3640),
.B(n_2005),
.Y(n_4000)
);

CKINVDCx8_ASAP7_75t_R g4001 ( 
.A(n_3428),
.Y(n_4001)
);

NOR2xp33_ASAP7_75t_L g4002 ( 
.A(n_3698),
.B(n_3676),
.Y(n_4002)
);

OAI22xp5_ASAP7_75t_L g4003 ( 
.A1(n_3652),
.A2(n_2190),
.B1(n_2203),
.B2(n_2180),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3562),
.Y(n_4004)
);

AOI21xp5_ASAP7_75t_L g4005 ( 
.A1(n_3696),
.A2(n_2137),
.B(n_2102),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3657),
.B(n_3430),
.Y(n_4006)
);

INVx2_ASAP7_75t_L g4007 ( 
.A(n_3563),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_3572),
.Y(n_4008)
);

OAI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_3431),
.A2(n_2261),
.B(n_2260),
.Y(n_4009)
);

HB1xp67_ASAP7_75t_L g4010 ( 
.A(n_3796),
.Y(n_4010)
);

OAI22xp5_ASAP7_75t_L g4011 ( 
.A1(n_3719),
.A2(n_3528),
.B1(n_3523),
.B2(n_3560),
.Y(n_4011)
);

INVxp33_ASAP7_75t_L g4012 ( 
.A(n_3817),
.Y(n_4012)
);

BUFx8_ASAP7_75t_SL g4013 ( 
.A(n_3865),
.Y(n_4013)
);

OAI22xp5_ASAP7_75t_L g4014 ( 
.A1(n_3728),
.A2(n_3434),
.B1(n_3429),
.B2(n_3502),
.Y(n_4014)
);

AOI22xp5_ASAP7_75t_L g4015 ( 
.A1(n_3745),
.A2(n_3734),
.B1(n_3809),
.B2(n_3834),
.Y(n_4015)
);

OAI22xp5_ASAP7_75t_L g4016 ( 
.A1(n_3744),
.A2(n_3702),
.B1(n_3491),
.B2(n_3540),
.Y(n_4016)
);

AOI22xp5_ASAP7_75t_L g4017 ( 
.A1(n_3734),
.A2(n_3638),
.B1(n_3504),
.B2(n_3648),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3857),
.B(n_3432),
.Y(n_4018)
);

AOI21xp5_ASAP7_75t_L g4019 ( 
.A1(n_3718),
.A2(n_3507),
.B(n_3696),
.Y(n_4019)
);

AOI21x1_ASAP7_75t_L g4020 ( 
.A1(n_3936),
.A2(n_3325),
.B(n_3411),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3739),
.B(n_3625),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3819),
.B(n_3465),
.Y(n_4022)
);

OA22x2_ASAP7_75t_L g4023 ( 
.A1(n_3908),
.A2(n_3730),
.B1(n_3899),
.B2(n_3923),
.Y(n_4023)
);

AOI21xp5_ASAP7_75t_L g4024 ( 
.A1(n_3720),
.A2(n_3709),
.B(n_3349),
.Y(n_4024)
);

OAI22xp5_ASAP7_75t_L g4025 ( 
.A1(n_3842),
.A2(n_3634),
.B1(n_3428),
.B2(n_3458),
.Y(n_4025)
);

BUFx2_ASAP7_75t_L g4026 ( 
.A(n_3804),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_3830),
.Y(n_4027)
);

NAND2x1_ASAP7_75t_L g4028 ( 
.A(n_3787),
.B(n_3556),
.Y(n_4028)
);

AOI21xp5_ASAP7_75t_L g4029 ( 
.A1(n_3994),
.A2(n_3349),
.B(n_3498),
.Y(n_4029)
);

AND2x2_ASAP7_75t_L g4030 ( 
.A(n_3876),
.B(n_3930),
.Y(n_4030)
);

BUFx6f_ASAP7_75t_L g4031 ( 
.A(n_3722),
.Y(n_4031)
);

AOI21xp5_ASAP7_75t_L g4032 ( 
.A1(n_3717),
.A2(n_3500),
.B(n_3498),
.Y(n_4032)
);

AND2x2_ASAP7_75t_L g4033 ( 
.A(n_3918),
.B(n_3584),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3763),
.B(n_3646),
.Y(n_4034)
);

CKINVDCx20_ASAP7_75t_R g4035 ( 
.A(n_3755),
.Y(n_4035)
);

OAI21xp33_ASAP7_75t_L g4036 ( 
.A1(n_3821),
.A2(n_3679),
.B(n_3597),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3765),
.B(n_3679),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_3831),
.Y(n_4038)
);

A2O1A1Ixp33_ASAP7_75t_L g4039 ( 
.A1(n_3740),
.A2(n_3487),
.B(n_3712),
.C(n_3646),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3947),
.B(n_3480),
.Y(n_4040)
);

BUFx6f_ASAP7_75t_L g4041 ( 
.A(n_3722),
.Y(n_4041)
);

A2O1A1Ixp33_ASAP7_75t_L g4042 ( 
.A1(n_3779),
.A2(n_3639),
.B(n_3674),
.C(n_3650),
.Y(n_4042)
);

OAI21xp33_ASAP7_75t_L g4043 ( 
.A1(n_3938),
.A2(n_1036),
.B(n_1035),
.Y(n_4043)
);

O2A1O1Ixp33_ASAP7_75t_SL g4044 ( 
.A1(n_3872),
.A2(n_3548),
.B(n_3516),
.C(n_3536),
.Y(n_4044)
);

AOI21xp5_ASAP7_75t_L g4045 ( 
.A1(n_3852),
.A2(n_3506),
.B(n_3500),
.Y(n_4045)
);

NAND2xp5_ASAP7_75t_SL g4046 ( 
.A(n_3929),
.B(n_3577),
.Y(n_4046)
);

NOR2xp33_ASAP7_75t_L g4047 ( 
.A(n_4002),
.B(n_3670),
.Y(n_4047)
);

AOI21xp5_ASAP7_75t_L g4048 ( 
.A1(n_3969),
.A2(n_3506),
.B(n_3530),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3750),
.Y(n_4049)
);

AOI21xp5_ASAP7_75t_L g4050 ( 
.A1(n_3724),
.A2(n_3541),
.B(n_3535),
.Y(n_4050)
);

AOI21xp5_ASAP7_75t_L g4051 ( 
.A1(n_3878),
.A2(n_3546),
.B(n_3544),
.Y(n_4051)
);

AOI21x1_ASAP7_75t_L g4052 ( 
.A1(n_3881),
.A2(n_3673),
.B(n_3665),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3771),
.B(n_3318),
.Y(n_4053)
);

OAI21xp5_ASAP7_75t_L g4054 ( 
.A1(n_3726),
.A2(n_3684),
.B(n_3678),
.Y(n_4054)
);

AOI21xp5_ASAP7_75t_L g4055 ( 
.A1(n_3886),
.A2(n_3588),
.B(n_3587),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3751),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3816),
.B(n_3677),
.Y(n_4057)
);

INVx4_ASAP7_75t_L g4058 ( 
.A(n_3722),
.Y(n_4058)
);

NOR2x1_ASAP7_75t_L g4059 ( 
.A(n_3838),
.B(n_3889),
.Y(n_4059)
);

AOI21xp5_ASAP7_75t_L g4060 ( 
.A1(n_3845),
.A2(n_3588),
.B(n_3587),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3877),
.Y(n_4061)
);

INVx3_ASAP7_75t_L g4062 ( 
.A(n_3790),
.Y(n_4062)
);

AND2x4_ASAP7_75t_L g4063 ( 
.A(n_3790),
.B(n_3524),
.Y(n_4063)
);

NOR2xp33_ASAP7_75t_L g4064 ( 
.A(n_3896),
.B(n_3343),
.Y(n_4064)
);

AOI21xp5_ASAP7_75t_L g4065 ( 
.A1(n_3807),
.A2(n_3675),
.B(n_3673),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3825),
.B(n_3593),
.Y(n_4066)
);

O2A1O1Ixp5_ASAP7_75t_L g4067 ( 
.A1(n_3731),
.A2(n_3475),
.B(n_3499),
.C(n_3479),
.Y(n_4067)
);

NOR2xp33_ASAP7_75t_L g4068 ( 
.A(n_3915),
.B(n_3373),
.Y(n_4068)
);

AOI21xp5_ASAP7_75t_L g4069 ( 
.A1(n_3803),
.A2(n_3675),
.B(n_3592),
.Y(n_4069)
);

AND2x4_ASAP7_75t_L g4070 ( 
.A(n_3838),
.B(n_3605),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_SL g4071 ( 
.A(n_3832),
.B(n_3596),
.Y(n_4071)
);

AOI21xp5_ASAP7_75t_L g4072 ( 
.A1(n_3785),
.A2(n_3501),
.B(n_3553),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3759),
.Y(n_4073)
);

AOI21xp5_ASAP7_75t_L g4074 ( 
.A1(n_3835),
.A2(n_3555),
.B(n_3554),
.Y(n_4074)
);

O2A1O1Ixp5_ASAP7_75t_L g4075 ( 
.A1(n_3949),
.A2(n_3408),
.B(n_3672),
.C(n_3662),
.Y(n_4075)
);

NOR2x1p5_ASAP7_75t_L g4076 ( 
.A(n_3927),
.B(n_3346),
.Y(n_4076)
);

AND2x2_ASAP7_75t_L g4077 ( 
.A(n_3766),
.B(n_3406),
.Y(n_4077)
);

AOI21xp5_ASAP7_75t_L g4078 ( 
.A1(n_3776),
.A2(n_3571),
.B(n_3565),
.Y(n_4078)
);

AOI21xp5_ASAP7_75t_L g4079 ( 
.A1(n_3874),
.A2(n_3602),
.B(n_3574),
.Y(n_4079)
);

AND2x2_ASAP7_75t_L g4080 ( 
.A(n_3837),
.B(n_3427),
.Y(n_4080)
);

AOI22xp5_ASAP7_75t_L g4081 ( 
.A1(n_3952),
.A2(n_3517),
.B1(n_3394),
.B2(n_3556),
.Y(n_4081)
);

NOR2x1_ASAP7_75t_L g4082 ( 
.A(n_3764),
.B(n_3667),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_3777),
.B(n_3693),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_SL g4084 ( 
.A(n_3792),
.B(n_3609),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_3890),
.Y(n_4085)
);

AOI21xp5_ASAP7_75t_L g4086 ( 
.A1(n_3721),
.A2(n_3603),
.B(n_3616),
.Y(n_4086)
);

OAI21xp5_ASAP7_75t_L g4087 ( 
.A1(n_3773),
.A2(n_3875),
.B(n_3742),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3955),
.Y(n_4088)
);

NOR2xp33_ASAP7_75t_L g4089 ( 
.A(n_3922),
.B(n_3441),
.Y(n_4089)
);

AND2x2_ASAP7_75t_L g4090 ( 
.A(n_3963),
.B(n_3449),
.Y(n_4090)
);

OAI22xp5_ASAP7_75t_L g4091 ( 
.A1(n_3769),
.A2(n_3687),
.B1(n_3697),
.B2(n_3681),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_SL g4092 ( 
.A(n_3984),
.B(n_3612),
.Y(n_4092)
);

AOI21xp5_ASAP7_75t_L g4093 ( 
.A1(n_3756),
.A2(n_3619),
.B(n_3618),
.Y(n_4093)
);

AOI221xp5_ASAP7_75t_SL g4094 ( 
.A1(n_3974),
.A2(n_3856),
.B1(n_3959),
.B2(n_3823),
.C(n_3820),
.Y(n_4094)
);

INVx3_ASAP7_75t_SL g4095 ( 
.A(n_3987),
.Y(n_4095)
);

AOI21xp5_ASAP7_75t_L g4096 ( 
.A1(n_3760),
.A2(n_3622),
.B(n_3621),
.Y(n_4096)
);

AOI21xp5_ASAP7_75t_L g4097 ( 
.A1(n_3972),
.A2(n_3645),
.B(n_3630),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_SL g4098 ( 
.A(n_3805),
.B(n_3620),
.Y(n_4098)
);

INVx2_ASAP7_75t_L g4099 ( 
.A(n_3990),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3767),
.B(n_3660),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_SL g4101 ( 
.A(n_3784),
.B(n_3661),
.Y(n_4101)
);

BUFx6f_ASAP7_75t_L g4102 ( 
.A(n_3737),
.Y(n_4102)
);

AND2x4_ASAP7_75t_SL g4103 ( 
.A(n_3737),
.B(n_3667),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3791),
.B(n_3700),
.Y(n_4104)
);

OAI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_3884),
.A2(n_3707),
.B1(n_3710),
.B2(n_3705),
.Y(n_4105)
);

AND2x6_ASAP7_75t_L g4106 ( 
.A(n_3901),
.B(n_3713),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_4004),
.Y(n_4107)
);

AOI21xp5_ASAP7_75t_L g4108 ( 
.A1(n_3822),
.A2(n_3663),
.B(n_3658),
.Y(n_4108)
);

INVx2_ASAP7_75t_L g4109 ( 
.A(n_4007),
.Y(n_4109)
);

OAI22xp5_ASAP7_75t_L g4110 ( 
.A1(n_3924),
.A2(n_3655),
.B1(n_3659),
.B2(n_3611),
.Y(n_4110)
);

AOI21xp5_ASAP7_75t_L g4111 ( 
.A1(n_3723),
.A2(n_3476),
.B(n_3691),
.Y(n_4111)
);

AND2x4_ASAP7_75t_L g4112 ( 
.A(n_3737),
.B(n_3346),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_3793),
.B(n_3727),
.Y(n_4113)
);

AOI22xp33_ASAP7_75t_L g4114 ( 
.A1(n_3997),
.A2(n_3517),
.B1(n_3556),
.B2(n_3455),
.Y(n_4114)
);

AOI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_3951),
.A2(n_3556),
.B1(n_3471),
.B2(n_3484),
.Y(n_4115)
);

BUFx6f_ASAP7_75t_L g4116 ( 
.A(n_3753),
.Y(n_4116)
);

INVx3_ASAP7_75t_L g4117 ( 
.A(n_3733),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_SL g4118 ( 
.A(n_3799),
.B(n_3691),
.Y(n_4118)
);

OAI22xp5_ASAP7_75t_L g4119 ( 
.A1(n_3924),
.A2(n_3496),
.B1(n_3497),
.B2(n_3494),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_3870),
.B(n_3456),
.Y(n_4120)
);

BUFx12f_ASAP7_75t_L g4121 ( 
.A(n_3725),
.Y(n_4121)
);

BUFx12f_ASAP7_75t_L g4122 ( 
.A(n_3725),
.Y(n_4122)
);

AOI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_3840),
.A2(n_3671),
.B(n_3664),
.Y(n_4123)
);

BUFx6f_ASAP7_75t_L g4124 ( 
.A(n_3753),
.Y(n_4124)
);

AOI22xp5_ASAP7_75t_L g4125 ( 
.A1(n_3900),
.A2(n_3556),
.B1(n_3508),
.B2(n_3493),
.Y(n_4125)
);

AOI21xp5_ASAP7_75t_L g4126 ( 
.A1(n_3781),
.A2(n_3680),
.B(n_3345),
.Y(n_4126)
);

NOR3xp33_ASAP7_75t_L g4127 ( 
.A(n_3891),
.B(n_1521),
.C(n_1518),
.Y(n_4127)
);

NOR2xp33_ASAP7_75t_L g4128 ( 
.A(n_3802),
.B(n_3413),
.Y(n_4128)
);

NOR2xp33_ASAP7_75t_L g4129 ( 
.A(n_3961),
.B(n_3839),
.Y(n_4129)
);

OAI22xp5_ASAP7_75t_L g4130 ( 
.A1(n_4001),
.A2(n_3447),
.B1(n_3413),
.B2(n_3590),
.Y(n_4130)
);

NOR2xp33_ASAP7_75t_SL g4131 ( 
.A(n_3729),
.B(n_3629),
.Y(n_4131)
);

A2O1A1Ixp33_ASAP7_75t_L g4132 ( 
.A1(n_3741),
.A2(n_3447),
.B(n_1175),
.C(n_1176),
.Y(n_4132)
);

INVx2_ASAP7_75t_SL g4133 ( 
.A(n_3815),
.Y(n_4133)
);

INVx3_ASAP7_75t_SL g4134 ( 
.A(n_3880),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_3797),
.B(n_1524),
.Y(n_4135)
);

A2O1A1Ixp33_ASAP7_75t_L g4136 ( 
.A1(n_3954),
.A2(n_1175),
.B(n_1176),
.C(n_1172),
.Y(n_4136)
);

INVx2_ASAP7_75t_L g4137 ( 
.A(n_4008),
.Y(n_4137)
);

AND2x4_ASAP7_75t_L g4138 ( 
.A(n_3753),
.B(n_3629),
.Y(n_4138)
);

AOI22xp5_ASAP7_75t_L g4139 ( 
.A1(n_3826),
.A2(n_1040),
.B1(n_1042),
.B2(n_1039),
.Y(n_4139)
);

BUFx6f_ASAP7_75t_L g4140 ( 
.A(n_3758),
.Y(n_4140)
);

HB1xp67_ASAP7_75t_L g4141 ( 
.A(n_3812),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_SL g4142 ( 
.A(n_3849),
.B(n_3629),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3761),
.Y(n_4143)
);

BUFx12f_ASAP7_75t_L g4144 ( 
.A(n_3880),
.Y(n_4144)
);

AOI33xp33_ASAP7_75t_L g4145 ( 
.A1(n_3860),
.A2(n_1200),
.A3(n_1186),
.B1(n_1201),
.B2(n_1189),
.B3(n_1181),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_3861),
.B(n_3345),
.Y(n_4146)
);

NOR2xp33_ASAP7_75t_L g4147 ( 
.A(n_3944),
.B(n_1047),
.Y(n_4147)
);

AND2x2_ASAP7_75t_L g4148 ( 
.A(n_3797),
.B(n_1526),
.Y(n_4148)
);

AOI21xp5_ASAP7_75t_L g4149 ( 
.A1(n_3732),
.A2(n_3345),
.B(n_2361),
.Y(n_4149)
);

OAI21xp5_ASAP7_75t_L g4150 ( 
.A1(n_3968),
.A2(n_3345),
.B(n_2364),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_SL g4151 ( 
.A(n_3849),
.B(n_1049),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_SL g4152 ( 
.A(n_3851),
.B(n_1050),
.Y(n_4152)
);

OAI22xp5_ASAP7_75t_L g4153 ( 
.A1(n_3859),
.A2(n_1052),
.B1(n_1053),
.B2(n_1051),
.Y(n_4153)
);

NOR2xp67_ASAP7_75t_SL g4154 ( 
.A(n_3903),
.B(n_1181),
.Y(n_4154)
);

AOI21xp5_ASAP7_75t_L g4155 ( 
.A1(n_3735),
.A2(n_3345),
.B(n_2370),
.Y(n_4155)
);

OAI21x1_ASAP7_75t_L g4156 ( 
.A1(n_3757),
.A2(n_2265),
.B(n_2263),
.Y(n_4156)
);

NOR2xp33_ASAP7_75t_L g4157 ( 
.A(n_3836),
.B(n_1059),
.Y(n_4157)
);

NOR2xp33_ASAP7_75t_SL g4158 ( 
.A(n_3754),
.B(n_3433),
.Y(n_4158)
);

NOR2xp67_ASAP7_75t_L g4159 ( 
.A(n_3801),
.B(n_2266),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_3848),
.B(n_1527),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3772),
.Y(n_4161)
);

AOI21xp5_ASAP7_75t_L g4162 ( 
.A1(n_3738),
.A2(n_3748),
.B(n_3747),
.Y(n_4162)
);

OAI22xp5_ASAP7_75t_L g4163 ( 
.A1(n_3893),
.A2(n_1061),
.B1(n_1067),
.B2(n_1060),
.Y(n_4163)
);

NOR2xp33_ASAP7_75t_L g4164 ( 
.A(n_3847),
.B(n_3800),
.Y(n_4164)
);

INVx4_ASAP7_75t_L g4165 ( 
.A(n_3758),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_3866),
.B(n_1068),
.Y(n_4166)
);

AOI22x1_ASAP7_75t_L g4167 ( 
.A1(n_3844),
.A2(n_1189),
.B1(n_1200),
.B2(n_1186),
.Y(n_4167)
);

OA22x2_ASAP7_75t_L g4168 ( 
.A1(n_3928),
.A2(n_1071),
.B1(n_1074),
.B2(n_1070),
.Y(n_4168)
);

O2A1O1Ixp33_ASAP7_75t_SL g4169 ( 
.A1(n_3746),
.A2(n_3752),
.B(n_3736),
.C(n_3965),
.Y(n_4169)
);

INVx2_ASAP7_75t_L g4170 ( 
.A(n_3778),
.Y(n_4170)
);

NOR2xp33_ASAP7_75t_R g4171 ( 
.A(n_3758),
.B(n_635),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_SL g4172 ( 
.A(n_3851),
.B(n_1075),
.Y(n_4172)
);

NOR2xp33_ASAP7_75t_L g4173 ( 
.A(n_3814),
.B(n_1076),
.Y(n_4173)
);

AOI21xp5_ASAP7_75t_L g4174 ( 
.A1(n_3768),
.A2(n_2371),
.B(n_2358),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_SL g4175 ( 
.A(n_3975),
.B(n_1077),
.Y(n_4175)
);

O2A1O1Ixp33_ASAP7_75t_SL g4176 ( 
.A1(n_3774),
.A2(n_1203),
.B(n_1205),
.C(n_1201),
.Y(n_4176)
);

NOR2xp67_ASAP7_75t_L g4177 ( 
.A(n_3787),
.B(n_2270),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_SL g4178 ( 
.A(n_3975),
.B(n_4006),
.Y(n_4178)
);

BUFx8_ASAP7_75t_L g4179 ( 
.A(n_3786),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_3789),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_3806),
.B(n_3775),
.Y(n_4181)
);

O2A1O1Ixp33_ASAP7_75t_L g4182 ( 
.A1(n_3780),
.A2(n_1205),
.B(n_1211),
.C(n_1203),
.Y(n_4182)
);

AOI21xp5_ASAP7_75t_L g4183 ( 
.A1(n_3770),
.A2(n_2376),
.B(n_2374),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_3811),
.B(n_1079),
.Y(n_4184)
);

AOI21xp5_ASAP7_75t_L g4185 ( 
.A1(n_3788),
.A2(n_2388),
.B(n_2378),
.Y(n_4185)
);

AOI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_3911),
.A2(n_2415),
.B(n_2411),
.Y(n_4186)
);

BUFx2_ASAP7_75t_L g4187 ( 
.A(n_3971),
.Y(n_4187)
);

AND2x2_ASAP7_75t_L g4188 ( 
.A(n_3898),
.B(n_1529),
.Y(n_4188)
);

AOI22x1_ASAP7_75t_L g4189 ( 
.A1(n_3813),
.A2(n_1213),
.B1(n_1215),
.B2(n_1211),
.Y(n_4189)
);

AOI22xp5_ASAP7_75t_L g4190 ( 
.A1(n_3954),
.A2(n_1083),
.B1(n_1084),
.B2(n_1080),
.Y(n_4190)
);

CKINVDCx10_ASAP7_75t_R g4191 ( 
.A(n_3786),
.Y(n_4191)
);

AOI21xp5_ASAP7_75t_L g4192 ( 
.A1(n_3795),
.A2(n_2421),
.B(n_2420),
.Y(n_4192)
);

AOI21xp5_ASAP7_75t_L g4193 ( 
.A1(n_3798),
.A2(n_2427),
.B(n_2423),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_3794),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_SL g4195 ( 
.A(n_3928),
.B(n_1085),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_3862),
.Y(n_4196)
);

AOI21xp5_ASAP7_75t_L g4197 ( 
.A1(n_3996),
.A2(n_2432),
.B(n_2431),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_SL g4198 ( 
.A(n_3898),
.B(n_1087),
.Y(n_4198)
);

OAI21xp5_ASAP7_75t_L g4199 ( 
.A1(n_3887),
.A2(n_2441),
.B(n_2437),
.Y(n_4199)
);

AOI21xp5_ASAP7_75t_L g4200 ( 
.A1(n_3998),
.A2(n_2445),
.B(n_2444),
.Y(n_4200)
);

AOI22xp33_ASAP7_75t_L g4201 ( 
.A1(n_3818),
.A2(n_1215),
.B1(n_1217),
.B2(n_1213),
.Y(n_4201)
);

INVx2_ASAP7_75t_L g4202 ( 
.A(n_3863),
.Y(n_4202)
);

OR2x6_ASAP7_75t_L g4203 ( 
.A(n_3786),
.B(n_1217),
.Y(n_4203)
);

NAND2xp33_ASAP7_75t_L g4204 ( 
.A(n_3867),
.B(n_3818),
.Y(n_4204)
);

AOI21xp5_ASAP7_75t_L g4205 ( 
.A1(n_4005),
.A2(n_2451),
.B(n_2448),
.Y(n_4205)
);

INVxp67_ASAP7_75t_L g4206 ( 
.A(n_3999),
.Y(n_4206)
);

OAI22xp5_ASAP7_75t_L g4207 ( 
.A1(n_3882),
.A2(n_1090),
.B1(n_1092),
.B2(n_1089),
.Y(n_4207)
);

INVx3_ASAP7_75t_L g4208 ( 
.A(n_3733),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_3841),
.B(n_1094),
.Y(n_4209)
);

AOI22xp5_ASAP7_75t_L g4210 ( 
.A1(n_3913),
.A2(n_1100),
.B1(n_1103),
.B2(n_1095),
.Y(n_4210)
);

AOI21xp5_ASAP7_75t_L g4211 ( 
.A1(n_3846),
.A2(n_2137),
.B(n_2102),
.Y(n_4211)
);

HB1xp67_ASAP7_75t_L g4212 ( 
.A(n_3888),
.Y(n_4212)
);

OAI21xp33_ASAP7_75t_L g4213 ( 
.A1(n_3906),
.A2(n_1107),
.B(n_1104),
.Y(n_4213)
);

NOR2xp33_ASAP7_75t_L g4214 ( 
.A(n_3919),
.B(n_1111),
.Y(n_4214)
);

AOI21xp5_ASAP7_75t_L g4215 ( 
.A1(n_3868),
.A2(n_2146),
.B(n_2137),
.Y(n_4215)
);

O2A1O1Ixp33_ASAP7_75t_L g4216 ( 
.A1(n_3976),
.A2(n_1219),
.B(n_1220),
.C(n_1218),
.Y(n_4216)
);

INVx2_ASAP7_75t_L g4217 ( 
.A(n_3895),
.Y(n_4217)
);

AOI21xp5_ASAP7_75t_L g4218 ( 
.A1(n_3869),
.A2(n_3905),
.B(n_3883),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_L g4219 ( 
.A(n_3897),
.B(n_1114),
.Y(n_4219)
);

OAI21xp5_ASAP7_75t_L g4220 ( 
.A1(n_3743),
.A2(n_2273),
.B(n_2272),
.Y(n_4220)
);

AOI22x1_ASAP7_75t_L g4221 ( 
.A1(n_3909),
.A2(n_1219),
.B1(n_1220),
.B2(n_1218),
.Y(n_4221)
);

OAI22xp5_ASAP7_75t_L g4222 ( 
.A1(n_3916),
.A2(n_1116),
.B1(n_1118),
.B2(n_1115),
.Y(n_4222)
);

OAI22xp5_ASAP7_75t_L g4223 ( 
.A1(n_3920),
.A2(n_3942),
.B1(n_3979),
.B2(n_3937),
.Y(n_4223)
);

O2A1O1Ixp5_ASAP7_75t_L g4224 ( 
.A1(n_3946),
.A2(n_1225),
.B(n_1231),
.C(n_1221),
.Y(n_4224)
);

AND2x2_ASAP7_75t_SL g4225 ( 
.A(n_3853),
.B(n_1221),
.Y(n_4225)
);

O2A1O1Ixp33_ASAP7_75t_L g4226 ( 
.A1(n_3925),
.A2(n_1231),
.B(n_1234),
.C(n_1225),
.Y(n_4226)
);

OAI21xp5_ASAP7_75t_L g4227 ( 
.A1(n_3894),
.A2(n_2278),
.B(n_2275),
.Y(n_4227)
);

BUFx4f_ASAP7_75t_L g4228 ( 
.A(n_3850),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3980),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_3982),
.Y(n_4230)
);

INVxp67_ASAP7_75t_L g4231 ( 
.A(n_3850),
.Y(n_4231)
);

AOI21xp5_ASAP7_75t_L g4232 ( 
.A1(n_3879),
.A2(n_2177),
.B(n_2146),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_3931),
.Y(n_4233)
);

INVx3_ASAP7_75t_L g4234 ( 
.A(n_3853),
.Y(n_4234)
);

OAI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_3933),
.A2(n_1122),
.B1(n_1125),
.B2(n_1120),
.Y(n_4235)
);

OAI22xp5_ASAP7_75t_L g4236 ( 
.A1(n_3843),
.A2(n_1136),
.B1(n_1137),
.B2(n_1127),
.Y(n_4236)
);

OAI21xp33_ASAP7_75t_SL g4237 ( 
.A1(n_3843),
.A2(n_1235),
.B(n_1234),
.Y(n_4237)
);

NOR2xp33_ASAP7_75t_L g4238 ( 
.A(n_3950),
.B(n_1142),
.Y(n_4238)
);

AOI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_3962),
.A2(n_2177),
.B(n_2146),
.Y(n_4239)
);

INVx1_ASAP7_75t_SL g4240 ( 
.A(n_3850),
.Y(n_4240)
);

OAI22xp5_ASAP7_75t_L g4241 ( 
.A1(n_3892),
.A2(n_1147),
.B1(n_1152),
.B2(n_1145),
.Y(n_4241)
);

INVx2_ASAP7_75t_L g4242 ( 
.A(n_3808),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_3810),
.B(n_1154),
.Y(n_4243)
);

BUFx6f_ASAP7_75t_L g4244 ( 
.A(n_3885),
.Y(n_4244)
);

OAI22xp5_ASAP7_75t_L g4245 ( 
.A1(n_3892),
.A2(n_1156),
.B1(n_1160),
.B2(n_1155),
.Y(n_4245)
);

BUFx8_ASAP7_75t_L g4246 ( 
.A(n_3885),
.Y(n_4246)
);

NOR2x1_ASAP7_75t_L g4247 ( 
.A(n_3901),
.B(n_2355),
.Y(n_4247)
);

AOI21xp5_ASAP7_75t_L g4248 ( 
.A1(n_3966),
.A2(n_2177),
.B(n_2146),
.Y(n_4248)
);

BUFx4f_ASAP7_75t_L g4249 ( 
.A(n_3885),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_3948),
.B(n_1161),
.Y(n_4250)
);

O2A1O1Ixp33_ASAP7_75t_L g4251 ( 
.A1(n_3762),
.A2(n_1235),
.B(n_1531),
.C(n_1530),
.Y(n_4251)
);

AND2x4_ASAP7_75t_L g4252 ( 
.A(n_3833),
.B(n_3914),
.Y(n_4252)
);

AND2x4_ASAP7_75t_L g4253 ( 
.A(n_3833),
.B(n_3914),
.Y(n_4253)
);

O2A1O1Ixp33_ASAP7_75t_L g4254 ( 
.A1(n_3827),
.A2(n_1533),
.B(n_1535),
.C(n_1532),
.Y(n_4254)
);

OAI22xp5_ASAP7_75t_L g4255 ( 
.A1(n_3824),
.A2(n_1167),
.B1(n_1169),
.B2(n_1164),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_3953),
.B(n_1170),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_3958),
.B(n_1171),
.Y(n_4257)
);

NOR2xp33_ASAP7_75t_L g4258 ( 
.A(n_3964),
.B(n_1173),
.Y(n_4258)
);

CKINVDCx11_ASAP7_75t_R g4259 ( 
.A(n_3932),
.Y(n_4259)
);

AOI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_3973),
.A2(n_2178),
.B(n_2177),
.Y(n_4260)
);

O2A1O1Ixp33_ASAP7_75t_L g4261 ( 
.A1(n_3977),
.A2(n_1539),
.B(n_1540),
.C(n_1536),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_3986),
.B(n_1174),
.Y(n_4262)
);

INVxp67_ASAP7_75t_R g4263 ( 
.A(n_3983),
.Y(n_4263)
);

NOR2xp67_ASAP7_75t_L g4264 ( 
.A(n_3939),
.B(n_2280),
.Y(n_4264)
);

CKINVDCx20_ASAP7_75t_R g4265 ( 
.A(n_3932),
.Y(n_4265)
);

AOI21xp5_ASAP7_75t_L g4266 ( 
.A1(n_3985),
.A2(n_2193),
.B(n_2178),
.Y(n_4266)
);

A2O1A1Ixp33_ASAP7_75t_L g4267 ( 
.A1(n_3906),
.A2(n_1179),
.B(n_1182),
.C(n_1177),
.Y(n_4267)
);

BUFx8_ASAP7_75t_L g4268 ( 
.A(n_3932),
.Y(n_4268)
);

BUFx3_ASAP7_75t_L g4269 ( 
.A(n_3970),
.Y(n_4269)
);

AOI21xp5_ASAP7_75t_L g4270 ( 
.A1(n_3988),
.A2(n_2193),
.B(n_2178),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_3989),
.B(n_1183),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_3991),
.B(n_1542),
.Y(n_4272)
);

BUFx8_ASAP7_75t_SL g4273 ( 
.A(n_3970),
.Y(n_4273)
);

NOR2x1_ASAP7_75t_SL g4274 ( 
.A(n_4016),
.B(n_3995),
.Y(n_4274)
);

INVx3_ASAP7_75t_L g4275 ( 
.A(n_4252),
.Y(n_4275)
);

OAI21x1_ASAP7_75t_L g4276 ( 
.A1(n_4156),
.A2(n_3828),
.B(n_3992),
.Y(n_4276)
);

AO32x2_ASAP7_75t_L g4277 ( 
.A1(n_4223),
.A2(n_4003),
.A3(n_3981),
.B1(n_3960),
.B2(n_3907),
.Y(n_4277)
);

OAI21x1_ASAP7_75t_L g4278 ( 
.A1(n_4162),
.A2(n_3921),
.B(n_3917),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4212),
.Y(n_4279)
);

NOR2xp33_ASAP7_75t_L g4280 ( 
.A(n_4012),
.B(n_3970),
.Y(n_4280)
);

BUFx2_ASAP7_75t_L g4281 ( 
.A(n_4265),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_4113),
.B(n_4181),
.Y(n_4282)
);

AOI221x1_ASAP7_75t_L g4283 ( 
.A1(n_4025),
.A2(n_3902),
.B1(n_3967),
.B2(n_3904),
.C(n_3873),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_4242),
.B(n_4000),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4049),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_4233),
.B(n_4018),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4030),
.B(n_3978),
.Y(n_4287)
);

AOI21xp5_ASAP7_75t_L g4288 ( 
.A1(n_4029),
.A2(n_3782),
.B(n_3871),
.Y(n_4288)
);

NOR2xp33_ASAP7_75t_L g4289 ( 
.A(n_4011),
.B(n_3978),
.Y(n_4289)
);

BUFx6f_ASAP7_75t_L g4290 ( 
.A(n_4259),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_4022),
.B(n_3978),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4056),
.Y(n_4292)
);

AO31x2_ASAP7_75t_L g4293 ( 
.A1(n_4218),
.A2(n_3956),
.A3(n_3943),
.B(n_3945),
.Y(n_4293)
);

BUFx2_ASAP7_75t_L g4294 ( 
.A(n_4010),
.Y(n_4294)
);

OAI21xp5_ASAP7_75t_L g4295 ( 
.A1(n_4094),
.A2(n_4224),
.B(n_4015),
.Y(n_4295)
);

INVx4_ASAP7_75t_L g4296 ( 
.A(n_4228),
.Y(n_4296)
);

INVx3_ASAP7_75t_L g4297 ( 
.A(n_4252),
.Y(n_4297)
);

OAI22xp5_ASAP7_75t_L g4298 ( 
.A1(n_4017),
.A2(n_3749),
.B1(n_3957),
.B2(n_3940),
.Y(n_4298)
);

NOR2xp33_ASAP7_75t_L g4299 ( 
.A(n_4021),
.B(n_3939),
.Y(n_4299)
);

NAND2xp33_ASAP7_75t_L g4300 ( 
.A(n_4059),
.B(n_3940),
.Y(n_4300)
);

AO31x2_ASAP7_75t_L g4301 ( 
.A1(n_4149),
.A2(n_4155),
.A3(n_4060),
.B(n_4024),
.Y(n_4301)
);

OAI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_4097),
.A2(n_3910),
.B(n_4009),
.Y(n_4302)
);

AOI21xp5_ASAP7_75t_L g4303 ( 
.A1(n_4048),
.A2(n_3855),
.B(n_3854),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_4083),
.B(n_1184),
.Y(n_4304)
);

AO31x2_ASAP7_75t_L g4305 ( 
.A1(n_4019),
.A2(n_4215),
.A3(n_4211),
.B(n_4051),
.Y(n_4305)
);

A2O1A1Ixp33_ASAP7_75t_L g4306 ( 
.A1(n_4145),
.A2(n_3957),
.B(n_3993),
.C(n_3783),
.Y(n_4306)
);

NAND2x1p5_ASAP7_75t_L g4307 ( 
.A(n_4228),
.B(n_3993),
.Y(n_4307)
);

A2O1A1Ixp33_ASAP7_75t_L g4308 ( 
.A1(n_4036),
.A2(n_3829),
.B(n_3864),
.C(n_3858),
.Y(n_4308)
);

OA21x2_ASAP7_75t_L g4309 ( 
.A1(n_4087),
.A2(n_3912),
.B(n_3926),
.Y(n_4309)
);

BUFx6f_ASAP7_75t_L g4310 ( 
.A(n_4249),
.Y(n_4310)
);

OAI22xp5_ASAP7_75t_L g4311 ( 
.A1(n_4064),
.A2(n_4046),
.B1(n_4114),
.B2(n_4081),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_4100),
.B(n_4068),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_4037),
.B(n_4104),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_4073),
.Y(n_4314)
);

OAI21x1_ASAP7_75t_L g4315 ( 
.A1(n_4197),
.A2(n_3935),
.B(n_3934),
.Y(n_4315)
);

OR2x2_ASAP7_75t_L g4316 ( 
.A(n_4026),
.B(n_1545),
.Y(n_4316)
);

OAI21x1_ASAP7_75t_L g4317 ( 
.A1(n_4200),
.A2(n_3941),
.B(n_2286),
.Y(n_4317)
);

AOI211x1_ASAP7_75t_L g4318 ( 
.A1(n_4014),
.A2(n_1551),
.B(n_1552),
.C(n_1547),
.Y(n_4318)
);

AOI221x1_ASAP7_75t_L g4319 ( 
.A1(n_4111),
.A2(n_1556),
.B1(n_1557),
.B2(n_1554),
.C(n_1553),
.Y(n_4319)
);

OAI22xp5_ASAP7_75t_L g4320 ( 
.A1(n_4023),
.A2(n_1187),
.B1(n_1191),
.B2(n_1185),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4143),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_4053),
.B(n_4040),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_4034),
.B(n_1558),
.Y(n_4323)
);

OAI21x1_ASAP7_75t_L g4324 ( 
.A1(n_4205),
.A2(n_2287),
.B(n_2283),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_4057),
.B(n_1194),
.Y(n_4325)
);

INVx2_ASAP7_75t_L g4326 ( 
.A(n_4170),
.Y(n_4326)
);

OAI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_4267),
.A2(n_1561),
.B(n_1560),
.Y(n_4327)
);

OAI21xp33_ASAP7_75t_L g4328 ( 
.A1(n_4213),
.A2(n_1198),
.B(n_1196),
.Y(n_4328)
);

OAI21x1_ASAP7_75t_L g4329 ( 
.A1(n_4174),
.A2(n_2292),
.B(n_2291),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4161),
.Y(n_4330)
);

OAI21xp5_ASAP7_75t_L g4331 ( 
.A1(n_4238),
.A2(n_1564),
.B(n_1562),
.Y(n_4331)
);

AOI21xp5_ASAP7_75t_L g4332 ( 
.A1(n_4045),
.A2(n_2309),
.B(n_2293),
.Y(n_4332)
);

AOI21xp5_ASAP7_75t_L g4333 ( 
.A1(n_4065),
.A2(n_4074),
.B(n_4032),
.Y(n_4333)
);

OAI21x1_ASAP7_75t_L g4334 ( 
.A1(n_4183),
.A2(n_2315),
.B(n_2311),
.Y(n_4334)
);

AOI21xp5_ASAP7_75t_L g4335 ( 
.A1(n_4078),
.A2(n_2318),
.B(n_2203),
.Y(n_4335)
);

INVx1_ASAP7_75t_SL g4336 ( 
.A(n_4187),
.Y(n_4336)
);

OAI21x1_ASAP7_75t_L g4337 ( 
.A1(n_4185),
.A2(n_2205),
.B(n_2190),
.Y(n_4337)
);

NAND2x1p5_ASAP7_75t_L g4338 ( 
.A(n_4249),
.B(n_2178),
.Y(n_4338)
);

INVx2_ASAP7_75t_L g4339 ( 
.A(n_4194),
.Y(n_4339)
);

INVx3_ASAP7_75t_L g4340 ( 
.A(n_4273),
.Y(n_4340)
);

AOI221x1_ASAP7_75t_L g4341 ( 
.A1(n_4136),
.A2(n_1568),
.B1(n_1569),
.B2(n_1567),
.C(n_1565),
.Y(n_4341)
);

OAI21x1_ASAP7_75t_L g4342 ( 
.A1(n_4050),
.A2(n_2224),
.B(n_2205),
.Y(n_4342)
);

OAI21xp5_ASAP7_75t_L g4343 ( 
.A1(n_4175),
.A2(n_1571),
.B(n_1570),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_L g4344 ( 
.A(n_4066),
.B(n_1199),
.Y(n_4344)
);

INVx5_ASAP7_75t_L g4345 ( 
.A(n_4106),
.Y(n_4345)
);

AOI22x1_ASAP7_75t_L g4346 ( 
.A1(n_4263),
.A2(n_1204),
.B1(n_1207),
.B2(n_1202),
.Y(n_4346)
);

NAND2xp5_ASAP7_75t_L g4347 ( 
.A(n_4120),
.B(n_1208),
.Y(n_4347)
);

HB1xp67_ASAP7_75t_L g4348 ( 
.A(n_4141),
.Y(n_4348)
);

NAND3xp33_ASAP7_75t_SL g4349 ( 
.A(n_4190),
.B(n_1212),
.C(n_1210),
.Y(n_4349)
);

OAI21x1_ASAP7_75t_L g4350 ( 
.A1(n_4186),
.A2(n_2282),
.B(n_2224),
.Y(n_4350)
);

OAI22x1_ASAP7_75t_L g4351 ( 
.A1(n_4167),
.A2(n_4033),
.B1(n_4071),
.B2(n_4092),
.Y(n_4351)
);

NAND3x1_ASAP7_75t_L g4352 ( 
.A(n_4047),
.B(n_1573),
.C(n_1572),
.Y(n_4352)
);

AOI21xp5_ASAP7_75t_L g4353 ( 
.A1(n_4079),
.A2(n_4096),
.B(n_4093),
.Y(n_4353)
);

AND2x2_ASAP7_75t_L g4354 ( 
.A(n_4090),
.B(n_1574),
.Y(n_4354)
);

AO31x2_ASAP7_75t_L g4355 ( 
.A1(n_4069),
.A2(n_1577),
.A3(n_1582),
.B(n_1576),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4180),
.Y(n_4356)
);

OAI21x1_ASAP7_75t_L g4357 ( 
.A1(n_4232),
.A2(n_2303),
.B(n_2282),
.Y(n_4357)
);

AOI21xp33_ASAP7_75t_L g4358 ( 
.A1(n_4195),
.A2(n_4178),
.B(n_4043),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_SL g4359 ( 
.A(n_4225),
.B(n_1583),
.Y(n_4359)
);

INVx2_ASAP7_75t_L g4360 ( 
.A(n_4196),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4229),
.Y(n_4361)
);

NOR2xp33_ASAP7_75t_L g4362 ( 
.A(n_4129),
.B(n_1209),
.Y(n_4362)
);

AO31x2_ASAP7_75t_L g4363 ( 
.A1(n_4055),
.A2(n_1585),
.A3(n_1586),
.B(n_1584),
.Y(n_4363)
);

AOI21xp5_ASAP7_75t_L g4364 ( 
.A1(n_4108),
.A2(n_2306),
.B(n_2303),
.Y(n_4364)
);

OAI21x1_ASAP7_75t_L g4365 ( 
.A1(n_4192),
.A2(n_2316),
.B(n_2306),
.Y(n_4365)
);

OAI21x1_ASAP7_75t_L g4366 ( 
.A1(n_4193),
.A2(n_2316),
.B(n_2355),
.Y(n_4366)
);

AOI221xp5_ASAP7_75t_L g4367 ( 
.A1(n_4236),
.A2(n_1227),
.B1(n_1238),
.B2(n_1216),
.C(n_1214),
.Y(n_4367)
);

AO31x2_ASAP7_75t_L g4368 ( 
.A1(n_4126),
.A2(n_1589),
.A3(n_1590),
.B(n_1588),
.Y(n_4368)
);

AND2x6_ASAP7_75t_L g4369 ( 
.A(n_4253),
.B(n_1591),
.Y(n_4369)
);

OAI21x1_ASAP7_75t_L g4370 ( 
.A1(n_4239),
.A2(n_2398),
.B(n_2360),
.Y(n_4370)
);

OA22x2_ASAP7_75t_L g4371 ( 
.A1(n_4203),
.A2(n_1594),
.B1(n_1595),
.B2(n_1592),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_SL g4372 ( 
.A(n_4082),
.B(n_1596),
.Y(n_4372)
);

NOR2xp67_ASAP7_75t_SL g4373 ( 
.A(n_4121),
.B(n_1601),
.Y(n_4373)
);

BUFx2_ASAP7_75t_L g4374 ( 
.A(n_4246),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4202),
.Y(n_4375)
);

OAI21xp5_ASAP7_75t_L g4376 ( 
.A1(n_4258),
.A2(n_1604),
.B(n_1602),
.Y(n_4376)
);

NOR2xp33_ASAP7_75t_L g4377 ( 
.A(n_4095),
.B(n_1606),
.Y(n_4377)
);

OAI21x1_ASAP7_75t_L g4378 ( 
.A1(n_4248),
.A2(n_2398),
.B(n_2360),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_4077),
.B(n_4080),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4230),
.Y(n_4380)
);

AND2x6_ASAP7_75t_SL g4381 ( 
.A(n_4147),
.B(n_1607),
.Y(n_4381)
);

CKINVDCx5p33_ASAP7_75t_R g4382 ( 
.A(n_4013),
.Y(n_4382)
);

INVxp67_ASAP7_75t_SL g4383 ( 
.A(n_4146),
.Y(n_4383)
);

OAI21x1_ASAP7_75t_L g4384 ( 
.A1(n_4260),
.A2(n_2408),
.B(n_2399),
.Y(n_4384)
);

AOI21xp5_ASAP7_75t_L g4385 ( 
.A1(n_4086),
.A2(n_2204),
.B(n_2193),
.Y(n_4385)
);

BUFx8_ASAP7_75t_SL g4386 ( 
.A(n_4035),
.Y(n_4386)
);

AO32x2_ASAP7_75t_L g4387 ( 
.A1(n_4091),
.A2(n_5),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_4387)
);

A2O1A1Ixp33_ASAP7_75t_L g4388 ( 
.A1(n_4237),
.A2(n_1609),
.B(n_1613),
.C(n_1608),
.Y(n_4388)
);

HB1xp67_ASAP7_75t_L g4389 ( 
.A(n_4217),
.Y(n_4389)
);

BUFx2_ASAP7_75t_L g4390 ( 
.A(n_4246),
.Y(n_4390)
);

OA21x2_ASAP7_75t_L g4391 ( 
.A1(n_4054),
.A2(n_1616),
.B(n_1615),
.Y(n_4391)
);

AND2x4_ASAP7_75t_L g4392 ( 
.A(n_4253),
.B(n_638),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4027),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4038),
.Y(n_4394)
);

NAND2x1p5_ASAP7_75t_L g4395 ( 
.A(n_4070),
.B(n_2193),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4061),
.Y(n_4396)
);

NOR2xp33_ASAP7_75t_L g4397 ( 
.A(n_4131),
.B(n_1619),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4085),
.Y(n_4398)
);

NOR2xp67_ASAP7_75t_L g4399 ( 
.A(n_4133),
.B(n_1621),
.Y(n_4399)
);

OAI21x1_ASAP7_75t_L g4400 ( 
.A1(n_4266),
.A2(n_2408),
.B(n_2399),
.Y(n_4400)
);

OAI21x1_ASAP7_75t_L g4401 ( 
.A1(n_4270),
.A2(n_2440),
.B(n_1624),
.Y(n_4401)
);

OAI21xp5_ASAP7_75t_L g4402 ( 
.A1(n_4214),
.A2(n_1625),
.B(n_1623),
.Y(n_4402)
);

BUFx6f_ASAP7_75t_L g4403 ( 
.A(n_4244),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_SL g4404 ( 
.A(n_4158),
.B(n_4164),
.Y(n_4404)
);

OAI21x1_ASAP7_75t_L g4405 ( 
.A1(n_4072),
.A2(n_2440),
.B(n_1628),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4088),
.Y(n_4406)
);

AOI21xp5_ASAP7_75t_L g4407 ( 
.A1(n_4123),
.A2(n_2213),
.B(n_2204),
.Y(n_4407)
);

INVx4_ASAP7_75t_L g4408 ( 
.A(n_4031),
.Y(n_4408)
);

OAI22xp5_ASAP7_75t_L g4409 ( 
.A1(n_4168),
.A2(n_1632),
.B1(n_1635),
.B2(n_1626),
.Y(n_4409)
);

OAI21x1_ASAP7_75t_SL g4410 ( 
.A1(n_4020),
.A2(n_4115),
.B(n_4216),
.Y(n_4410)
);

O2A1O1Ixp5_ASAP7_75t_SL g4411 ( 
.A1(n_4234),
.A2(n_1645),
.B(n_1646),
.C(n_1640),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_L g4412 ( 
.A(n_4209),
.B(n_1649),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_4098),
.B(n_1653),
.Y(n_4413)
);

OAI21xp5_ASAP7_75t_L g4414 ( 
.A1(n_4039),
.A2(n_1662),
.B(n_1659),
.Y(n_4414)
);

OAI21x1_ASAP7_75t_L g4415 ( 
.A1(n_4052),
.A2(n_1664),
.B(n_1663),
.Y(n_4415)
);

INVx2_ASAP7_75t_L g4416 ( 
.A(n_4099),
.Y(n_4416)
);

AO31x2_ASAP7_75t_L g4417 ( 
.A1(n_4110),
.A2(n_1666),
.A3(n_1670),
.B(n_1665),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_SL g4418 ( 
.A(n_4119),
.B(n_1671),
.Y(n_4418)
);

NAND3xp33_ASAP7_75t_L g4419 ( 
.A(n_4241),
.B(n_1677),
.C(n_1676),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_L g4420 ( 
.A(n_4101),
.B(n_1679),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_L g4421 ( 
.A(n_4084),
.B(n_2005),
.Y(n_4421)
);

OAI21x1_ASAP7_75t_L g4422 ( 
.A1(n_4220),
.A2(n_2213),
.B(n_2204),
.Y(n_4422)
);

OAI21x1_ASAP7_75t_L g4423 ( 
.A1(n_4150),
.A2(n_2213),
.B(n_2204),
.Y(n_4423)
);

AOI21xp5_ASAP7_75t_L g4424 ( 
.A1(n_4044),
.A2(n_2214),
.B(n_2213),
.Y(n_4424)
);

NOR2xp33_ASAP7_75t_L g4425 ( 
.A(n_4151),
.B(n_639),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_SL g4426 ( 
.A(n_4128),
.B(n_2020),
.Y(n_4426)
);

AND2x4_ASAP7_75t_L g4427 ( 
.A(n_4234),
.B(n_640),
.Y(n_4427)
);

AO31x2_ASAP7_75t_L g4428 ( 
.A1(n_4105),
.A2(n_4042),
.A3(n_4089),
.B(n_4132),
.Y(n_4428)
);

NOR2xp33_ASAP7_75t_L g4429 ( 
.A(n_4152),
.B(n_4172),
.Y(n_4429)
);

NOR2x1_ASAP7_75t_SL g4430 ( 
.A(n_4203),
.B(n_4142),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_L g4431 ( 
.A(n_4107),
.B(n_2024),
.Y(n_4431)
);

OAI21xp33_ASAP7_75t_SL g4432 ( 
.A1(n_4118),
.A2(n_4),
.B(n_5),
.Y(n_4432)
);

BUFx2_ASAP7_75t_L g4433 ( 
.A(n_4268),
.Y(n_4433)
);

AO22x2_ASAP7_75t_L g4434 ( 
.A1(n_4028),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_4434)
);

BUFx3_ASAP7_75t_L g4435 ( 
.A(n_4122),
.Y(n_4435)
);

CKINVDCx5p33_ASAP7_75t_R g4436 ( 
.A(n_4191),
.Y(n_4436)
);

AOI21xp5_ASAP7_75t_L g4437 ( 
.A1(n_4169),
.A2(n_2221),
.B(n_2214),
.Y(n_4437)
);

BUFx3_ASAP7_75t_L g4438 ( 
.A(n_4144),
.Y(n_4438)
);

NOR2x1_ASAP7_75t_SL g4439 ( 
.A(n_4160),
.B(n_2214),
.Y(n_4439)
);

NAND3xp33_ASAP7_75t_L g4440 ( 
.A(n_4245),
.B(n_2028),
.C(n_2024),
.Y(n_4440)
);

OAI21xp5_ASAP7_75t_L g4441 ( 
.A1(n_4166),
.A2(n_1777),
.B(n_1895),
.Y(n_4441)
);

AO31x2_ASAP7_75t_L g4442 ( 
.A1(n_4130),
.A2(n_2221),
.A3(n_2226),
.B(n_2214),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_4109),
.B(n_2024),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_4137),
.B(n_2024),
.Y(n_4444)
);

NAND3xp33_ASAP7_75t_L g4445 ( 
.A(n_4182),
.B(n_2028),
.C(n_1989),
.Y(n_4445)
);

OAI21xp5_ASAP7_75t_L g4446 ( 
.A1(n_4219),
.A2(n_1898),
.B(n_1895),
.Y(n_4446)
);

NOR2xp33_ASAP7_75t_L g4447 ( 
.A(n_4198),
.B(n_641),
.Y(n_4447)
);

OAI22xp5_ASAP7_75t_L g4448 ( 
.A1(n_4159),
.A2(n_2221),
.B1(n_2231),
.B2(n_2226),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_4135),
.Y(n_4449)
);

AOI21xp5_ASAP7_75t_L g4450 ( 
.A1(n_4204),
.A2(n_2226),
.B(n_2221),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_L g4451 ( 
.A(n_4250),
.B(n_2028),
.Y(n_4451)
);

AOI21xp5_ASAP7_75t_L g4452 ( 
.A1(n_4199),
.A2(n_2231),
.B(n_2226),
.Y(n_4452)
);

NOR2xp33_ASAP7_75t_L g4453 ( 
.A(n_4157),
.B(n_642),
.Y(n_4453)
);

OA22x2_ASAP7_75t_L g4454 ( 
.A1(n_4139),
.A2(n_11),
.B1(n_7),
.B2(n_8),
.Y(n_4454)
);

NOR2xp67_ASAP7_75t_L g4455 ( 
.A(n_4058),
.B(n_645),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4148),
.Y(n_4456)
);

OAI21xp5_ASAP7_75t_L g4457 ( 
.A1(n_4173),
.A2(n_1898),
.B(n_1895),
.Y(n_4457)
);

CKINVDCx5p33_ASAP7_75t_R g4458 ( 
.A(n_4134),
.Y(n_4458)
);

INVx3_ASAP7_75t_L g4459 ( 
.A(n_4062),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4075),
.Y(n_4460)
);

AOI21xp5_ASAP7_75t_L g4461 ( 
.A1(n_4067),
.A2(n_2256),
.B(n_2231),
.Y(n_4461)
);

AOI21xp5_ASAP7_75t_L g4462 ( 
.A1(n_4176),
.A2(n_2256),
.B(n_2231),
.Y(n_4462)
);

BUFx2_ASAP7_75t_L g4463 ( 
.A(n_4268),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_SL g4464 ( 
.A(n_4177),
.B(n_2028),
.Y(n_4464)
);

BUFx2_ASAP7_75t_L g4465 ( 
.A(n_4269),
.Y(n_4465)
);

AOI21xp5_ASAP7_75t_L g4466 ( 
.A1(n_4227),
.A2(n_2269),
.B(n_2256),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4243),
.B(n_11),
.Y(n_4467)
);

OAI21x1_ASAP7_75t_L g4468 ( 
.A1(n_4189),
.A2(n_4125),
.B(n_4247),
.Y(n_4468)
);

OAI21xp33_ASAP7_75t_L g4469 ( 
.A1(n_4201),
.A2(n_1989),
.B(n_1988),
.Y(n_4469)
);

OAI21xp5_ASAP7_75t_L g4470 ( 
.A1(n_4256),
.A2(n_1898),
.B(n_1895),
.Y(n_4470)
);

AOI21x1_ASAP7_75t_L g4471 ( 
.A1(n_4264),
.A2(n_2269),
.B(n_2256),
.Y(n_4471)
);

HB1xp67_ASAP7_75t_L g4472 ( 
.A(n_4206),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4117),
.Y(n_4473)
);

OAI21x1_ASAP7_75t_L g4474 ( 
.A1(n_4251),
.A2(n_2279),
.B(n_2269),
.Y(n_4474)
);

AOI22xp5_ASAP7_75t_L g4475 ( 
.A1(n_4127),
.A2(n_1989),
.B1(n_1988),
.B2(n_1875),
.Y(n_4475)
);

BUFx2_ASAP7_75t_L g4476 ( 
.A(n_4231),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_L g4477 ( 
.A(n_4272),
.B(n_12),
.Y(n_4477)
);

OAI21x1_ASAP7_75t_L g4478 ( 
.A1(n_4221),
.A2(n_2279),
.B(n_2269),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_4188),
.B(n_12),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_4117),
.B(n_4208),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4226),
.Y(n_4481)
);

NAND2x1p5_ASAP7_75t_L g4482 ( 
.A(n_4070),
.B(n_2279),
.Y(n_4482)
);

BUFx6f_ASAP7_75t_L g4483 ( 
.A(n_4244),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_L g4484 ( 
.A(n_4208),
.B(n_13),
.Y(n_4484)
);

AND2x2_ASAP7_75t_L g4485 ( 
.A(n_4062),
.B(n_4063),
.Y(n_4485)
);

A2O1A1Ixp33_ASAP7_75t_L g4486 ( 
.A1(n_4261),
.A2(n_17),
.B(n_14),
.C(n_15),
.Y(n_4486)
);

BUFx6f_ASAP7_75t_L g4487 ( 
.A(n_4244),
.Y(n_4487)
);

AOI21xp5_ASAP7_75t_L g4488 ( 
.A1(n_4257),
.A2(n_4271),
.B(n_4262),
.Y(n_4488)
);

NOR2x1_ASAP7_75t_SL g4489 ( 
.A(n_4031),
.B(n_2279),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_4063),
.B(n_14),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_4184),
.B(n_15),
.Y(n_4491)
);

AND2x2_ASAP7_75t_L g4492 ( 
.A(n_4240),
.B(n_646),
.Y(n_4492)
);

OAI21xp5_ASAP7_75t_L g4493 ( 
.A1(n_4255),
.A2(n_1925),
.B(n_1898),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_L g4494 ( 
.A(n_4153),
.B(n_17),
.Y(n_4494)
);

HB1xp67_ASAP7_75t_L g4495 ( 
.A(n_4138),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_4112),
.Y(n_4496)
);

AO31x2_ASAP7_75t_L g4497 ( 
.A1(n_4235),
.A2(n_2295),
.A3(n_2300),
.B(n_2289),
.Y(n_4497)
);

INVx2_ASAP7_75t_L g4498 ( 
.A(n_4112),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_4210),
.B(n_18),
.Y(n_4499)
);

AOI21xp33_ASAP7_75t_L g4500 ( 
.A1(n_4254),
.A2(n_1989),
.B(n_2289),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4138),
.B(n_650),
.Y(n_4501)
);

OAI21x1_ASAP7_75t_L g4502 ( 
.A1(n_4076),
.A2(n_2295),
.B(n_2289),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4106),
.Y(n_4503)
);

INVx2_ASAP7_75t_SL g4504 ( 
.A(n_4179),
.Y(n_4504)
);

OAI21x1_ASAP7_75t_L g4505 ( 
.A1(n_4106),
.A2(n_2295),
.B(n_2289),
.Y(n_4505)
);

AND2x2_ASAP7_75t_SL g4506 ( 
.A(n_4058),
.B(n_1874),
.Y(n_4506)
);

OAI21x1_ASAP7_75t_L g4507 ( 
.A1(n_4106),
.A2(n_4222),
.B(n_4207),
.Y(n_4507)
);

OAI21xp5_ASAP7_75t_L g4508 ( 
.A1(n_4163),
.A2(n_1937),
.B(n_1925),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_SL g4509 ( 
.A(n_4171),
.B(n_1874),
.Y(n_4509)
);

INVx3_ASAP7_75t_L g4510 ( 
.A(n_4165),
.Y(n_4510)
);

OAI21x1_ASAP7_75t_SL g4511 ( 
.A1(n_4165),
.A2(n_4179),
.B(n_4041),
.Y(n_4511)
);

INVx1_ASAP7_75t_L g4512 ( 
.A(n_4031),
.Y(n_4512)
);

AND2x4_ASAP7_75t_L g4513 ( 
.A(n_4041),
.B(n_651),
.Y(n_4513)
);

AOI21xp5_ASAP7_75t_L g4514 ( 
.A1(n_4103),
.A2(n_2300),
.B(n_2295),
.Y(n_4514)
);

AOI22x1_ASAP7_75t_L g4515 ( 
.A1(n_4041),
.A2(n_2314),
.B1(n_2300),
.B2(n_2319),
.Y(n_4515)
);

AOI21x1_ASAP7_75t_L g4516 ( 
.A1(n_4154),
.A2(n_2314),
.B(n_2300),
.Y(n_4516)
);

OAI21x1_ASAP7_75t_L g4517 ( 
.A1(n_4102),
.A2(n_2314),
.B(n_1875),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_L g4518 ( 
.A(n_4102),
.B(n_18),
.Y(n_4518)
);

AO31x2_ASAP7_75t_L g4519 ( 
.A1(n_4102),
.A2(n_2314),
.A3(n_656),
.B(n_659),
.Y(n_4519)
);

NOR2xp33_ASAP7_75t_L g4520 ( 
.A(n_4116),
.B(n_655),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_4116),
.B(n_19),
.Y(n_4521)
);

AOI21xp5_ASAP7_75t_L g4522 ( 
.A1(n_4116),
.A2(n_4140),
.B(n_4124),
.Y(n_4522)
);

OAI22xp5_ASAP7_75t_L g4523 ( 
.A1(n_4124),
.A2(n_2328),
.B1(n_2332),
.B2(n_2319),
.Y(n_4523)
);

AOI21xp5_ASAP7_75t_L g4524 ( 
.A1(n_4124),
.A2(n_2328),
.B(n_2319),
.Y(n_4524)
);

OAI21x1_ASAP7_75t_L g4525 ( 
.A1(n_4140),
.A2(n_1875),
.B(n_1874),
.Y(n_4525)
);

OAI21x1_ASAP7_75t_L g4526 ( 
.A1(n_4140),
.A2(n_1875),
.B(n_1874),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_SL g4527 ( 
.A(n_4282),
.B(n_1925),
.Y(n_4527)
);

INVx2_ASAP7_75t_L g4528 ( 
.A(n_4326),
.Y(n_4528)
);

AO21x1_ASAP7_75t_L g4529 ( 
.A1(n_4311),
.A2(n_20),
.B(n_21),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4285),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_4339),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_4279),
.Y(n_4532)
);

AND2x2_ASAP7_75t_L g4533 ( 
.A(n_4287),
.B(n_20),
.Y(n_4533)
);

AOI21xp5_ASAP7_75t_L g4534 ( 
.A1(n_4353),
.A2(n_2328),
.B(n_2319),
.Y(n_4534)
);

NAND2xp5_ASAP7_75t_L g4535 ( 
.A(n_4313),
.B(n_21),
.Y(n_4535)
);

AOI21xp5_ASAP7_75t_L g4536 ( 
.A1(n_4333),
.A2(n_2332),
.B(n_2328),
.Y(n_4536)
);

NAND2x1p5_ASAP7_75t_L g4537 ( 
.A(n_4345),
.B(n_2332),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_4312),
.B(n_22),
.Y(n_4538)
);

AND2x2_ASAP7_75t_L g4539 ( 
.A(n_4383),
.B(n_23),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4389),
.B(n_23),
.Y(n_4540)
);

AND2x2_ASAP7_75t_L g4541 ( 
.A(n_4322),
.B(n_24),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4292),
.Y(n_4542)
);

BUFx2_ASAP7_75t_L g4543 ( 
.A(n_4294),
.Y(n_4543)
);

AOI22xp33_ASAP7_75t_L g4544 ( 
.A1(n_4349),
.A2(n_1937),
.B1(n_1940),
.B2(n_1925),
.Y(n_4544)
);

AOI21xp5_ASAP7_75t_L g4545 ( 
.A1(n_4457),
.A2(n_4302),
.B(n_4508),
.Y(n_4545)
);

BUFx2_ASAP7_75t_L g4546 ( 
.A(n_4348),
.Y(n_4546)
);

AND2x2_ASAP7_75t_L g4547 ( 
.A(n_4485),
.B(n_24),
.Y(n_4547)
);

CKINVDCx5p33_ASAP7_75t_R g4548 ( 
.A(n_4386),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4314),
.Y(n_4549)
);

INVx3_ASAP7_75t_L g4550 ( 
.A(n_4473),
.Y(n_4550)
);

INVx2_ASAP7_75t_SL g4551 ( 
.A(n_4290),
.Y(n_4551)
);

NAND3xp33_ASAP7_75t_L g4552 ( 
.A(n_4295),
.B(n_1940),
.C(n_1937),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_4321),
.Y(n_4553)
);

BUFx2_ASAP7_75t_L g4554 ( 
.A(n_4495),
.Y(n_4554)
);

AND2x4_ASAP7_75t_L g4555 ( 
.A(n_4503),
.B(n_662),
.Y(n_4555)
);

BUFx3_ASAP7_75t_L g4556 ( 
.A(n_4458),
.Y(n_4556)
);

AOI22xp33_ASAP7_75t_L g4557 ( 
.A1(n_4358),
.A2(n_1940),
.B1(n_1941),
.B2(n_1937),
.Y(n_4557)
);

CKINVDCx5p33_ASAP7_75t_R g4558 ( 
.A(n_4382),
.Y(n_4558)
);

OAI21xp33_ASAP7_75t_L g4559 ( 
.A1(n_4494),
.A2(n_25),
.B(n_26),
.Y(n_4559)
);

AND2x4_ASAP7_75t_L g4560 ( 
.A(n_4345),
.B(n_665),
.Y(n_4560)
);

AND2x4_ASAP7_75t_L g4561 ( 
.A(n_4345),
.B(n_668),
.Y(n_4561)
);

AOI21xp5_ASAP7_75t_L g4562 ( 
.A1(n_4493),
.A2(n_2333),
.B(n_2332),
.Y(n_4562)
);

NOR2xp33_ASAP7_75t_L g4563 ( 
.A(n_4381),
.B(n_4379),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4299),
.B(n_26),
.Y(n_4564)
);

AOI21xp5_ASAP7_75t_L g4565 ( 
.A1(n_4452),
.A2(n_2347),
.B(n_2333),
.Y(n_4565)
);

BUFx12f_ASAP7_75t_L g4566 ( 
.A(n_4436),
.Y(n_4566)
);

AND2x2_ASAP7_75t_L g4567 ( 
.A(n_4330),
.B(n_28),
.Y(n_4567)
);

NAND2xp5_ASAP7_75t_L g4568 ( 
.A(n_4286),
.B(n_28),
.Y(n_4568)
);

BUFx12f_ASAP7_75t_L g4569 ( 
.A(n_4290),
.Y(n_4569)
);

NAND2xp5_ASAP7_75t_L g4570 ( 
.A(n_4360),
.B(n_29),
.Y(n_4570)
);

AND2x4_ASAP7_75t_L g4571 ( 
.A(n_4356),
.B(n_669),
.Y(n_4571)
);

NAND2xp5_ASAP7_75t_L g4572 ( 
.A(n_4375),
.B(n_4393),
.Y(n_4572)
);

NAND2x1p5_ASAP7_75t_L g4573 ( 
.A(n_4509),
.B(n_2333),
.Y(n_4573)
);

NOR2xp67_ASAP7_75t_L g4574 ( 
.A(n_4316),
.B(n_30),
.Y(n_4574)
);

INVx2_ASAP7_75t_SL g4575 ( 
.A(n_4290),
.Y(n_4575)
);

INVx5_ASAP7_75t_L g4576 ( 
.A(n_4369),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4361),
.Y(n_4577)
);

OAI22xp5_ASAP7_75t_L g4578 ( 
.A1(n_4404),
.A2(n_2347),
.B1(n_2372),
.B2(n_2333),
.Y(n_4578)
);

AO32x1_ASAP7_75t_L g4579 ( 
.A1(n_4460),
.A2(n_34),
.A3(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_4579)
);

AND2x4_ASAP7_75t_L g4580 ( 
.A(n_4380),
.B(n_670),
.Y(n_4580)
);

AOI21xp5_ASAP7_75t_L g4581 ( 
.A1(n_4288),
.A2(n_4446),
.B(n_4470),
.Y(n_4581)
);

AOI21xp5_ASAP7_75t_L g4582 ( 
.A1(n_4303),
.A2(n_2372),
.B(n_2347),
.Y(n_4582)
);

NOR2xp33_ASAP7_75t_L g4583 ( 
.A(n_4362),
.B(n_32),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_L g4584 ( 
.A(n_4394),
.B(n_35),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4396),
.Y(n_4585)
);

INVx2_ASAP7_75t_L g4586 ( 
.A(n_4398),
.Y(n_4586)
);

NOR2xp33_ASAP7_75t_L g4587 ( 
.A(n_4281),
.B(n_36),
.Y(n_4587)
);

CKINVDCx20_ASAP7_75t_R g4588 ( 
.A(n_4435),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_4406),
.B(n_36),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4416),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4449),
.Y(n_4591)
);

AO21x2_ASAP7_75t_L g4592 ( 
.A1(n_4424),
.A2(n_37),
.B(n_39),
.Y(n_4592)
);

AOI22xp33_ASAP7_75t_L g4593 ( 
.A1(n_4454),
.A2(n_1941),
.B1(n_1940),
.B2(n_1715),
.Y(n_4593)
);

INVx2_ASAP7_75t_L g4594 ( 
.A(n_4291),
.Y(n_4594)
);

INVx3_ASAP7_75t_L g4595 ( 
.A(n_4408),
.Y(n_4595)
);

INVxp67_ASAP7_75t_L g4596 ( 
.A(n_4472),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4456),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_4387),
.Y(n_4598)
);

NOR2xp67_ASAP7_75t_L g4599 ( 
.A(n_4488),
.B(n_39),
.Y(n_4599)
);

HB1xp67_ASAP7_75t_L g4600 ( 
.A(n_4336),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_4480),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4512),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_4284),
.B(n_40),
.Y(n_4603)
);

OAI22xp5_ASAP7_75t_L g4604 ( 
.A1(n_4429),
.A2(n_2347),
.B1(n_2375),
.B2(n_2372),
.Y(n_4604)
);

BUFx6f_ASAP7_75t_SL g4605 ( 
.A(n_4504),
.Y(n_4605)
);

NAND2xp5_ASAP7_75t_L g4606 ( 
.A(n_4354),
.B(n_40),
.Y(n_4606)
);

NOR2xp33_ASAP7_75t_L g4607 ( 
.A(n_4280),
.B(n_41),
.Y(n_4607)
);

INVx2_ASAP7_75t_SL g4608 ( 
.A(n_4403),
.Y(n_4608)
);

BUFx6f_ASAP7_75t_L g4609 ( 
.A(n_4310),
.Y(n_4609)
);

AND2x2_ASAP7_75t_L g4610 ( 
.A(n_4275),
.B(n_41),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4387),
.Y(n_4611)
);

NOR2xp33_ASAP7_75t_L g4612 ( 
.A(n_4377),
.B(n_42),
.Y(n_4612)
);

OR2x2_ASAP7_75t_L g4613 ( 
.A(n_4417),
.B(n_42),
.Y(n_4613)
);

OAI22xp5_ASAP7_75t_L g4614 ( 
.A1(n_4499),
.A2(n_4453),
.B1(n_4289),
.B2(n_4486),
.Y(n_4614)
);

OAI21x1_ASAP7_75t_L g4615 ( 
.A1(n_4385),
.A2(n_4276),
.B(n_4315),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4387),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4434),
.Y(n_4617)
);

AOI222xp33_ASAP7_75t_L g4618 ( 
.A1(n_4402),
.A2(n_73),
.B1(n_54),
.B2(n_84),
.C1(n_64),
.C2(n_43),
.Y(n_4618)
);

O2A1O1Ixp33_ASAP7_75t_SL g4619 ( 
.A1(n_4359),
.A2(n_54),
.B(n_64),
.C(n_43),
.Y(n_4619)
);

AND2x2_ASAP7_75t_SL g4620 ( 
.A(n_4300),
.B(n_45),
.Y(n_4620)
);

INVx4_ASAP7_75t_SL g4621 ( 
.A(n_4369),
.Y(n_4621)
);

AND2x2_ASAP7_75t_L g4622 ( 
.A(n_4275),
.B(n_46),
.Y(n_4622)
);

AND2x6_ASAP7_75t_L g4623 ( 
.A(n_4459),
.B(n_2372),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_4323),
.B(n_46),
.Y(n_4624)
);

AOI21xp33_ASAP7_75t_SL g4625 ( 
.A1(n_4397),
.A2(n_47),
.B(n_49),
.Y(n_4625)
);

NOR3xp33_ASAP7_75t_L g4626 ( 
.A(n_4432),
.B(n_49),
.C(n_50),
.Y(n_4626)
);

NOR2xp33_ASAP7_75t_SL g4627 ( 
.A(n_4296),
.B(n_1941),
.Y(n_4627)
);

NAND2xp5_ASAP7_75t_SL g4628 ( 
.A(n_4351),
.B(n_1941),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_4459),
.Y(n_4629)
);

OR2x2_ASAP7_75t_L g4630 ( 
.A(n_4417),
.B(n_51),
.Y(n_4630)
);

INVx3_ASAP7_75t_L g4631 ( 
.A(n_4408),
.Y(n_4631)
);

OR2x2_ASAP7_75t_L g4632 ( 
.A(n_4417),
.B(n_51),
.Y(n_4632)
);

HB1xp67_ASAP7_75t_L g4633 ( 
.A(n_4428),
.Y(n_4633)
);

INVx2_ASAP7_75t_L g4634 ( 
.A(n_4496),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_L g4635 ( 
.A(n_4347),
.B(n_53),
.Y(n_4635)
);

AND2x4_ASAP7_75t_L g4636 ( 
.A(n_4297),
.B(n_671),
.Y(n_4636)
);

NAND2xp33_ASAP7_75t_SL g4637 ( 
.A(n_4310),
.B(n_53),
.Y(n_4637)
);

NOR2xp33_ASAP7_75t_L g4638 ( 
.A(n_4412),
.B(n_55),
.Y(n_4638)
);

O2A1O1Ixp33_ASAP7_75t_SL g4639 ( 
.A1(n_4467),
.A2(n_67),
.B(n_75),
.C(n_55),
.Y(n_4639)
);

OAI21xp5_ASAP7_75t_L g4640 ( 
.A1(n_4331),
.A2(n_2030),
.B(n_2006),
.Y(n_4640)
);

CKINVDCx5p33_ASAP7_75t_R g4641 ( 
.A(n_4438),
.Y(n_4641)
);

BUFx2_ASAP7_75t_L g4642 ( 
.A(n_4465),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4434),
.Y(n_4643)
);

INVx2_ASAP7_75t_L g4644 ( 
.A(n_4498),
.Y(n_4644)
);

BUFx3_ASAP7_75t_L g4645 ( 
.A(n_4340),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4304),
.B(n_56),
.Y(n_4646)
);

INVx5_ASAP7_75t_L g4647 ( 
.A(n_4369),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4403),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4355),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4325),
.B(n_56),
.Y(n_4650)
);

AND2x2_ASAP7_75t_L g4651 ( 
.A(n_4297),
.B(n_58),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_4476),
.B(n_58),
.Y(n_4652)
);

NAND2xp5_ASAP7_75t_L g4653 ( 
.A(n_4344),
.B(n_60),
.Y(n_4653)
);

OAI22xp5_ASAP7_75t_L g4654 ( 
.A1(n_4399),
.A2(n_2379),
.B1(n_2391),
.B2(n_2375),
.Y(n_4654)
);

O2A1O1Ixp33_ASAP7_75t_L g4655 ( 
.A1(n_4306),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_4655)
);

INVx4_ASAP7_75t_L g4656 ( 
.A(n_4369),
.Y(n_4656)
);

NOR2xp33_ASAP7_75t_L g4657 ( 
.A(n_4477),
.B(n_61),
.Y(n_4657)
);

NOR2xp33_ASAP7_75t_L g4658 ( 
.A(n_4479),
.B(n_66),
.Y(n_4658)
);

BUFx2_ASAP7_75t_L g4659 ( 
.A(n_4374),
.Y(n_4659)
);

OAI22xp5_ASAP7_75t_L g4660 ( 
.A1(n_4371),
.A2(n_2379),
.B1(n_2391),
.B2(n_2375),
.Y(n_4660)
);

INVx1_ASAP7_75t_SL g4661 ( 
.A(n_4390),
.Y(n_4661)
);

INVxp67_ASAP7_75t_SL g4662 ( 
.A(n_4274),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4490),
.B(n_66),
.Y(n_4663)
);

INVx2_ASAP7_75t_L g4664 ( 
.A(n_4403),
.Y(n_4664)
);

INVx2_ASAP7_75t_SL g4665 ( 
.A(n_4483),
.Y(n_4665)
);

A2O1A1Ixp33_ASAP7_75t_L g4666 ( 
.A1(n_4447),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_4666)
);

O2A1O1Ixp33_ASAP7_75t_L g4667 ( 
.A1(n_4414),
.A2(n_4491),
.B(n_4320),
.C(n_4328),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_L g4668 ( 
.A(n_4428),
.B(n_68),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4355),
.Y(n_4669)
);

AOI22xp5_ASAP7_75t_L g4670 ( 
.A1(n_4425),
.A2(n_2030),
.B1(n_2006),
.B2(n_2375),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4355),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4428),
.B(n_70),
.Y(n_4672)
);

AND2x4_ASAP7_75t_L g4673 ( 
.A(n_4430),
.B(n_672),
.Y(n_4673)
);

BUFx6f_ASAP7_75t_L g4674 ( 
.A(n_4310),
.Y(n_4674)
);

BUFx6f_ASAP7_75t_L g4675 ( 
.A(n_4483),
.Y(n_4675)
);

BUFx3_ASAP7_75t_L g4676 ( 
.A(n_4433),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4368),
.Y(n_4677)
);

CKINVDCx20_ASAP7_75t_R g4678 ( 
.A(n_4463),
.Y(n_4678)
);

AOI21xp5_ASAP7_75t_L g4679 ( 
.A1(n_4450),
.A2(n_4441),
.B(n_4437),
.Y(n_4679)
);

INVx2_ASAP7_75t_SL g4680 ( 
.A(n_4483),
.Y(n_4680)
);

AOI21xp5_ASAP7_75t_L g4681 ( 
.A1(n_4466),
.A2(n_2391),
.B(n_2379),
.Y(n_4681)
);

OR2x2_ASAP7_75t_L g4682 ( 
.A(n_4368),
.B(n_70),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_4368),
.Y(n_4683)
);

INVxp67_ASAP7_75t_SL g4684 ( 
.A(n_4391),
.Y(n_4684)
);

INVxp67_ASAP7_75t_L g4685 ( 
.A(n_4487),
.Y(n_4685)
);

BUFx6f_ASAP7_75t_L g4686 ( 
.A(n_4487),
.Y(n_4686)
);

OA21x2_ASAP7_75t_L g4687 ( 
.A1(n_4319),
.A2(n_71),
.B(n_72),
.Y(n_4687)
);

AOI21xp5_ASAP7_75t_L g4688 ( 
.A1(n_4308),
.A2(n_2391),
.B(n_2379),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4415),
.Y(n_4689)
);

BUFx2_ASAP7_75t_L g4690 ( 
.A(n_4487),
.Y(n_4690)
);

BUFx3_ASAP7_75t_L g4691 ( 
.A(n_4511),
.Y(n_4691)
);

AND2x2_ASAP7_75t_L g4692 ( 
.A(n_4518),
.B(n_71),
.Y(n_4692)
);

AOI21xp5_ASAP7_75t_L g4693 ( 
.A1(n_4462),
.A2(n_2400),
.B(n_2397),
.Y(n_4693)
);

INVx2_ASAP7_75t_SL g4694 ( 
.A(n_4510),
.Y(n_4694)
);

BUFx12f_ASAP7_75t_L g4695 ( 
.A(n_4296),
.Y(n_4695)
);

CKINVDCx5p33_ASAP7_75t_R g4696 ( 
.A(n_4522),
.Y(n_4696)
);

AND2x4_ASAP7_75t_L g4697 ( 
.A(n_4519),
.B(n_676),
.Y(n_4697)
);

NAND2xp5_ASAP7_75t_SL g4698 ( 
.A(n_4298),
.B(n_2006),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_L g4699 ( 
.A(n_4484),
.B(n_73),
.Y(n_4699)
);

OR2x2_ASAP7_75t_L g4700 ( 
.A(n_4413),
.B(n_74),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4363),
.Y(n_4701)
);

INVx3_ASAP7_75t_L g4702 ( 
.A(n_4427),
.Y(n_4702)
);

INVx3_ASAP7_75t_L g4703 ( 
.A(n_4427),
.Y(n_4703)
);

AOI22xp33_ASAP7_75t_L g4704 ( 
.A1(n_4481),
.A2(n_1715),
.B1(n_1694),
.B2(n_2006),
.Y(n_4704)
);

O2A1O1Ixp33_ASAP7_75t_L g4705 ( 
.A1(n_4327),
.A2(n_79),
.B(n_76),
.C(n_77),
.Y(n_4705)
);

AOI21xp5_ASAP7_75t_L g4706 ( 
.A1(n_4440),
.A2(n_2400),
.B(n_2397),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_L g4707 ( 
.A(n_4420),
.B(n_77),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4363),
.Y(n_4708)
);

AOI21xp5_ASAP7_75t_L g4709 ( 
.A1(n_4391),
.A2(n_2400),
.B(n_2397),
.Y(n_4709)
);

BUFx2_ASAP7_75t_L g4710 ( 
.A(n_4519),
.Y(n_4710)
);

BUFx2_ASAP7_75t_L g4711 ( 
.A(n_4519),
.Y(n_4711)
);

AO32x1_ASAP7_75t_L g4712 ( 
.A1(n_4448),
.A2(n_83),
.A3(n_79),
.B1(n_80),
.B2(n_84),
.Y(n_4712)
);

NAND2xp5_ASAP7_75t_L g4713 ( 
.A(n_4451),
.B(n_83),
.Y(n_4713)
);

BUFx3_ASAP7_75t_L g4714 ( 
.A(n_4392),
.Y(n_4714)
);

OR2x2_ASAP7_75t_L g4715 ( 
.A(n_4426),
.B(n_86),
.Y(n_4715)
);

CKINVDCx20_ASAP7_75t_R g4716 ( 
.A(n_4501),
.Y(n_4716)
);

AOI21xp5_ASAP7_75t_L g4717 ( 
.A1(n_4407),
.A2(n_2400),
.B(n_2397),
.Y(n_4717)
);

INVx2_ASAP7_75t_SL g4718 ( 
.A(n_4513),
.Y(n_4718)
);

AND2x4_ASAP7_75t_L g4719 ( 
.A(n_4392),
.B(n_4513),
.Y(n_4719)
);

OR2x2_ASAP7_75t_L g4720 ( 
.A(n_4421),
.B(n_86),
.Y(n_4720)
);

NOR3xp33_ASAP7_75t_L g4721 ( 
.A(n_4376),
.B(n_87),
.C(n_88),
.Y(n_4721)
);

CKINVDCx20_ASAP7_75t_R g4722 ( 
.A(n_4492),
.Y(n_4722)
);

OR2x2_ASAP7_75t_L g4723 ( 
.A(n_4521),
.B(n_88),
.Y(n_4723)
);

INVx2_ASAP7_75t_SL g4724 ( 
.A(n_4307),
.Y(n_4724)
);

AND2x2_ASAP7_75t_L g4725 ( 
.A(n_4520),
.B(n_89),
.Y(n_4725)
);

INVx5_ASAP7_75t_L g4726 ( 
.A(n_4439),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4352),
.B(n_90),
.Y(n_4727)
);

AND2x2_ASAP7_75t_L g4728 ( 
.A(n_4309),
.B(n_90),
.Y(n_4728)
);

A2O1A1Ixp33_ASAP7_75t_L g4729 ( 
.A1(n_4507),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_4729)
);

BUFx2_ASAP7_75t_L g4730 ( 
.A(n_4442),
.Y(n_4730)
);

AOI22xp33_ASAP7_75t_SL g4731 ( 
.A1(n_4346),
.A2(n_95),
.B1(n_92),
.B2(n_94),
.Y(n_4731)
);

AOI21xp5_ASAP7_75t_L g4732 ( 
.A1(n_4332),
.A2(n_2433),
.B(n_2412),
.Y(n_4732)
);

INVx5_ASAP7_75t_L g4733 ( 
.A(n_4489),
.Y(n_4733)
);

AOI222xp33_ASAP7_75t_L g4734 ( 
.A1(n_4367),
.A2(n_96),
.B1(n_98),
.B2(n_94),
.C1(n_95),
.C2(n_97),
.Y(n_4734)
);

OAI21xp33_ASAP7_75t_L g4735 ( 
.A1(n_4419),
.A2(n_97),
.B(n_99),
.Y(n_4735)
);

INVx4_ASAP7_75t_L g4736 ( 
.A(n_4506),
.Y(n_4736)
);

A2O1A1Ixp33_ASAP7_75t_SL g4737 ( 
.A1(n_4373),
.A2(n_104),
.B(n_101),
.C(n_103),
.Y(n_4737)
);

CKINVDCx5p33_ASAP7_75t_R g4738 ( 
.A(n_4409),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4363),
.Y(n_4739)
);

INVx2_ASAP7_75t_L g4740 ( 
.A(n_4442),
.Y(n_4740)
);

INVxp67_ASAP7_75t_L g4741 ( 
.A(n_4372),
.Y(n_4741)
);

CKINVDCx20_ASAP7_75t_R g4742 ( 
.A(n_4343),
.Y(n_4742)
);

OR2x2_ASAP7_75t_L g4743 ( 
.A(n_4431),
.B(n_104),
.Y(n_4743)
);

INVxp67_ASAP7_75t_L g4744 ( 
.A(n_4418),
.Y(n_4744)
);

INVx2_ASAP7_75t_SL g4745 ( 
.A(n_4395),
.Y(n_4745)
);

INVx2_ASAP7_75t_L g4746 ( 
.A(n_4442),
.Y(n_4746)
);

AOI22xp33_ASAP7_75t_L g4747 ( 
.A1(n_4410),
.A2(n_1715),
.B1(n_1694),
.B2(n_2030),
.Y(n_4747)
);

NOR2xp33_ASAP7_75t_L g4748 ( 
.A(n_4388),
.B(n_105),
.Y(n_4748)
);

INVx3_ASAP7_75t_L g4749 ( 
.A(n_4505),
.Y(n_4749)
);

NOR2xp33_ASAP7_75t_R g4750 ( 
.A(n_4516),
.B(n_4471),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4309),
.B(n_106),
.Y(n_4751)
);

INVx2_ASAP7_75t_L g4752 ( 
.A(n_4497),
.Y(n_4752)
);

AND2x2_ASAP7_75t_L g4753 ( 
.A(n_4497),
.B(n_107),
.Y(n_4753)
);

HB1xp67_ASAP7_75t_L g4754 ( 
.A(n_4497),
.Y(n_4754)
);

AOI21xp5_ASAP7_75t_L g4755 ( 
.A1(n_4278),
.A2(n_4464),
.B(n_4469),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_L g4756 ( 
.A(n_4318),
.B(n_4283),
.Y(n_4756)
);

AOI221x1_ASAP7_75t_L g4757 ( 
.A1(n_4461),
.A2(n_111),
.B1(n_108),
.B2(n_109),
.C(n_112),
.Y(n_4757)
);

BUFx3_ASAP7_75t_L g4758 ( 
.A(n_4482),
.Y(n_4758)
);

BUFx4_ASAP7_75t_SL g4759 ( 
.A(n_4445),
.Y(n_4759)
);

AND2x2_ASAP7_75t_L g4760 ( 
.A(n_4468),
.B(n_108),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4443),
.Y(n_4761)
);

AOI21xp5_ASAP7_75t_L g4762 ( 
.A1(n_4364),
.A2(n_2433),
.B(n_2412),
.Y(n_4762)
);

HB1xp67_ASAP7_75t_L g4763 ( 
.A(n_4305),
.Y(n_4763)
);

BUFx3_ASAP7_75t_L g4764 ( 
.A(n_4338),
.Y(n_4764)
);

OAI21x1_ASAP7_75t_L g4765 ( 
.A1(n_4342),
.A2(n_681),
.B(n_678),
.Y(n_4765)
);

INVx2_ASAP7_75t_SL g4766 ( 
.A(n_4502),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_4444),
.B(n_112),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4305),
.Y(n_4768)
);

INVx3_ASAP7_75t_L g4769 ( 
.A(n_4517),
.Y(n_4769)
);

AOI21xp33_ASAP7_75t_SL g4770 ( 
.A1(n_4475),
.A2(n_114),
.B(n_116),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4305),
.Y(n_4771)
);

CKINVDCx5p33_ASAP7_75t_R g4772 ( 
.A(n_4524),
.Y(n_4772)
);

AND2x4_ASAP7_75t_L g4773 ( 
.A(n_4455),
.B(n_684),
.Y(n_4773)
);

INVx1_ASAP7_75t_SL g4774 ( 
.A(n_4514),
.Y(n_4774)
);

AND2x4_ASAP7_75t_L g4775 ( 
.A(n_4525),
.B(n_4526),
.Y(n_4775)
);

BUFx2_ASAP7_75t_SL g4776 ( 
.A(n_4588),
.Y(n_4776)
);

INVx2_ASAP7_75t_L g4777 ( 
.A(n_4602),
.Y(n_4777)
);

OAI22xp5_ASAP7_75t_L g4778 ( 
.A1(n_4742),
.A2(n_4515),
.B1(n_4523),
.B2(n_4335),
.Y(n_4778)
);

HB1xp67_ASAP7_75t_L g4779 ( 
.A(n_4546),
.Y(n_4779)
);

OAI22xp33_ASAP7_75t_L g4780 ( 
.A1(n_4614),
.A2(n_4341),
.B1(n_4500),
.B2(n_4277),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4530),
.Y(n_4781)
);

AOI22xp5_ASAP7_75t_L g4782 ( 
.A1(n_4721),
.A2(n_4474),
.B1(n_4422),
.B2(n_4423),
.Y(n_4782)
);

NAND2x1p5_ASAP7_75t_L g4783 ( 
.A(n_4576),
.B(n_4405),
.Y(n_4783)
);

OAI22xp5_ASAP7_75t_L g4784 ( 
.A1(n_4738),
.A2(n_4277),
.B1(n_4411),
.B2(n_4478),
.Y(n_4784)
);

CKINVDCx20_ASAP7_75t_R g4785 ( 
.A(n_4548),
.Y(n_4785)
);

INVx6_ASAP7_75t_L g4786 ( 
.A(n_4566),
.Y(n_4786)
);

HB1xp67_ASAP7_75t_L g4787 ( 
.A(n_4554),
.Y(n_4787)
);

AOI22xp33_ASAP7_75t_L g4788 ( 
.A1(n_4618),
.A2(n_4401),
.B1(n_4317),
.B2(n_4324),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4530),
.Y(n_4789)
);

CKINVDCx11_ASAP7_75t_R g4790 ( 
.A(n_4678),
.Y(n_4790)
);

INVx5_ASAP7_75t_L g4791 ( 
.A(n_4728),
.Y(n_4791)
);

AOI22xp33_ASAP7_75t_L g4792 ( 
.A1(n_4583),
.A2(n_4734),
.B1(n_4529),
.B2(n_4559),
.Y(n_4792)
);

INVx1_ASAP7_75t_SL g4793 ( 
.A(n_4543),
.Y(n_4793)
);

AOI22xp33_ASAP7_75t_L g4794 ( 
.A1(n_4626),
.A2(n_4334),
.B1(n_4329),
.B2(n_4350),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4542),
.Y(n_4795)
);

INVx8_ASAP7_75t_L g4796 ( 
.A(n_4569),
.Y(n_4796)
);

INVxp67_ASAP7_75t_SL g4797 ( 
.A(n_4633),
.Y(n_4797)
);

INVx4_ASAP7_75t_L g4798 ( 
.A(n_4696),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4549),
.Y(n_4799)
);

OAI22xp5_ASAP7_75t_L g4800 ( 
.A1(n_4620),
.A2(n_4277),
.B1(n_4301),
.B2(n_117),
.Y(n_4800)
);

INVx1_ASAP7_75t_SL g4801 ( 
.A(n_4642),
.Y(n_4801)
);

AOI22xp33_ASAP7_75t_SL g4802 ( 
.A1(n_4748),
.A2(n_4357),
.B1(n_4378),
.B2(n_4370),
.Y(n_4802)
);

INVx2_ASAP7_75t_L g4803 ( 
.A(n_4553),
.Y(n_4803)
);

AOI22xp33_ASAP7_75t_L g4804 ( 
.A1(n_4612),
.A2(n_4365),
.B1(n_4366),
.B2(n_4337),
.Y(n_4804)
);

INVxp67_ASAP7_75t_SL g4805 ( 
.A(n_4596),
.Y(n_4805)
);

AOI22xp33_ASAP7_75t_L g4806 ( 
.A1(n_4735),
.A2(n_4400),
.B1(n_4384),
.B2(n_1715),
.Y(n_4806)
);

AND2x2_ASAP7_75t_L g4807 ( 
.A(n_4600),
.B(n_4293),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4577),
.Y(n_4808)
);

BUFx2_ASAP7_75t_L g4809 ( 
.A(n_4690),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_4532),
.Y(n_4810)
);

BUFx3_ASAP7_75t_L g4811 ( 
.A(n_4556),
.Y(n_4811)
);

BUFx10_ASAP7_75t_L g4812 ( 
.A(n_4605),
.Y(n_4812)
);

CKINVDCx5p33_ASAP7_75t_R g4813 ( 
.A(n_4558),
.Y(n_4813)
);

INVx2_ASAP7_75t_L g4814 ( 
.A(n_4586),
.Y(n_4814)
);

AOI22xp33_ASAP7_75t_L g4815 ( 
.A1(n_4563),
.A2(n_1694),
.B1(n_2030),
.B2(n_2412),
.Y(n_4815)
);

BUFx6f_ASAP7_75t_L g4816 ( 
.A(n_4675),
.Y(n_4816)
);

BUFx12f_ASAP7_75t_L g4817 ( 
.A(n_4641),
.Y(n_4817)
);

AOI22xp33_ASAP7_75t_L g4818 ( 
.A1(n_4637),
.A2(n_1694),
.B1(n_2433),
.B2(n_2412),
.Y(n_4818)
);

BUFx12f_ASAP7_75t_L g4819 ( 
.A(n_4551),
.Y(n_4819)
);

AOI22xp33_ASAP7_75t_L g4820 ( 
.A1(n_4731),
.A2(n_2443),
.B1(n_2433),
.B2(n_118),
.Y(n_4820)
);

AOI22xp33_ASAP7_75t_SL g4821 ( 
.A1(n_4668),
.A2(n_4301),
.B1(n_118),
.B2(n_114),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4585),
.Y(n_4822)
);

INVxp67_ASAP7_75t_SL g4823 ( 
.A(n_4550),
.Y(n_4823)
);

INVx4_ASAP7_75t_L g4824 ( 
.A(n_4576),
.Y(n_4824)
);

AOI22xp33_ASAP7_75t_L g4825 ( 
.A1(n_4638),
.A2(n_2443),
.B1(n_120),
.B2(n_116),
.Y(n_4825)
);

CKINVDCx5p33_ASAP7_75t_R g4826 ( 
.A(n_4605),
.Y(n_4826)
);

OAI22xp33_ASAP7_75t_L g4827 ( 
.A1(n_4727),
.A2(n_4757),
.B1(n_4599),
.B2(n_4647),
.Y(n_4827)
);

INVx3_ASAP7_75t_L g4828 ( 
.A(n_4691),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4591),
.Y(n_4829)
);

BUFx12f_ASAP7_75t_L g4830 ( 
.A(n_4575),
.Y(n_4830)
);

AND2x4_ASAP7_75t_SL g4831 ( 
.A(n_4719),
.B(n_2443),
.Y(n_4831)
);

AOI22xp33_ASAP7_75t_SL g4832 ( 
.A1(n_4672),
.A2(n_4301),
.B1(n_121),
.B2(n_119),
.Y(n_4832)
);

OAI22xp5_ASAP7_75t_L g4833 ( 
.A1(n_4666),
.A2(n_122),
.B1(n_119),
.B2(n_120),
.Y(n_4833)
);

HB1xp67_ASAP7_75t_L g4834 ( 
.A(n_4601),
.Y(n_4834)
);

AOI22xp33_ASAP7_75t_SL g4835 ( 
.A1(n_4576),
.A2(n_4647),
.B1(n_4687),
.B2(n_4545),
.Y(n_4835)
);

OAI22xp5_ASAP7_75t_L g4836 ( 
.A1(n_4593),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_4836)
);

INVx1_ASAP7_75t_L g4837 ( 
.A(n_4597),
.Y(n_4837)
);

OAI22xp33_ASAP7_75t_L g4838 ( 
.A1(n_4647),
.A2(n_4293),
.B1(n_126),
.B2(n_124),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4572),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4590),
.Y(n_4840)
);

BUFx12f_ASAP7_75t_L g4841 ( 
.A(n_4695),
.Y(n_4841)
);

AOI22xp33_ASAP7_75t_L g4842 ( 
.A1(n_4628),
.A2(n_2443),
.B1(n_127),
.B2(n_125),
.Y(n_4842)
);

BUFx6f_ASAP7_75t_L g4843 ( 
.A(n_4675),
.Y(n_4843)
);

AOI22xp33_ASAP7_75t_L g4844 ( 
.A1(n_4657),
.A2(n_129),
.B1(n_126),
.B2(n_127),
.Y(n_4844)
);

INVx3_ASAP7_75t_L g4845 ( 
.A(n_4550),
.Y(n_4845)
);

BUFx3_ASAP7_75t_L g4846 ( 
.A(n_4645),
.Y(n_4846)
);

BUFx3_ASAP7_75t_L g4847 ( 
.A(n_4676),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4528),
.Y(n_4848)
);

OAI22xp5_ASAP7_75t_SL g4849 ( 
.A1(n_4587),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4531),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_4617),
.Y(n_4851)
);

BUFx2_ASAP7_75t_SL g4852 ( 
.A(n_4722),
.Y(n_4852)
);

OAI22xp5_ASAP7_75t_L g4853 ( 
.A1(n_4744),
.A2(n_4667),
.B1(n_4655),
.B2(n_4705),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_4643),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4594),
.Y(n_4855)
);

BUFx3_ASAP7_75t_L g4856 ( 
.A(n_4659),
.Y(n_4856)
);

AOI22xp33_ASAP7_75t_L g4857 ( 
.A1(n_4658),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_4857)
);

AOI22xp33_ASAP7_75t_L g4858 ( 
.A1(n_4725),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4761),
.Y(n_4859)
);

INVx6_ASAP7_75t_L g4860 ( 
.A(n_4609),
.Y(n_4860)
);

INVx2_ASAP7_75t_L g4861 ( 
.A(n_4629),
.Y(n_4861)
);

AOI22xp33_ASAP7_75t_L g4862 ( 
.A1(n_4698),
.A2(n_138),
.B1(n_135),
.B2(n_136),
.Y(n_4862)
);

OAI22xp5_ASAP7_75t_L g4863 ( 
.A1(n_4741),
.A2(n_141),
.B1(n_138),
.B2(n_140),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4634),
.Y(n_4864)
);

INVx2_ASAP7_75t_L g4865 ( 
.A(n_4644),
.Y(n_4865)
);

AOI22xp33_ASAP7_75t_L g4866 ( 
.A1(n_4760),
.A2(n_4607),
.B1(n_4656),
.B2(n_4756),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4751),
.Y(n_4867)
);

AOI22xp33_ASAP7_75t_L g4868 ( 
.A1(n_4656),
.A2(n_144),
.B1(n_141),
.B2(n_142),
.Y(n_4868)
);

CKINVDCx8_ASAP7_75t_R g4869 ( 
.A(n_4609),
.Y(n_4869)
);

AOI22xp33_ASAP7_75t_SL g4870 ( 
.A1(n_4687),
.A2(n_145),
.B1(n_142),
.B2(n_144),
.Y(n_4870)
);

CKINVDCx20_ASAP7_75t_R g4871 ( 
.A(n_4716),
.Y(n_4871)
);

INVxp67_ASAP7_75t_SL g4872 ( 
.A(n_4763),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4701),
.Y(n_4873)
);

OAI21xp5_ASAP7_75t_L g4874 ( 
.A1(n_4729),
.A2(n_4293),
.B(n_145),
.Y(n_4874)
);

INVx2_ASAP7_75t_L g4875 ( 
.A(n_4648),
.Y(n_4875)
);

BUFx6f_ASAP7_75t_L g4876 ( 
.A(n_4675),
.Y(n_4876)
);

NAND2x1p5_ASAP7_75t_L g4877 ( 
.A(n_4736),
.B(n_1838),
.Y(n_4877)
);

BUFx3_ASAP7_75t_L g4878 ( 
.A(n_4609),
.Y(n_4878)
);

BUFx12f_ASAP7_75t_L g4879 ( 
.A(n_4723),
.Y(n_4879)
);

BUFx6f_ASAP7_75t_SL g4880 ( 
.A(n_4673),
.Y(n_4880)
);

CKINVDCx11_ASAP7_75t_R g4881 ( 
.A(n_4661),
.Y(n_4881)
);

INVx1_ASAP7_75t_L g4882 ( 
.A(n_4708),
.Y(n_4882)
);

AOI22xp33_ASAP7_75t_L g4883 ( 
.A1(n_4692),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_L g4884 ( 
.A(n_4539),
.B(n_4568),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4739),
.Y(n_4885)
);

CKINVDCx11_ASAP7_75t_R g4886 ( 
.A(n_4674),
.Y(n_4886)
);

INVx3_ASAP7_75t_L g4887 ( 
.A(n_4595),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4677),
.Y(n_4888)
);

CKINVDCx5p33_ASAP7_75t_R g4889 ( 
.A(n_4674),
.Y(n_4889)
);

AOI22xp33_ASAP7_75t_L g4890 ( 
.A1(n_4564),
.A2(n_150),
.B1(n_146),
.B2(n_148),
.Y(n_4890)
);

AOI22xp33_ASAP7_75t_SL g4891 ( 
.A1(n_4697),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_4891)
);

CKINVDCx5p33_ASAP7_75t_R g4892 ( 
.A(n_4674),
.Y(n_4892)
);

AOI22xp33_ASAP7_75t_L g4893 ( 
.A1(n_4673),
.A2(n_155),
.B1(n_152),
.B2(n_153),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4535),
.B(n_155),
.Y(n_4894)
);

INVx1_ASAP7_75t_L g4895 ( 
.A(n_4683),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4649),
.Y(n_4896)
);

AOI22xp33_ASAP7_75t_L g4897 ( 
.A1(n_4697),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_4897)
);

BUFx4f_ASAP7_75t_SL g4898 ( 
.A(n_4686),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4649),
.Y(n_4899)
);

AOI22xp33_ASAP7_75t_L g4900 ( 
.A1(n_4571),
.A2(n_4580),
.B1(n_4630),
.B2(n_4613),
.Y(n_4900)
);

INVx2_ASAP7_75t_L g4901 ( 
.A(n_4664),
.Y(n_4901)
);

INVx6_ASAP7_75t_L g4902 ( 
.A(n_4686),
.Y(n_4902)
);

INVx2_ASAP7_75t_L g4903 ( 
.A(n_4740),
.Y(n_4903)
);

INVx2_ASAP7_75t_L g4904 ( 
.A(n_4746),
.Y(n_4904)
);

BUFx4f_ASAP7_75t_SL g4905 ( 
.A(n_4686),
.Y(n_4905)
);

INVx3_ASAP7_75t_L g4906 ( 
.A(n_4595),
.Y(n_4906)
);

INVx1_ASAP7_75t_SL g4907 ( 
.A(n_4710),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4669),
.Y(n_4908)
);

INVx6_ASAP7_75t_L g4909 ( 
.A(n_4719),
.Y(n_4909)
);

AOI22xp33_ASAP7_75t_L g4910 ( 
.A1(n_4571),
.A2(n_164),
.B1(n_161),
.B2(n_163),
.Y(n_4910)
);

CKINVDCx11_ASAP7_75t_R g4911 ( 
.A(n_4621),
.Y(n_4911)
);

BUFx12f_ASAP7_75t_L g4912 ( 
.A(n_4720),
.Y(n_4912)
);

AND2x4_ASAP7_75t_L g4913 ( 
.A(n_4662),
.B(n_164),
.Y(n_4913)
);

BUFx12f_ASAP7_75t_L g4914 ( 
.A(n_4700),
.Y(n_4914)
);

NAND2xp5_ASAP7_75t_L g4915 ( 
.A(n_4540),
.B(n_165),
.Y(n_4915)
);

INVx2_ASAP7_75t_L g4916 ( 
.A(n_4752),
.Y(n_4916)
);

HB1xp67_ASAP7_75t_L g4917 ( 
.A(n_4711),
.Y(n_4917)
);

INVx4_ASAP7_75t_L g4918 ( 
.A(n_4631),
.Y(n_4918)
);

BUFx6f_ASAP7_75t_L g4919 ( 
.A(n_4631),
.Y(n_4919)
);

INVx2_ASAP7_75t_L g4920 ( 
.A(n_4730),
.Y(n_4920)
);

CKINVDCx20_ASAP7_75t_R g4921 ( 
.A(n_4714),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_4671),
.Y(n_4922)
);

CKINVDCx11_ASAP7_75t_R g4923 ( 
.A(n_4621),
.Y(n_4923)
);

AOI22xp33_ASAP7_75t_L g4924 ( 
.A1(n_4580),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_4924)
);

OAI22xp33_ASAP7_75t_L g4925 ( 
.A1(n_4770),
.A2(n_171),
.B1(n_168),
.B2(n_170),
.Y(n_4925)
);

OAI22xp33_ASAP7_75t_L g4926 ( 
.A1(n_4625),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4598),
.Y(n_4927)
);

INVx1_ASAP7_75t_L g4928 ( 
.A(n_4611),
.Y(n_4928)
);

BUFx10_ASAP7_75t_L g4929 ( 
.A(n_4560),
.Y(n_4929)
);

CKINVDCx11_ASAP7_75t_R g4930 ( 
.A(n_4555),
.Y(n_4930)
);

AOI22xp33_ASAP7_75t_L g4931 ( 
.A1(n_4632),
.A2(n_175),
.B1(n_172),
.B2(n_174),
.Y(n_4931)
);

OAI21xp5_ASAP7_75t_L g4932 ( 
.A1(n_4581),
.A2(n_174),
.B(n_175),
.Y(n_4932)
);

INVx6_ASAP7_75t_L g4933 ( 
.A(n_4533),
.Y(n_4933)
);

AOI22xp33_ASAP7_75t_L g4934 ( 
.A1(n_4574),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_4934)
);

INVx2_ASAP7_75t_L g4935 ( 
.A(n_4771),
.Y(n_4935)
);

CKINVDCx16_ASAP7_75t_R g4936 ( 
.A(n_4547),
.Y(n_4936)
);

AOI22xp33_ASAP7_75t_L g4937 ( 
.A1(n_4555),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_4937)
);

INVx2_ASAP7_75t_L g4938 ( 
.A(n_4768),
.Y(n_4938)
);

AOI22xp5_ASAP7_75t_L g4939 ( 
.A1(n_4639),
.A2(n_183),
.B1(n_180),
.B2(n_181),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4616),
.Y(n_4940)
);

INVx2_ASAP7_75t_L g4941 ( 
.A(n_4766),
.Y(n_4941)
);

OAI22xp5_ASAP7_75t_L g4942 ( 
.A1(n_4736),
.A2(n_184),
.B1(n_181),
.B2(n_183),
.Y(n_4942)
);

INVx2_ASAP7_75t_L g4943 ( 
.A(n_4754),
.Y(n_4943)
);

INVx1_ASAP7_75t_SL g4944 ( 
.A(n_4774),
.Y(n_4944)
);

AOI22xp33_ASAP7_75t_L g4945 ( 
.A1(n_4527),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4753),
.Y(n_4946)
);

CKINVDCx6p67_ASAP7_75t_R g4947 ( 
.A(n_4606),
.Y(n_4947)
);

AOI22xp5_ASAP7_75t_L g4948 ( 
.A1(n_4646),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_4948)
);

CKINVDCx5p33_ASAP7_75t_R g4949 ( 
.A(n_4608),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4682),
.Y(n_4950)
);

BUFx2_ASAP7_75t_SL g4951 ( 
.A(n_4694),
.Y(n_4951)
);

AOI22xp33_ASAP7_75t_L g4952 ( 
.A1(n_4635),
.A2(n_190),
.B1(n_187),
.B2(n_189),
.Y(n_4952)
);

BUFx12f_ASAP7_75t_L g4953 ( 
.A(n_4652),
.Y(n_4953)
);

OR2x2_ASAP7_75t_L g4954 ( 
.A(n_4743),
.B(n_189),
.Y(n_4954)
);

CKINVDCx20_ASAP7_75t_R g4955 ( 
.A(n_4718),
.Y(n_4955)
);

INVx8_ASAP7_75t_L g4956 ( 
.A(n_4560),
.Y(n_4956)
);

AOI22xp33_ASAP7_75t_L g4957 ( 
.A1(n_4541),
.A2(n_193),
.B1(n_190),
.B2(n_192),
.Y(n_4957)
);

OAI22xp5_ASAP7_75t_L g4958 ( 
.A1(n_4772),
.A2(n_4715),
.B1(n_4544),
.B2(n_4747),
.Y(n_4958)
);

AOI22xp33_ASAP7_75t_SL g4959 ( 
.A1(n_4592),
.A2(n_195),
.B1(n_192),
.B2(n_193),
.Y(n_4959)
);

AOI22xp33_ASAP7_75t_SL g4960 ( 
.A1(n_4640),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_4960)
);

AOI22xp5_ASAP7_75t_L g4961 ( 
.A1(n_4650),
.A2(n_199),
.B1(n_196),
.B2(n_198),
.Y(n_4961)
);

INVx2_ASAP7_75t_L g4962 ( 
.A(n_4769),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4584),
.Y(n_4963)
);

INVx2_ASAP7_75t_L g4964 ( 
.A(n_4769),
.Y(n_4964)
);

OAI22xp5_ASAP7_75t_L g4965 ( 
.A1(n_4713),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4589),
.Y(n_4966)
);

OAI22xp5_ASAP7_75t_L g4967 ( 
.A1(n_4792),
.A2(n_4702),
.B1(n_4703),
.B2(n_4670),
.Y(n_4967)
);

INVx3_ASAP7_75t_L g4968 ( 
.A(n_4828),
.Y(n_4968)
);

OR2x2_ASAP7_75t_L g4969 ( 
.A(n_4867),
.B(n_4684),
.Y(n_4969)
);

BUFx3_ASAP7_75t_L g4970 ( 
.A(n_4817),
.Y(n_4970)
);

NAND2xp5_ASAP7_75t_L g4971 ( 
.A(n_4805),
.B(n_4538),
.Y(n_4971)
);

OR2x2_ASAP7_75t_L g4972 ( 
.A(n_4851),
.B(n_4854),
.Y(n_4972)
);

AND2x6_ASAP7_75t_L g4973 ( 
.A(n_4913),
.B(n_4561),
.Y(n_4973)
);

CKINVDCx14_ASAP7_75t_R g4974 ( 
.A(n_4790),
.Y(n_4974)
);

AOI221xp5_ASAP7_75t_L g4975 ( 
.A1(n_4853),
.A2(n_4619),
.B1(n_4653),
.B2(n_4699),
.C(n_4663),
.Y(n_4975)
);

OA21x2_ASAP7_75t_L g4976 ( 
.A1(n_4896),
.A2(n_4615),
.B(n_4709),
.Y(n_4976)
);

AOI21xp5_ASAP7_75t_SL g4977 ( 
.A1(n_4932),
.A2(n_4561),
.B(n_4552),
.Y(n_4977)
);

AOI21xp5_ASAP7_75t_L g4978 ( 
.A1(n_4874),
.A2(n_4562),
.B(n_4688),
.Y(n_4978)
);

INVx2_ASAP7_75t_L g4979 ( 
.A(n_4859),
.Y(n_4979)
);

AND2x4_ASAP7_75t_L g4980 ( 
.A(n_4791),
.B(n_4665),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_L g4981 ( 
.A(n_4839),
.B(n_4567),
.Y(n_4981)
);

AND2x2_ASAP7_75t_L g4982 ( 
.A(n_4787),
.B(n_4702),
.Y(n_4982)
);

AND2x2_ASAP7_75t_L g4983 ( 
.A(n_4779),
.B(n_4703),
.Y(n_4983)
);

BUFx2_ASAP7_75t_L g4984 ( 
.A(n_4828),
.Y(n_4984)
);

AND2x4_ASAP7_75t_L g4985 ( 
.A(n_4791),
.B(n_4680),
.Y(n_4985)
);

INVx2_ASAP7_75t_L g4986 ( 
.A(n_4777),
.Y(n_4986)
);

AOI22xp33_ASAP7_75t_L g4987 ( 
.A1(n_4833),
.A2(n_4773),
.B1(n_4624),
.B2(n_4636),
.Y(n_4987)
);

AOI21xp5_ASAP7_75t_SL g4988 ( 
.A1(n_4800),
.A2(n_4773),
.B(n_4537),
.Y(n_4988)
);

AND2x2_ASAP7_75t_L g4989 ( 
.A(n_4793),
.B(n_4685),
.Y(n_4989)
);

AND2x2_ASAP7_75t_L g4990 ( 
.A(n_4793),
.B(n_4749),
.Y(n_4990)
);

NAND2xp5_ASAP7_75t_L g4991 ( 
.A(n_4946),
.B(n_4755),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4899),
.Y(n_4992)
);

AND2x2_ASAP7_75t_L g4993 ( 
.A(n_4809),
.B(n_4749),
.Y(n_4993)
);

OR2x2_ASAP7_75t_L g4994 ( 
.A(n_4807),
.B(n_4689),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4781),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4789),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4944),
.B(n_4603),
.Y(n_4997)
);

NAND2x1_ASAP7_75t_L g4998 ( 
.A(n_4824),
.B(n_4623),
.Y(n_4998)
);

NAND2xp5_ASAP7_75t_L g4999 ( 
.A(n_4944),
.B(n_4570),
.Y(n_4999)
);

AND2x2_ASAP7_75t_L g5000 ( 
.A(n_4801),
.B(n_4726),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_4834),
.B(n_4536),
.Y(n_5001)
);

INVx1_ASAP7_75t_SL g5002 ( 
.A(n_4881),
.Y(n_5002)
);

AND2x4_ASAP7_75t_L g5003 ( 
.A(n_4791),
.B(n_4887),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_4801),
.B(n_4726),
.Y(n_5004)
);

INVx1_ASAP7_75t_L g5005 ( 
.A(n_4795),
.Y(n_5005)
);

AND2x2_ASAP7_75t_L g5006 ( 
.A(n_4856),
.B(n_4726),
.Y(n_5006)
);

AND2x4_ASAP7_75t_L g5007 ( 
.A(n_4887),
.B(n_4724),
.Y(n_5007)
);

NOR2xp67_ASAP7_75t_L g5008 ( 
.A(n_4798),
.B(n_4733),
.Y(n_5008)
);

HB1xp67_ASAP7_75t_L g5009 ( 
.A(n_4917),
.Y(n_5009)
);

OAI22xp5_ASAP7_75t_L g5010 ( 
.A1(n_4939),
.A2(n_4573),
.B1(n_4660),
.B2(n_4767),
.Y(n_5010)
);

CKINVDCx16_ASAP7_75t_R g5011 ( 
.A(n_4871),
.Y(n_5011)
);

INVx1_ASAP7_75t_L g5012 ( 
.A(n_4799),
.Y(n_5012)
);

O2A1O1Ixp5_ASAP7_75t_L g5013 ( 
.A1(n_4827),
.A2(n_4838),
.B(n_4780),
.C(n_4950),
.Y(n_5013)
);

OR2x6_ASAP7_75t_L g5014 ( 
.A(n_4956),
.B(n_4745),
.Y(n_5014)
);

NOR2xp33_ASAP7_75t_SL g5015 ( 
.A(n_4798),
.B(n_4636),
.Y(n_5015)
);

O2A1O1Ixp33_ASAP7_75t_L g5016 ( 
.A1(n_4925),
.A2(n_4737),
.B(n_4707),
.C(n_4610),
.Y(n_5016)
);

BUFx2_ASAP7_75t_L g5017 ( 
.A(n_4918),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_4808),
.Y(n_5018)
);

AND2x4_ASAP7_75t_L g5019 ( 
.A(n_4906),
.B(n_4758),
.Y(n_5019)
);

A2O1A1Ixp33_ASAP7_75t_SL g5020 ( 
.A1(n_4815),
.A2(n_4534),
.B(n_4651),
.C(n_4622),
.Y(n_5020)
);

INVx2_ASAP7_75t_L g5021 ( 
.A(n_4803),
.Y(n_5021)
);

BUFx4f_ASAP7_75t_L g5022 ( 
.A(n_4841),
.Y(n_5022)
);

AOI21xp5_ASAP7_75t_SL g5023 ( 
.A1(n_4824),
.A2(n_4679),
.B(n_4578),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4822),
.Y(n_5024)
);

NAND2xp5_ASAP7_75t_L g5025 ( 
.A(n_4855),
.B(n_4582),
.Y(n_5025)
);

AOI21x1_ASAP7_75t_SL g5026 ( 
.A1(n_4913),
.A2(n_4894),
.B(n_4884),
.Y(n_5026)
);

OR2x2_ASAP7_75t_L g5027 ( 
.A(n_4927),
.B(n_4681),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_4810),
.Y(n_5028)
);

AND2x2_ASAP7_75t_L g5029 ( 
.A(n_4909),
.B(n_4775),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_L g5030 ( 
.A(n_4963),
.B(n_4565),
.Y(n_5030)
);

AND2x2_ASAP7_75t_L g5031 ( 
.A(n_4909),
.B(n_4775),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_4966),
.B(n_4762),
.Y(n_5032)
);

O2A1O1Ixp33_ASAP7_75t_L g5033 ( 
.A1(n_4926),
.A2(n_4654),
.B(n_4604),
.C(n_4706),
.Y(n_5033)
);

AOI211xp5_ASAP7_75t_L g5034 ( 
.A1(n_4849),
.A2(n_4732),
.B(n_4717),
.C(n_4627),
.Y(n_5034)
);

AOI21x1_ASAP7_75t_SL g5035 ( 
.A1(n_4915),
.A2(n_4579),
.B(n_4712),
.Y(n_5035)
);

BUFx12f_ASAP7_75t_L g5036 ( 
.A(n_4813),
.Y(n_5036)
);

AOI21x1_ASAP7_75t_SL g5037 ( 
.A1(n_4911),
.A2(n_4579),
.B(n_4712),
.Y(n_5037)
);

AOI21x1_ASAP7_75t_SL g5038 ( 
.A1(n_4923),
.A2(n_4579),
.B(n_4712),
.Y(n_5038)
);

AOI21xp5_ASAP7_75t_SL g5039 ( 
.A1(n_4880),
.A2(n_4764),
.B(n_4759),
.Y(n_5039)
);

HB1xp67_ASAP7_75t_L g5040 ( 
.A(n_4907),
.Y(n_5040)
);

AND2x2_ASAP7_75t_L g5041 ( 
.A(n_4823),
.B(n_4733),
.Y(n_5041)
);

AND2x4_ASAP7_75t_L g5042 ( 
.A(n_4906),
.B(n_4733),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_4848),
.B(n_4704),
.Y(n_5043)
);

OAI22xp5_ASAP7_75t_L g5044 ( 
.A1(n_4939),
.A2(n_4557),
.B1(n_4693),
.B2(n_4750),
.Y(n_5044)
);

NOR2xp67_ASAP7_75t_L g5045 ( 
.A(n_4826),
.B(n_4918),
.Y(n_5045)
);

AOI21xp5_ASAP7_75t_SL g5046 ( 
.A1(n_4880),
.A2(n_4623),
.B(n_4765),
.Y(n_5046)
);

AND2x2_ASAP7_75t_L g5047 ( 
.A(n_4847),
.B(n_4623),
.Y(n_5047)
);

AND2x4_ASAP7_75t_L g5048 ( 
.A(n_4845),
.B(n_4623),
.Y(n_5048)
);

AND2x4_ASAP7_75t_L g5049 ( 
.A(n_4845),
.B(n_201),
.Y(n_5049)
);

AND2x2_ASAP7_75t_L g5050 ( 
.A(n_4951),
.B(n_202),
.Y(n_5050)
);

AND2x2_ASAP7_75t_L g5051 ( 
.A(n_4875),
.B(n_206),
.Y(n_5051)
);

O2A1O1Ixp33_ASAP7_75t_L g5052 ( 
.A1(n_4965),
.A2(n_209),
.B(n_207),
.C(n_208),
.Y(n_5052)
);

INVx5_ASAP7_75t_L g5053 ( 
.A(n_4812),
.Y(n_5053)
);

AND2x2_ASAP7_75t_L g5054 ( 
.A(n_4901),
.B(n_207),
.Y(n_5054)
);

INVx2_ASAP7_75t_L g5055 ( 
.A(n_4814),
.Y(n_5055)
);

O2A1O1Ixp33_ASAP7_75t_L g5056 ( 
.A1(n_4942),
.A2(n_210),
.B(n_208),
.C(n_209),
.Y(n_5056)
);

OAI22xp5_ASAP7_75t_L g5057 ( 
.A1(n_4900),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_5057)
);

AND2x2_ASAP7_75t_L g5058 ( 
.A(n_4861),
.B(n_211),
.Y(n_5058)
);

O2A1O1Ixp33_ASAP7_75t_L g5059 ( 
.A1(n_4863),
.A2(n_214),
.B(n_212),
.C(n_213),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_4829),
.Y(n_5060)
);

O2A1O1Ixp5_ASAP7_75t_L g5061 ( 
.A1(n_4784),
.A2(n_216),
.B(n_213),
.C(n_215),
.Y(n_5061)
);

AOI21x1_ASAP7_75t_SL g5062 ( 
.A1(n_4835),
.A2(n_215),
.B(n_218),
.Y(n_5062)
);

INVx1_ASAP7_75t_L g5063 ( 
.A(n_4837),
.Y(n_5063)
);

AOI21x1_ASAP7_75t_SL g5064 ( 
.A1(n_4849),
.A2(n_220),
.B(n_221),
.Y(n_5064)
);

NOR2xp67_ASAP7_75t_L g5065 ( 
.A(n_4962),
.B(n_220),
.Y(n_5065)
);

AOI21xp5_ASAP7_75t_L g5066 ( 
.A1(n_4960),
.A2(n_1849),
.B(n_1838),
.Y(n_5066)
);

NOR2xp67_ASAP7_75t_L g5067 ( 
.A(n_4964),
.B(n_221),
.Y(n_5067)
);

NAND2xp5_ASAP7_75t_L g5068 ( 
.A(n_4850),
.B(n_222),
.Y(n_5068)
);

AND2x2_ASAP7_75t_L g5069 ( 
.A(n_4936),
.B(n_222),
.Y(n_5069)
);

AND2x2_ASAP7_75t_L g5070 ( 
.A(n_4852),
.B(n_223),
.Y(n_5070)
);

AOI21xp5_ASAP7_75t_L g5071 ( 
.A1(n_4821),
.A2(n_1849),
.B(n_1838),
.Y(n_5071)
);

HB1xp67_ASAP7_75t_L g5072 ( 
.A(n_4907),
.Y(n_5072)
);

HB1xp67_ASAP7_75t_L g5073 ( 
.A(n_4920),
.Y(n_5073)
);

OR2x2_ASAP7_75t_L g5074 ( 
.A(n_4928),
.B(n_223),
.Y(n_5074)
);

AND2x2_ASAP7_75t_L g5075 ( 
.A(n_4840),
.B(n_224),
.Y(n_5075)
);

HB1xp67_ASAP7_75t_L g5076 ( 
.A(n_4943),
.Y(n_5076)
);

AND2x2_ASAP7_75t_L g5077 ( 
.A(n_4864),
.B(n_224),
.Y(n_5077)
);

AND2x2_ASAP7_75t_L g5078 ( 
.A(n_4947),
.B(n_226),
.Y(n_5078)
);

BUFx2_ASAP7_75t_L g5079 ( 
.A(n_4919),
.Y(n_5079)
);

OAI22xp5_ASAP7_75t_L g5080 ( 
.A1(n_4959),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.Y(n_5080)
);

AOI211xp5_ASAP7_75t_L g5081 ( 
.A1(n_4948),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_5081)
);

O2A1O1Ixp33_ASAP7_75t_L g5082 ( 
.A1(n_4958),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_5082)
);

O2A1O1Ixp5_ASAP7_75t_L g5083 ( 
.A1(n_4940),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_5083)
);

AND2x4_ASAP7_75t_L g5084 ( 
.A(n_4941),
.B(n_234),
.Y(n_5084)
);

O2A1O1Ixp33_ASAP7_75t_L g5085 ( 
.A1(n_4836),
.A2(n_238),
.B(n_235),
.C(n_236),
.Y(n_5085)
);

AOI21xp5_ASAP7_75t_L g5086 ( 
.A1(n_4832),
.A2(n_1849),
.B(n_1838),
.Y(n_5086)
);

INVx3_ASAP7_75t_L g5087 ( 
.A(n_4919),
.Y(n_5087)
);

OAI211xp5_ASAP7_75t_L g5088 ( 
.A1(n_4948),
.A2(n_241),
.B(n_238),
.C(n_239),
.Y(n_5088)
);

NAND2xp5_ASAP7_75t_L g5089 ( 
.A(n_4865),
.B(n_239),
.Y(n_5089)
);

OR2x2_ASAP7_75t_L g5090 ( 
.A(n_4797),
.B(n_4872),
.Y(n_5090)
);

AND2x2_ASAP7_75t_L g5091 ( 
.A(n_4846),
.B(n_243),
.Y(n_5091)
);

OR2x2_ASAP7_75t_L g5092 ( 
.A(n_4873),
.B(n_243),
.Y(n_5092)
);

NAND2xp5_ASAP7_75t_L g5093 ( 
.A(n_4866),
.B(n_244),
.Y(n_5093)
);

OAI22xp5_ASAP7_75t_L g5094 ( 
.A1(n_4931),
.A2(n_248),
.B1(n_244),
.B2(n_246),
.Y(n_5094)
);

BUFx12f_ASAP7_75t_L g5095 ( 
.A(n_4812),
.Y(n_5095)
);

O2A1O1Ixp33_ASAP7_75t_L g5096 ( 
.A1(n_4844),
.A2(n_249),
.B(n_246),
.C(n_248),
.Y(n_5096)
);

BUFx2_ASAP7_75t_L g5097 ( 
.A(n_4919),
.Y(n_5097)
);

CKINVDCx20_ASAP7_75t_R g5098 ( 
.A(n_4785),
.Y(n_5098)
);

HB1xp67_ASAP7_75t_L g5099 ( 
.A(n_4882),
.Y(n_5099)
);

AOI21xp5_ASAP7_75t_SL g5100 ( 
.A1(n_4778),
.A2(n_249),
.B(n_250),
.Y(n_5100)
);

BUFx6f_ASAP7_75t_L g5101 ( 
.A(n_4886),
.Y(n_5101)
);

AOI21xp5_ASAP7_75t_SL g5102 ( 
.A1(n_4877),
.A2(n_251),
.B(n_256),
.Y(n_5102)
);

OAI22xp5_ASAP7_75t_SL g5103 ( 
.A1(n_4921),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_5103)
);

OAI22xp5_ASAP7_75t_L g5104 ( 
.A1(n_4961),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_5104)
);

OA21x2_ASAP7_75t_L g5105 ( 
.A1(n_4885),
.A2(n_260),
.B(n_261),
.Y(n_5105)
);

OAI22xp5_ASAP7_75t_L g5106 ( 
.A1(n_4961),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_5106)
);

AOI21x1_ASAP7_75t_SL g5107 ( 
.A1(n_4796),
.A2(n_262),
.B(n_263),
.Y(n_5107)
);

AND2x2_ASAP7_75t_L g5108 ( 
.A(n_4776),
.B(n_264),
.Y(n_5108)
);

AOI21xp5_ASAP7_75t_SL g5109 ( 
.A1(n_4811),
.A2(n_265),
.B(n_266),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_4888),
.Y(n_5110)
);

NAND2xp5_ASAP7_75t_L g5111 ( 
.A(n_4895),
.B(n_265),
.Y(n_5111)
);

OA21x2_ASAP7_75t_L g5112 ( 
.A1(n_4908),
.A2(n_267),
.B(n_268),
.Y(n_5112)
);

HB1xp67_ASAP7_75t_L g5113 ( 
.A(n_4922),
.Y(n_5113)
);

OAI22xp5_ASAP7_75t_L g5114 ( 
.A1(n_4870),
.A2(n_272),
.B1(n_269),
.B2(n_271),
.Y(n_5114)
);

INVx2_ASAP7_75t_L g5115 ( 
.A(n_4972),
.Y(n_5115)
);

NAND2x1p5_ASAP7_75t_L g5116 ( 
.A(n_4980),
.B(n_4878),
.Y(n_5116)
);

AO31x2_ASAP7_75t_L g5117 ( 
.A1(n_4978),
.A2(n_4935),
.A3(n_4904),
.B(n_4916),
.Y(n_5117)
);

AND2x2_ASAP7_75t_L g5118 ( 
.A(n_5029),
.B(n_4933),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_5110),
.Y(n_5119)
);

AND2x2_ASAP7_75t_L g5120 ( 
.A(n_5031),
.B(n_4933),
.Y(n_5120)
);

AO31x2_ASAP7_75t_L g5121 ( 
.A1(n_4992),
.A2(n_4903),
.A3(n_4938),
.B(n_4869),
.Y(n_5121)
);

OR2x6_ASAP7_75t_L g5122 ( 
.A(n_5039),
.B(n_4956),
.Y(n_5122)
);

CKINVDCx16_ASAP7_75t_R g5123 ( 
.A(n_4974),
.Y(n_5123)
);

INVx2_ASAP7_75t_L g5124 ( 
.A(n_4990),
.Y(n_5124)
);

BUFx12f_ASAP7_75t_L g5125 ( 
.A(n_5101),
.Y(n_5125)
);

HB1xp67_ASAP7_75t_L g5126 ( 
.A(n_5040),
.Y(n_5126)
);

AOI22xp33_ASAP7_75t_SL g5127 ( 
.A1(n_5088),
.A2(n_4914),
.B1(n_4912),
.B2(n_4879),
.Y(n_5127)
);

AND2x4_ASAP7_75t_L g5128 ( 
.A(n_5045),
.B(n_4816),
.Y(n_5128)
);

AOI22xp33_ASAP7_75t_SL g5129 ( 
.A1(n_5104),
.A2(n_4956),
.B1(n_4953),
.B2(n_4955),
.Y(n_5129)
);

CKINVDCx16_ASAP7_75t_R g5130 ( 
.A(n_5011),
.Y(n_5130)
);

AND2x2_ASAP7_75t_L g5131 ( 
.A(n_5000),
.B(n_5004),
.Y(n_5131)
);

INVx2_ASAP7_75t_L g5132 ( 
.A(n_4993),
.Y(n_5132)
);

OR2x2_ASAP7_75t_L g5133 ( 
.A(n_4969),
.B(n_4954),
.Y(n_5133)
);

OAI22xp5_ASAP7_75t_L g5134 ( 
.A1(n_5081),
.A2(n_4897),
.B1(n_4891),
.B2(n_4893),
.Y(n_5134)
);

BUFx10_ASAP7_75t_L g5135 ( 
.A(n_5101),
.Y(n_5135)
);

OR2x2_ASAP7_75t_L g5136 ( 
.A(n_4991),
.B(n_4782),
.Y(n_5136)
);

OR2x2_ASAP7_75t_L g5137 ( 
.A(n_5001),
.B(n_4782),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_5110),
.Y(n_5138)
);

OAI22xp5_ASAP7_75t_L g5139 ( 
.A1(n_4977),
.A2(n_4868),
.B1(n_4825),
.B2(n_4910),
.Y(n_5139)
);

INVx2_ASAP7_75t_L g5140 ( 
.A(n_5041),
.Y(n_5140)
);

NAND2xp5_ASAP7_75t_L g5141 ( 
.A(n_5030),
.B(n_4997),
.Y(n_5141)
);

AOI21xp5_ASAP7_75t_L g5142 ( 
.A1(n_5100),
.A2(n_4857),
.B(n_4788),
.Y(n_5142)
);

HB1xp67_ASAP7_75t_L g5143 ( 
.A(n_5072),
.Y(n_5143)
);

BUFx2_ASAP7_75t_L g5144 ( 
.A(n_4984),
.Y(n_5144)
);

AND2x2_ASAP7_75t_L g5145 ( 
.A(n_5006),
.B(n_4949),
.Y(n_5145)
);

OAI21xp5_ASAP7_75t_L g5146 ( 
.A1(n_5013),
.A2(n_4952),
.B(n_4934),
.Y(n_5146)
);

OAI22xp5_ASAP7_75t_L g5147 ( 
.A1(n_4988),
.A2(n_4924),
.B1(n_4820),
.B2(n_4937),
.Y(n_5147)
);

NOR2xp33_ASAP7_75t_R g5148 ( 
.A(n_5101),
.B(n_4796),
.Y(n_5148)
);

AND2x2_ASAP7_75t_L g5149 ( 
.A(n_4982),
.B(n_4889),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_5099),
.Y(n_5150)
);

INVx2_ASAP7_75t_L g5151 ( 
.A(n_5090),
.Y(n_5151)
);

CKINVDCx5p33_ASAP7_75t_R g5152 ( 
.A(n_5098),
.Y(n_5152)
);

NOR3xp33_ASAP7_75t_SL g5153 ( 
.A(n_5103),
.B(n_4892),
.C(n_4796),
.Y(n_5153)
);

HB1xp67_ASAP7_75t_L g5154 ( 
.A(n_5009),
.Y(n_5154)
);

BUFx12f_ASAP7_75t_L g5155 ( 
.A(n_5095),
.Y(n_5155)
);

OAI22xp5_ASAP7_75t_L g5156 ( 
.A1(n_4987),
.A2(n_4842),
.B1(n_4818),
.B2(n_4862),
.Y(n_5156)
);

AOI22xp5_ASAP7_75t_L g5157 ( 
.A1(n_5106),
.A2(n_4930),
.B1(n_4883),
.B2(n_4858),
.Y(n_5157)
);

BUFx2_ASAP7_75t_L g5158 ( 
.A(n_4980),
.Y(n_5158)
);

INVxp67_ASAP7_75t_L g5159 ( 
.A(n_4971),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_5113),
.Y(n_5160)
);

AOI22xp33_ASAP7_75t_L g5161 ( 
.A1(n_5114),
.A2(n_4957),
.B1(n_4890),
.B2(n_4794),
.Y(n_5161)
);

CKINVDCx16_ASAP7_75t_R g5162 ( 
.A(n_5036),
.Y(n_5162)
);

AND2x2_ASAP7_75t_L g5163 ( 
.A(n_4983),
.B(n_4786),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_4992),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_4995),
.Y(n_5165)
);

HB1xp67_ASAP7_75t_L g5166 ( 
.A(n_5076),
.Y(n_5166)
);

BUFx6f_ASAP7_75t_L g5167 ( 
.A(n_5053),
.Y(n_5167)
);

AND2x2_ASAP7_75t_L g5168 ( 
.A(n_5079),
.B(n_4786),
.Y(n_5168)
);

OR2x6_ASAP7_75t_L g5169 ( 
.A(n_5046),
.B(n_4819),
.Y(n_5169)
);

AND2x2_ASAP7_75t_L g5170 ( 
.A(n_5097),
.B(n_4830),
.Y(n_5170)
);

INVx1_ASAP7_75t_L g5171 ( 
.A(n_4996),
.Y(n_5171)
);

HB1xp67_ASAP7_75t_L g5172 ( 
.A(n_4994),
.Y(n_5172)
);

INVx2_ASAP7_75t_L g5173 ( 
.A(n_5017),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_5005),
.Y(n_5174)
);

BUFx6f_ASAP7_75t_L g5175 ( 
.A(n_5053),
.Y(n_5175)
);

NAND2xp33_ASAP7_75t_R g5176 ( 
.A(n_5069),
.B(n_5078),
.Y(n_5176)
);

BUFx12f_ASAP7_75t_L g5177 ( 
.A(n_5108),
.Y(n_5177)
);

INVx1_ASAP7_75t_L g5178 ( 
.A(n_5012),
.Y(n_5178)
);

INVx2_ASAP7_75t_L g5179 ( 
.A(n_4979),
.Y(n_5179)
);

HB1xp67_ASAP7_75t_L g5180 ( 
.A(n_5027),
.Y(n_5180)
);

INVx11_ASAP7_75t_L g5181 ( 
.A(n_4973),
.Y(n_5181)
);

INVx2_ASAP7_75t_L g5182 ( 
.A(n_5003),
.Y(n_5182)
);

AO31x2_ASAP7_75t_L g5183 ( 
.A1(n_5032),
.A2(n_4902),
.A3(n_4860),
.B(n_4898),
.Y(n_5183)
);

INVx1_ASAP7_75t_L g5184 ( 
.A(n_5018),
.Y(n_5184)
);

OAI21x1_ASAP7_75t_L g5185 ( 
.A1(n_5025),
.A2(n_4783),
.B(n_4804),
.Y(n_5185)
);

NAND2xp5_ASAP7_75t_L g5186 ( 
.A(n_4999),
.B(n_4816),
.Y(n_5186)
);

CKINVDCx16_ASAP7_75t_R g5187 ( 
.A(n_5015),
.Y(n_5187)
);

AND2x2_ASAP7_75t_L g5188 ( 
.A(n_4989),
.B(n_4929),
.Y(n_5188)
);

HB1xp67_ASAP7_75t_L g5189 ( 
.A(n_5073),
.Y(n_5189)
);

AND2x2_ASAP7_75t_L g5190 ( 
.A(n_5003),
.B(n_4985),
.Y(n_5190)
);

O2A1O1Ixp5_ASAP7_75t_L g5191 ( 
.A1(n_5061),
.A2(n_4929),
.B(n_4905),
.C(n_4902),
.Y(n_5191)
);

NOR2xp33_ASAP7_75t_R g5192 ( 
.A(n_5022),
.B(n_4860),
.Y(n_5192)
);

NOR2xp33_ASAP7_75t_L g5193 ( 
.A(n_5053),
.B(n_4816),
.Y(n_5193)
);

AOI22xp33_ASAP7_75t_L g5194 ( 
.A1(n_5071),
.A2(n_4945),
.B1(n_4802),
.B2(n_4806),
.Y(n_5194)
);

INVx1_ASAP7_75t_SL g5195 ( 
.A(n_5002),
.Y(n_5195)
);

INVx2_ASAP7_75t_L g5196 ( 
.A(n_5021),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_5024),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_5028),
.Y(n_5198)
);

INVx3_ASAP7_75t_L g5199 ( 
.A(n_4985),
.Y(n_5199)
);

OR2x2_ASAP7_75t_L g5200 ( 
.A(n_4986),
.B(n_4843),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_5060),
.Y(n_5201)
);

INVx2_ASAP7_75t_L g5202 ( 
.A(n_4968),
.Y(n_5202)
);

OR2x6_ASAP7_75t_L g5203 ( 
.A(n_5008),
.B(n_5023),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_5063),
.Y(n_5204)
);

INVx2_ASAP7_75t_L g5205 ( 
.A(n_4968),
.Y(n_5205)
);

BUFx3_ASAP7_75t_L g5206 ( 
.A(n_4970),
.Y(n_5206)
);

CKINVDCx5p33_ASAP7_75t_R g5207 ( 
.A(n_5022),
.Y(n_5207)
);

OR2x2_ASAP7_75t_L g5208 ( 
.A(n_5055),
.B(n_4843),
.Y(n_5208)
);

INVx8_ASAP7_75t_L g5209 ( 
.A(n_5050),
.Y(n_5209)
);

AND2x4_ASAP7_75t_L g5210 ( 
.A(n_5014),
.B(n_4876),
.Y(n_5210)
);

INVx3_ASAP7_75t_L g5211 ( 
.A(n_5042),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_5111),
.Y(n_5212)
);

NOR2xp33_ASAP7_75t_R g5213 ( 
.A(n_5070),
.B(n_272),
.Y(n_5213)
);

CKINVDCx16_ASAP7_75t_R g5214 ( 
.A(n_4973),
.Y(n_5214)
);

OR2x2_ASAP7_75t_L g5215 ( 
.A(n_4981),
.B(n_4843),
.Y(n_5215)
);

AOI22xp33_ASAP7_75t_L g5216 ( 
.A1(n_5086),
.A2(n_4831),
.B1(n_4876),
.B2(n_1849),
.Y(n_5216)
);

AND2x2_ASAP7_75t_L g5217 ( 
.A(n_5019),
.B(n_4876),
.Y(n_5217)
);

NAND2xp5_ASAP7_75t_L g5218 ( 
.A(n_5043),
.B(n_273),
.Y(n_5218)
);

CKINVDCx16_ASAP7_75t_R g5219 ( 
.A(n_4973),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_5092),
.Y(n_5220)
);

NAND3xp33_ASAP7_75t_SL g5221 ( 
.A(n_5082),
.B(n_5093),
.C(n_5034),
.Y(n_5221)
);

AND2x2_ASAP7_75t_L g5222 ( 
.A(n_5019),
.B(n_274),
.Y(n_5222)
);

NOR2xp33_ASAP7_75t_R g5223 ( 
.A(n_4973),
.B(n_274),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_L g5224 ( 
.A(n_5007),
.B(n_275),
.Y(n_5224)
);

AND2x4_ASAP7_75t_L g5225 ( 
.A(n_5014),
.B(n_275),
.Y(n_5225)
);

NAND2xp5_ASAP7_75t_L g5226 ( 
.A(n_5007),
.B(n_276),
.Y(n_5226)
);

AOI22xp33_ASAP7_75t_SL g5227 ( 
.A1(n_5057),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_5074),
.Y(n_5228)
);

NAND2xp33_ASAP7_75t_L g5229 ( 
.A(n_5080),
.B(n_279),
.Y(n_5229)
);

AOI22xp33_ASAP7_75t_SL g5230 ( 
.A1(n_5094),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_5230)
);

NOR3xp33_ASAP7_75t_SL g5231 ( 
.A(n_4975),
.B(n_281),
.C(n_282),
.Y(n_5231)
);

OAI22xp33_ASAP7_75t_L g5232 ( 
.A1(n_4967),
.A2(n_5044),
.B1(n_5010),
.B2(n_5105),
.Y(n_5232)
);

CKINVDCx5p33_ASAP7_75t_R g5233 ( 
.A(n_5087),
.Y(n_5233)
);

NAND3xp33_ASAP7_75t_SL g5234 ( 
.A(n_5016),
.B(n_284),
.C(n_285),
.Y(n_5234)
);

AOI22xp33_ASAP7_75t_L g5235 ( 
.A1(n_5066),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_5235)
);

AOI22xp33_ASAP7_75t_L g5236 ( 
.A1(n_5105),
.A2(n_291),
.B1(n_288),
.B2(n_289),
.Y(n_5236)
);

INVx2_ASAP7_75t_L g5237 ( 
.A(n_5087),
.Y(n_5237)
);

INVx2_ASAP7_75t_L g5238 ( 
.A(n_5042),
.Y(n_5238)
);

BUFx6f_ASAP7_75t_L g5239 ( 
.A(n_5084),
.Y(n_5239)
);

CKINVDCx11_ASAP7_75t_R g5240 ( 
.A(n_5049),
.Y(n_5240)
);

INVx2_ASAP7_75t_L g5241 ( 
.A(n_5084),
.Y(n_5241)
);

AO32x2_ASAP7_75t_L g5242 ( 
.A1(n_5035),
.A2(n_292),
.A3(n_289),
.B1(n_291),
.B2(n_293),
.Y(n_5242)
);

XNOR2xp5_ASAP7_75t_L g5243 ( 
.A(n_5091),
.B(n_295),
.Y(n_5243)
);

INVx2_ASAP7_75t_L g5244 ( 
.A(n_5077),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_5112),
.Y(n_5245)
);

OAI22xp5_ASAP7_75t_L g5246 ( 
.A1(n_5109),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_5246)
);

OR2x2_ASAP7_75t_L g5247 ( 
.A(n_5068),
.B(n_297),
.Y(n_5247)
);

NAND2xp33_ASAP7_75t_R g5248 ( 
.A(n_5049),
.B(n_298),
.Y(n_5248)
);

BUFx2_ASAP7_75t_L g5249 ( 
.A(n_5048),
.Y(n_5249)
);

INVx2_ASAP7_75t_SL g5250 ( 
.A(n_5047),
.Y(n_5250)
);

INVx1_ASAP7_75t_L g5251 ( 
.A(n_5112),
.Y(n_5251)
);

AND2x4_ASAP7_75t_L g5252 ( 
.A(n_5048),
.B(n_298),
.Y(n_5252)
);

AND2x4_ASAP7_75t_L g5253 ( 
.A(n_4998),
.B(n_299),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_5089),
.Y(n_5254)
);

BUFx6f_ASAP7_75t_L g5255 ( 
.A(n_5051),
.Y(n_5255)
);

OAI21xp5_ASAP7_75t_L g5256 ( 
.A1(n_5083),
.A2(n_5052),
.B(n_5065),
.Y(n_5256)
);

INVx2_ASAP7_75t_L g5257 ( 
.A(n_5058),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_5119),
.Y(n_5258)
);

INVx4_ASAP7_75t_L g5259 ( 
.A(n_5125),
.Y(n_5259)
);

INVx2_ASAP7_75t_L g5260 ( 
.A(n_5158),
.Y(n_5260)
);

INVx2_ASAP7_75t_L g5261 ( 
.A(n_5237),
.Y(n_5261)
);

OR2x6_ASAP7_75t_L g5262 ( 
.A(n_5169),
.B(n_5102),
.Y(n_5262)
);

AOI21x1_ASAP7_75t_L g5263 ( 
.A1(n_5169),
.A2(n_5203),
.B(n_5122),
.Y(n_5263)
);

AO21x2_ASAP7_75t_L g5264 ( 
.A1(n_5245),
.A2(n_5075),
.B(n_5054),
.Y(n_5264)
);

AO21x2_ASAP7_75t_L g5265 ( 
.A1(n_5251),
.A2(n_5067),
.B(n_5056),
.Y(n_5265)
);

INVx3_ASAP7_75t_L g5266 ( 
.A(n_5167),
.Y(n_5266)
);

AOI211xp5_ASAP7_75t_L g5267 ( 
.A1(n_5234),
.A2(n_5096),
.B(n_5059),
.C(n_5085),
.Y(n_5267)
);

INVx1_ASAP7_75t_L g5268 ( 
.A(n_5138),
.Y(n_5268)
);

BUFx3_ASAP7_75t_L g5269 ( 
.A(n_5135),
.Y(n_5269)
);

AO21x2_ASAP7_75t_L g5270 ( 
.A1(n_5232),
.A2(n_5020),
.B(n_5037),
.Y(n_5270)
);

INVx1_ASAP7_75t_SL g5271 ( 
.A(n_5223),
.Y(n_5271)
);

AND2x2_ASAP7_75t_L g5272 ( 
.A(n_5214),
.B(n_4976),
.Y(n_5272)
);

NAND3xp33_ASAP7_75t_L g5273 ( 
.A(n_5231),
.B(n_5229),
.C(n_5146),
.Y(n_5273)
);

BUFx3_ASAP7_75t_L g5274 ( 
.A(n_5135),
.Y(n_5274)
);

BUFx6f_ASAP7_75t_L g5275 ( 
.A(n_5167),
.Y(n_5275)
);

INVx1_ASAP7_75t_L g5276 ( 
.A(n_5164),
.Y(n_5276)
);

AOI21xp5_ASAP7_75t_SL g5277 ( 
.A1(n_5203),
.A2(n_5033),
.B(n_5062),
.Y(n_5277)
);

OA21x2_ASAP7_75t_L g5278 ( 
.A1(n_5185),
.A2(n_5038),
.B(n_5026),
.Y(n_5278)
);

OR2x6_ASAP7_75t_L g5279 ( 
.A(n_5122),
.B(n_5064),
.Y(n_5279)
);

INVx2_ASAP7_75t_SL g5280 ( 
.A(n_5167),
.Y(n_5280)
);

BUFx6f_ASAP7_75t_L g5281 ( 
.A(n_5175),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_5165),
.Y(n_5282)
);

AO21x2_ASAP7_75t_L g5283 ( 
.A1(n_5224),
.A2(n_5107),
.B(n_4976),
.Y(n_5283)
);

OR2x2_ASAP7_75t_L g5284 ( 
.A(n_5180),
.B(n_300),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_5171),
.Y(n_5285)
);

INVx3_ASAP7_75t_SL g5286 ( 
.A(n_5207),
.Y(n_5286)
);

BUFx3_ASAP7_75t_L g5287 ( 
.A(n_5155),
.Y(n_5287)
);

INVx2_ASAP7_75t_L g5288 ( 
.A(n_5131),
.Y(n_5288)
);

NAND2xp5_ASAP7_75t_L g5289 ( 
.A(n_5159),
.B(n_300),
.Y(n_5289)
);

HB1xp67_ASAP7_75t_L g5290 ( 
.A(n_5126),
.Y(n_5290)
);

AND2x2_ASAP7_75t_L g5291 ( 
.A(n_5219),
.B(n_301),
.Y(n_5291)
);

INVx2_ASAP7_75t_L g5292 ( 
.A(n_5183),
.Y(n_5292)
);

INVx2_ASAP7_75t_L g5293 ( 
.A(n_5183),
.Y(n_5293)
);

NAND2xp5_ASAP7_75t_L g5294 ( 
.A(n_5136),
.B(n_302),
.Y(n_5294)
);

AND2x2_ASAP7_75t_L g5295 ( 
.A(n_5190),
.B(n_303),
.Y(n_5295)
);

AND2x2_ASAP7_75t_L g5296 ( 
.A(n_5249),
.B(n_305),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_5174),
.Y(n_5297)
);

AND2x2_ASAP7_75t_L g5298 ( 
.A(n_5187),
.B(n_305),
.Y(n_5298)
);

OR2x2_ASAP7_75t_L g5299 ( 
.A(n_5133),
.B(n_307),
.Y(n_5299)
);

AND2x2_ASAP7_75t_L g5300 ( 
.A(n_5238),
.B(n_307),
.Y(n_5300)
);

AND2x2_ASAP7_75t_L g5301 ( 
.A(n_5182),
.B(n_308),
.Y(n_5301)
);

AO21x2_ASAP7_75t_L g5302 ( 
.A1(n_5226),
.A2(n_308),
.B(n_309),
.Y(n_5302)
);

INVx1_ASAP7_75t_L g5303 ( 
.A(n_5178),
.Y(n_5303)
);

INVx1_ASAP7_75t_L g5304 ( 
.A(n_5184),
.Y(n_5304)
);

INVx2_ASAP7_75t_L g5305 ( 
.A(n_5183),
.Y(n_5305)
);

AND2x2_ASAP7_75t_L g5306 ( 
.A(n_5116),
.B(n_309),
.Y(n_5306)
);

INVx2_ASAP7_75t_L g5307 ( 
.A(n_5199),
.Y(n_5307)
);

AOI22xp33_ASAP7_75t_L g5308 ( 
.A1(n_5221),
.A2(n_5134),
.B1(n_5142),
.B2(n_5139),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_5197),
.Y(n_5309)
);

OAI21xp5_ASAP7_75t_L g5310 ( 
.A1(n_5256),
.A2(n_310),
.B(n_311),
.Y(n_5310)
);

INVx2_ASAP7_75t_L g5311 ( 
.A(n_5199),
.Y(n_5311)
);

INVx3_ASAP7_75t_L g5312 ( 
.A(n_5175),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_5198),
.Y(n_5313)
);

INVx2_ASAP7_75t_L g5314 ( 
.A(n_5140),
.Y(n_5314)
);

AND2x2_ASAP7_75t_L g5315 ( 
.A(n_5211),
.B(n_310),
.Y(n_5315)
);

INVx2_ASAP7_75t_L g5316 ( 
.A(n_5144),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_5201),
.Y(n_5317)
);

OAI21xp5_ASAP7_75t_L g5318 ( 
.A1(n_5191),
.A2(n_313),
.B(n_314),
.Y(n_5318)
);

AND2x4_ASAP7_75t_L g5319 ( 
.A(n_5211),
.B(n_314),
.Y(n_5319)
);

HB1xp67_ASAP7_75t_L g5320 ( 
.A(n_5143),
.Y(n_5320)
);

A2O1A1Ixp33_ASAP7_75t_L g5321 ( 
.A1(n_5153),
.A2(n_317),
.B(n_315),
.C(n_316),
.Y(n_5321)
);

NAND2xp5_ASAP7_75t_L g5322 ( 
.A(n_5141),
.B(n_316),
.Y(n_5322)
);

NOR2x1_ASAP7_75t_L g5323 ( 
.A(n_5175),
.B(n_318),
.Y(n_5323)
);

BUFx6f_ASAP7_75t_L g5324 ( 
.A(n_5206),
.Y(n_5324)
);

INVx2_ASAP7_75t_L g5325 ( 
.A(n_5202),
.Y(n_5325)
);

BUFx6f_ASAP7_75t_L g5326 ( 
.A(n_5253),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_5204),
.Y(n_5327)
);

HB1xp67_ASAP7_75t_L g5328 ( 
.A(n_5154),
.Y(n_5328)
);

NOR2x1_ASAP7_75t_L g5329 ( 
.A(n_5253),
.B(n_319),
.Y(n_5329)
);

AO21x2_ASAP7_75t_L g5330 ( 
.A1(n_5213),
.A2(n_319),
.B(n_320),
.Y(n_5330)
);

BUFx2_ASAP7_75t_L g5331 ( 
.A(n_5192),
.Y(n_5331)
);

OAI222xp33_ASAP7_75t_L g5332 ( 
.A1(n_5127),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.C1(n_325),
.C2(n_327),
.Y(n_5332)
);

HB1xp67_ASAP7_75t_L g5333 ( 
.A(n_5166),
.Y(n_5333)
);

INVx1_ASAP7_75t_L g5334 ( 
.A(n_5150),
.Y(n_5334)
);

AO21x2_ASAP7_75t_L g5335 ( 
.A1(n_5218),
.A2(n_325),
.B(n_329),
.Y(n_5335)
);

BUFx2_ASAP7_75t_L g5336 ( 
.A(n_5177),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_5160),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_5115),
.Y(n_5338)
);

OR2x2_ASAP7_75t_L g5339 ( 
.A(n_5151),
.B(n_329),
.Y(n_5339)
);

BUFx3_ASAP7_75t_L g5340 ( 
.A(n_5209),
.Y(n_5340)
);

INVx3_ASAP7_75t_L g5341 ( 
.A(n_5181),
.Y(n_5341)
);

AND2x2_ASAP7_75t_L g5342 ( 
.A(n_5217),
.B(n_330),
.Y(n_5342)
);

INVxp67_ASAP7_75t_L g5343 ( 
.A(n_5248),
.Y(n_5343)
);

AND2x2_ASAP7_75t_L g5344 ( 
.A(n_5168),
.B(n_330),
.Y(n_5344)
);

OR2x2_ASAP7_75t_L g5345 ( 
.A(n_5137),
.B(n_5220),
.Y(n_5345)
);

AOI21x1_ASAP7_75t_L g5346 ( 
.A1(n_5128),
.A2(n_5222),
.B(n_5170),
.Y(n_5346)
);

AOI22xp33_ASAP7_75t_SL g5347 ( 
.A1(n_5147),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_5179),
.Y(n_5348)
);

AND2x4_ASAP7_75t_SL g5349 ( 
.A(n_5128),
.B(n_331),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_5228),
.Y(n_5350)
);

AO21x2_ASAP7_75t_L g5351 ( 
.A1(n_5246),
.A2(n_332),
.B(n_334),
.Y(n_5351)
);

AND2x4_ASAP7_75t_L g5352 ( 
.A(n_5173),
.B(n_336),
.Y(n_5352)
);

INVx2_ASAP7_75t_L g5353 ( 
.A(n_5205),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5189),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_5196),
.Y(n_5355)
);

AO21x2_ASAP7_75t_L g5356 ( 
.A1(n_5193),
.A2(n_5212),
.B(n_5243),
.Y(n_5356)
);

BUFx3_ASAP7_75t_L g5357 ( 
.A(n_5209),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_5254),
.Y(n_5358)
);

INVxp67_ASAP7_75t_L g5359 ( 
.A(n_5176),
.Y(n_5359)
);

AOI21xp5_ASAP7_75t_SL g5360 ( 
.A1(n_5225),
.A2(n_337),
.B(n_338),
.Y(n_5360)
);

OA222x2_ASAP7_75t_L g5361 ( 
.A1(n_5132),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.C1(n_341),
.C2(n_342),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_5172),
.Y(n_5362)
);

OR2x2_ASAP7_75t_L g5363 ( 
.A(n_5215),
.B(n_343),
.Y(n_5363)
);

OR2x2_ASAP7_75t_L g5364 ( 
.A(n_5244),
.B(n_344),
.Y(n_5364)
);

OR2x6_ASAP7_75t_L g5365 ( 
.A(n_5225),
.B(n_344),
.Y(n_5365)
);

AO21x2_ASAP7_75t_L g5366 ( 
.A1(n_5148),
.A2(n_345),
.B(n_346),
.Y(n_5366)
);

BUFx2_ASAP7_75t_L g5367 ( 
.A(n_5130),
.Y(n_5367)
);

AND2x2_ASAP7_75t_L g5368 ( 
.A(n_5124),
.B(n_346),
.Y(n_5368)
);

OAI221xp5_ASAP7_75t_L g5369 ( 
.A1(n_5157),
.A2(n_350),
.B1(n_347),
.B2(n_348),
.C(n_351),
.Y(n_5369)
);

INVx1_ASAP7_75t_L g5370 ( 
.A(n_5333),
.Y(n_5370)
);

AND2x4_ASAP7_75t_SL g5371 ( 
.A(n_5326),
.B(n_5239),
.Y(n_5371)
);

HB1xp67_ASAP7_75t_L g5372 ( 
.A(n_5290),
.Y(n_5372)
);

INVx2_ASAP7_75t_L g5373 ( 
.A(n_5367),
.Y(n_5373)
);

INVx2_ASAP7_75t_L g5374 ( 
.A(n_5326),
.Y(n_5374)
);

INVx3_ASAP7_75t_L g5375 ( 
.A(n_5326),
.Y(n_5375)
);

AND2x2_ASAP7_75t_L g5376 ( 
.A(n_5340),
.B(n_5123),
.Y(n_5376)
);

INVx1_ASAP7_75t_L g5377 ( 
.A(n_5333),
.Y(n_5377)
);

INVx2_ASAP7_75t_L g5378 ( 
.A(n_5264),
.Y(n_5378)
);

INVx2_ASAP7_75t_L g5379 ( 
.A(n_5264),
.Y(n_5379)
);

NOR2xp33_ASAP7_75t_L g5380 ( 
.A(n_5343),
.B(n_5195),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_5328),
.Y(n_5381)
);

OAI22xp5_ASAP7_75t_L g5382 ( 
.A1(n_5308),
.A2(n_5129),
.B1(n_5194),
.B2(n_5161),
.Y(n_5382)
);

AND2x2_ASAP7_75t_L g5383 ( 
.A(n_5340),
.B(n_5210),
.Y(n_5383)
);

INVx1_ASAP7_75t_SL g5384 ( 
.A(n_5286),
.Y(n_5384)
);

NAND2xp5_ASAP7_75t_L g5385 ( 
.A(n_5359),
.B(n_5241),
.Y(n_5385)
);

INVx2_ASAP7_75t_L g5386 ( 
.A(n_5290),
.Y(n_5386)
);

INVx1_ASAP7_75t_L g5387 ( 
.A(n_5328),
.Y(n_5387)
);

NOR2xp33_ASAP7_75t_L g5388 ( 
.A(n_5343),
.B(n_5162),
.Y(n_5388)
);

INVx2_ASAP7_75t_L g5389 ( 
.A(n_5320),
.Y(n_5389)
);

BUFx3_ASAP7_75t_L g5390 ( 
.A(n_5324),
.Y(n_5390)
);

AND2x2_ASAP7_75t_L g5391 ( 
.A(n_5357),
.B(n_5210),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_5320),
.Y(n_5392)
);

OAI22xp5_ASAP7_75t_L g5393 ( 
.A1(n_5308),
.A2(n_5236),
.B1(n_5235),
.B2(n_5239),
.Y(n_5393)
);

AND2x2_ASAP7_75t_L g5394 ( 
.A(n_5263),
.B(n_5163),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_5258),
.Y(n_5395)
);

OAI21xp5_ASAP7_75t_L g5396 ( 
.A1(n_5273),
.A2(n_5230),
.B(n_5227),
.Y(n_5396)
);

NAND2xp5_ASAP7_75t_L g5397 ( 
.A(n_5359),
.B(n_5257),
.Y(n_5397)
);

OR2x2_ASAP7_75t_L g5398 ( 
.A(n_5345),
.B(n_5186),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_5268),
.Y(n_5399)
);

NAND2xp5_ASAP7_75t_L g5400 ( 
.A(n_5294),
.B(n_5255),
.Y(n_5400)
);

OAI21xp5_ASAP7_75t_SL g5401 ( 
.A1(n_5273),
.A2(n_5310),
.B(n_5347),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_5276),
.Y(n_5402)
);

NAND2xp5_ASAP7_75t_L g5403 ( 
.A(n_5294),
.B(n_5255),
.Y(n_5403)
);

INVx2_ASAP7_75t_L g5404 ( 
.A(n_5316),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5282),
.Y(n_5405)
);

BUFx2_ASAP7_75t_L g5406 ( 
.A(n_5331),
.Y(n_5406)
);

INVx1_ASAP7_75t_L g5407 ( 
.A(n_5285),
.Y(n_5407)
);

AND2x4_ASAP7_75t_L g5408 ( 
.A(n_5266),
.B(n_5252),
.Y(n_5408)
);

HB1xp67_ASAP7_75t_L g5409 ( 
.A(n_5354),
.Y(n_5409)
);

AND2x4_ASAP7_75t_L g5410 ( 
.A(n_5266),
.B(n_5252),
.Y(n_5410)
);

AND2x2_ASAP7_75t_L g5411 ( 
.A(n_5357),
.B(n_5188),
.Y(n_5411)
);

NAND2xp5_ASAP7_75t_L g5412 ( 
.A(n_5265),
.B(n_5255),
.Y(n_5412)
);

AND2x2_ASAP7_75t_L g5413 ( 
.A(n_5288),
.B(n_5118),
.Y(n_5413)
);

AND2x2_ASAP7_75t_L g5414 ( 
.A(n_5312),
.B(n_5307),
.Y(n_5414)
);

HB1xp67_ASAP7_75t_L g5415 ( 
.A(n_5362),
.Y(n_5415)
);

BUFx2_ASAP7_75t_L g5416 ( 
.A(n_5269),
.Y(n_5416)
);

AND2x2_ASAP7_75t_L g5417 ( 
.A(n_5312),
.B(n_5120),
.Y(n_5417)
);

AND2x2_ASAP7_75t_L g5418 ( 
.A(n_5346),
.B(n_5250),
.Y(n_5418)
);

NAND2xp5_ASAP7_75t_L g5419 ( 
.A(n_5265),
.B(n_5239),
.Y(n_5419)
);

AND2x4_ASAP7_75t_L g5420 ( 
.A(n_5260),
.B(n_5117),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_5297),
.Y(n_5421)
);

AOI22xp33_ASAP7_75t_L g5422 ( 
.A1(n_5356),
.A2(n_5156),
.B1(n_5247),
.B2(n_5240),
.Y(n_5422)
);

INVx2_ASAP7_75t_L g5423 ( 
.A(n_5275),
.Y(n_5423)
);

NAND2xp5_ASAP7_75t_SL g5424 ( 
.A(n_5318),
.B(n_5152),
.Y(n_5424)
);

NAND2xp5_ASAP7_75t_L g5425 ( 
.A(n_5270),
.B(n_5200),
.Y(n_5425)
);

OR2x2_ASAP7_75t_L g5426 ( 
.A(n_5338),
.B(n_5208),
.Y(n_5426)
);

CKINVDCx8_ASAP7_75t_R g5427 ( 
.A(n_5365),
.Y(n_5427)
);

INVx2_ASAP7_75t_L g5428 ( 
.A(n_5275),
.Y(n_5428)
);

OR2x2_ASAP7_75t_L g5429 ( 
.A(n_5314),
.B(n_5117),
.Y(n_5429)
);

AOI22xp33_ASAP7_75t_SL g5430 ( 
.A1(n_5356),
.A2(n_5233),
.B1(n_5149),
.B2(n_5145),
.Y(n_5430)
);

INVx1_ASAP7_75t_SL g5431 ( 
.A(n_5286),
.Y(n_5431)
);

AOI22xp33_ASAP7_75t_SL g5432 ( 
.A1(n_5270),
.A2(n_5242),
.B1(n_5117),
.B2(n_5216),
.Y(n_5432)
);

BUFx2_ASAP7_75t_L g5433 ( 
.A(n_5269),
.Y(n_5433)
);

AND2x2_ASAP7_75t_L g5434 ( 
.A(n_5341),
.B(n_5121),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5303),
.Y(n_5435)
);

AOI222xp33_ASAP7_75t_L g5436 ( 
.A1(n_5310),
.A2(n_5369),
.B1(n_5318),
.B2(n_5332),
.C1(n_5321),
.C2(n_5289),
.Y(n_5436)
);

AOI22xp33_ASAP7_75t_L g5437 ( 
.A1(n_5369),
.A2(n_5242),
.B1(n_353),
.B2(n_347),
.Y(n_5437)
);

AND2x2_ASAP7_75t_L g5438 ( 
.A(n_5341),
.B(n_5121),
.Y(n_5438)
);

AND2x4_ASAP7_75t_L g5439 ( 
.A(n_5280),
.B(n_5121),
.Y(n_5439)
);

INVx2_ASAP7_75t_L g5440 ( 
.A(n_5275),
.Y(n_5440)
);

INVx1_ASAP7_75t_SL g5441 ( 
.A(n_5271),
.Y(n_5441)
);

AND2x2_ASAP7_75t_L g5442 ( 
.A(n_5336),
.B(n_5242),
.Y(n_5442)
);

INVx2_ASAP7_75t_L g5443 ( 
.A(n_5281),
.Y(n_5443)
);

AOI22xp33_ASAP7_75t_L g5444 ( 
.A1(n_5422),
.A2(n_5347),
.B1(n_5279),
.B2(n_5351),
.Y(n_5444)
);

BUFx3_ASAP7_75t_L g5445 ( 
.A(n_5406),
.Y(n_5445)
);

AND2x2_ASAP7_75t_L g5446 ( 
.A(n_5376),
.B(n_5274),
.Y(n_5446)
);

BUFx3_ASAP7_75t_L g5447 ( 
.A(n_5390),
.Y(n_5447)
);

INVx3_ASAP7_75t_L g5448 ( 
.A(n_5390),
.Y(n_5448)
);

INVx3_ASAP7_75t_L g5449 ( 
.A(n_5371),
.Y(n_5449)
);

AND2x2_ASAP7_75t_L g5450 ( 
.A(n_5373),
.B(n_5274),
.Y(n_5450)
);

AND2x2_ASAP7_75t_L g5451 ( 
.A(n_5373),
.B(n_5287),
.Y(n_5451)
);

NAND2xp5_ASAP7_75t_SL g5452 ( 
.A(n_5436),
.B(n_5281),
.Y(n_5452)
);

AO21x1_ASAP7_75t_SL g5453 ( 
.A1(n_5419),
.A2(n_5332),
.B(n_5350),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_5372),
.Y(n_5454)
);

OAI211xp5_ASAP7_75t_L g5455 ( 
.A1(n_5401),
.A2(n_5321),
.B(n_5267),
.C(n_5277),
.Y(n_5455)
);

AND2x2_ASAP7_75t_L g5456 ( 
.A(n_5388),
.B(n_5287),
.Y(n_5456)
);

AO21x2_ASAP7_75t_L g5457 ( 
.A1(n_5412),
.A2(n_5289),
.B(n_5292),
.Y(n_5457)
);

NAND4xp25_ASAP7_75t_SL g5458 ( 
.A(n_5422),
.B(n_5267),
.C(n_5360),
.D(n_5271),
.Y(n_5458)
);

NAND3xp33_ASAP7_75t_L g5459 ( 
.A(n_5437),
.B(n_5279),
.C(n_5329),
.Y(n_5459)
);

AND2x2_ASAP7_75t_L g5460 ( 
.A(n_5388),
.B(n_5281),
.Y(n_5460)
);

AOI22xp33_ASAP7_75t_SL g5461 ( 
.A1(n_5382),
.A2(n_5278),
.B1(n_5330),
.B2(n_5279),
.Y(n_5461)
);

INVx2_ASAP7_75t_L g5462 ( 
.A(n_5375),
.Y(n_5462)
);

INVx1_ASAP7_75t_L g5463 ( 
.A(n_5372),
.Y(n_5463)
);

HB1xp67_ASAP7_75t_L g5464 ( 
.A(n_5386),
.Y(n_5464)
);

NAND2xp5_ASAP7_75t_L g5465 ( 
.A(n_5380),
.B(n_5330),
.Y(n_5465)
);

OR2x6_ASAP7_75t_L g5466 ( 
.A(n_5416),
.B(n_5259),
.Y(n_5466)
);

HB1xp67_ASAP7_75t_L g5467 ( 
.A(n_5386),
.Y(n_5467)
);

NAND2xp5_ASAP7_75t_L g5468 ( 
.A(n_5380),
.B(n_5441),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_5389),
.Y(n_5469)
);

NOR2xp33_ASAP7_75t_R g5470 ( 
.A(n_5427),
.B(n_5259),
.Y(n_5470)
);

HB1xp67_ASAP7_75t_L g5471 ( 
.A(n_5389),
.Y(n_5471)
);

INVx5_ASAP7_75t_L g5472 ( 
.A(n_5375),
.Y(n_5472)
);

AND2x4_ASAP7_75t_SL g5473 ( 
.A(n_5408),
.B(n_5262),
.Y(n_5473)
);

AOI22xp33_ASAP7_75t_L g5474 ( 
.A1(n_5424),
.A2(n_5351),
.B1(n_5366),
.B2(n_5298),
.Y(n_5474)
);

INVx3_ASAP7_75t_L g5475 ( 
.A(n_5371),
.Y(n_5475)
);

OAI211xp5_ASAP7_75t_SL g5476 ( 
.A1(n_5396),
.A2(n_5322),
.B(n_5323),
.C(n_5358),
.Y(n_5476)
);

AND2x4_ASAP7_75t_L g5477 ( 
.A(n_5375),
.B(n_5262),
.Y(n_5477)
);

INVx5_ASAP7_75t_L g5478 ( 
.A(n_5433),
.Y(n_5478)
);

OAI21xp5_ASAP7_75t_L g5479 ( 
.A1(n_5424),
.A2(n_5278),
.B(n_5262),
.Y(n_5479)
);

AOI22xp33_ASAP7_75t_L g5480 ( 
.A1(n_5430),
.A2(n_5366),
.B1(n_5283),
.B2(n_5291),
.Y(n_5480)
);

INVx2_ASAP7_75t_L g5481 ( 
.A(n_5427),
.Y(n_5481)
);

OAI22xp5_ASAP7_75t_L g5482 ( 
.A1(n_5437),
.A2(n_5311),
.B1(n_5337),
.B2(n_5334),
.Y(n_5482)
);

OAI211xp5_ASAP7_75t_L g5483 ( 
.A1(n_5432),
.A2(n_5322),
.B(n_5293),
.C(n_5305),
.Y(n_5483)
);

AOI22xp33_ASAP7_75t_L g5484 ( 
.A1(n_5393),
.A2(n_5283),
.B1(n_5335),
.B2(n_5302),
.Y(n_5484)
);

NAND3xp33_ASAP7_75t_SL g5485 ( 
.A(n_5442),
.B(n_5284),
.C(n_5306),
.Y(n_5485)
);

OAI221xp5_ASAP7_75t_L g5486 ( 
.A1(n_5385),
.A2(n_5365),
.B1(n_5272),
.B2(n_5339),
.C(n_5299),
.Y(n_5486)
);

AND2x4_ASAP7_75t_L g5487 ( 
.A(n_5383),
.B(n_5349),
.Y(n_5487)
);

AOI221xp5_ASAP7_75t_L g5488 ( 
.A1(n_5409),
.A2(n_5335),
.B1(n_5302),
.B2(n_5296),
.C(n_5352),
.Y(n_5488)
);

INVx2_ASAP7_75t_L g5489 ( 
.A(n_5408),
.Y(n_5489)
);

INVx1_ASAP7_75t_L g5490 ( 
.A(n_5464),
.Y(n_5490)
);

AND2x2_ASAP7_75t_L g5491 ( 
.A(n_5456),
.B(n_5394),
.Y(n_5491)
);

INVx2_ASAP7_75t_L g5492 ( 
.A(n_5478),
.Y(n_5492)
);

BUFx2_ASAP7_75t_L g5493 ( 
.A(n_5470),
.Y(n_5493)
);

OR2x2_ASAP7_75t_L g5494 ( 
.A(n_5454),
.B(n_5370),
.Y(n_5494)
);

INVxp33_ASAP7_75t_L g5495 ( 
.A(n_5470),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5464),
.Y(n_5496)
);

NAND2xp5_ASAP7_75t_L g5497 ( 
.A(n_5445),
.B(n_5481),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_5467),
.Y(n_5498)
);

AND2x2_ASAP7_75t_L g5499 ( 
.A(n_5446),
.B(n_5394),
.Y(n_5499)
);

AND2x2_ASAP7_75t_L g5500 ( 
.A(n_5451),
.B(n_5414),
.Y(n_5500)
);

INVx5_ASAP7_75t_L g5501 ( 
.A(n_5466),
.Y(n_5501)
);

AND2x2_ASAP7_75t_L g5502 ( 
.A(n_5460),
.B(n_5414),
.Y(n_5502)
);

INVx2_ASAP7_75t_L g5503 ( 
.A(n_5478),
.Y(n_5503)
);

HB1xp67_ASAP7_75t_L g5504 ( 
.A(n_5478),
.Y(n_5504)
);

NAND2xp5_ASAP7_75t_L g5505 ( 
.A(n_5445),
.B(n_5374),
.Y(n_5505)
);

AND2x2_ASAP7_75t_L g5506 ( 
.A(n_5466),
.B(n_5449),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_5467),
.Y(n_5507)
);

INVx1_ASAP7_75t_L g5508 ( 
.A(n_5471),
.Y(n_5508)
);

NAND2xp5_ASAP7_75t_L g5509 ( 
.A(n_5481),
.B(n_5374),
.Y(n_5509)
);

INVx2_ASAP7_75t_L g5510 ( 
.A(n_5478),
.Y(n_5510)
);

INVx1_ASAP7_75t_L g5511 ( 
.A(n_5471),
.Y(n_5511)
);

INVx1_ASAP7_75t_L g5512 ( 
.A(n_5463),
.Y(n_5512)
);

AND2x2_ASAP7_75t_L g5513 ( 
.A(n_5466),
.B(n_5423),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_5469),
.Y(n_5514)
);

AND2x4_ASAP7_75t_L g5515 ( 
.A(n_5472),
.B(n_5423),
.Y(n_5515)
);

AND2x2_ASAP7_75t_L g5516 ( 
.A(n_5449),
.B(n_5428),
.Y(n_5516)
);

AND2x2_ASAP7_75t_L g5517 ( 
.A(n_5475),
.B(n_5428),
.Y(n_5517)
);

INVx1_ASAP7_75t_L g5518 ( 
.A(n_5462),
.Y(n_5518)
);

NAND3xp33_ASAP7_75t_L g5519 ( 
.A(n_5461),
.B(n_5381),
.C(n_5377),
.Y(n_5519)
);

INVx1_ASAP7_75t_L g5520 ( 
.A(n_5462),
.Y(n_5520)
);

AND2x2_ASAP7_75t_L g5521 ( 
.A(n_5475),
.B(n_5448),
.Y(n_5521)
);

NAND2xp5_ASAP7_75t_L g5522 ( 
.A(n_5474),
.B(n_5440),
.Y(n_5522)
);

NOR2xp33_ASAP7_75t_L g5523 ( 
.A(n_5495),
.B(n_5455),
.Y(n_5523)
);

AND2x2_ASAP7_75t_L g5524 ( 
.A(n_5491),
.B(n_5487),
.Y(n_5524)
);

OR2x2_ASAP7_75t_L g5525 ( 
.A(n_5509),
.B(n_5485),
.Y(n_5525)
);

OR2x2_ASAP7_75t_L g5526 ( 
.A(n_5497),
.B(n_5468),
.Y(n_5526)
);

AND2x2_ASAP7_75t_L g5527 ( 
.A(n_5491),
.B(n_5487),
.Y(n_5527)
);

NAND2xp5_ASAP7_75t_L g5528 ( 
.A(n_5516),
.B(n_5517),
.Y(n_5528)
);

AND2x2_ASAP7_75t_SL g5529 ( 
.A(n_5493),
.B(n_5480),
.Y(n_5529)
);

HB1xp67_ASAP7_75t_L g5530 ( 
.A(n_5504),
.Y(n_5530)
);

INVx1_ASAP7_75t_L g5531 ( 
.A(n_5490),
.Y(n_5531)
);

AND2x2_ASAP7_75t_L g5532 ( 
.A(n_5499),
.B(n_5448),
.Y(n_5532)
);

INVx1_ASAP7_75t_SL g5533 ( 
.A(n_5493),
.Y(n_5533)
);

NAND2x1_ASAP7_75t_L g5534 ( 
.A(n_5515),
.B(n_5477),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_5490),
.Y(n_5535)
);

NAND2xp5_ASAP7_75t_L g5536 ( 
.A(n_5516),
.B(n_5474),
.Y(n_5536)
);

AND2x4_ASAP7_75t_L g5537 ( 
.A(n_5501),
.B(n_5515),
.Y(n_5537)
);

NAND2xp5_ASAP7_75t_L g5538 ( 
.A(n_5517),
.B(n_5447),
.Y(n_5538)
);

AND2x2_ASAP7_75t_L g5539 ( 
.A(n_5499),
.B(n_5450),
.Y(n_5539)
);

BUFx2_ASAP7_75t_SL g5540 ( 
.A(n_5501),
.Y(n_5540)
);

NAND2xp5_ASAP7_75t_L g5541 ( 
.A(n_5521),
.B(n_5447),
.Y(n_5541)
);

INVx2_ASAP7_75t_L g5542 ( 
.A(n_5501),
.Y(n_5542)
);

INVx2_ASAP7_75t_L g5543 ( 
.A(n_5501),
.Y(n_5543)
);

AND2x2_ASAP7_75t_L g5544 ( 
.A(n_5502),
.B(n_5391),
.Y(n_5544)
);

NAND2xp5_ASAP7_75t_L g5545 ( 
.A(n_5521),
.B(n_5500),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_5530),
.Y(n_5546)
);

NAND2xp5_ASAP7_75t_L g5547 ( 
.A(n_5532),
.B(n_5533),
.Y(n_5547)
);

INVx1_ASAP7_75t_L g5548 ( 
.A(n_5530),
.Y(n_5548)
);

AND2x2_ASAP7_75t_L g5549 ( 
.A(n_5532),
.B(n_5502),
.Y(n_5549)
);

OR2x2_ASAP7_75t_L g5550 ( 
.A(n_5528),
.B(n_5452),
.Y(n_5550)
);

OAI21xp33_ASAP7_75t_L g5551 ( 
.A1(n_5529),
.A2(n_5452),
.B(n_5458),
.Y(n_5551)
);

INVx1_ASAP7_75t_SL g5552 ( 
.A(n_5540),
.Y(n_5552)
);

OR2x2_ASAP7_75t_L g5553 ( 
.A(n_5536),
.B(n_5522),
.Y(n_5553)
);

AND2x2_ASAP7_75t_L g5554 ( 
.A(n_5544),
.B(n_5500),
.Y(n_5554)
);

INVx2_ASAP7_75t_L g5555 ( 
.A(n_5537),
.Y(n_5555)
);

OAI211xp5_ASAP7_75t_L g5556 ( 
.A1(n_5523),
.A2(n_5480),
.B(n_5519),
.C(n_5483),
.Y(n_5556)
);

AOI22xp33_ASAP7_75t_SL g5557 ( 
.A1(n_5529),
.A2(n_5479),
.B1(n_5459),
.B2(n_5473),
.Y(n_5557)
);

OAI21xp5_ASAP7_75t_L g5558 ( 
.A1(n_5523),
.A2(n_5444),
.B(n_5484),
.Y(n_5558)
);

INVx2_ASAP7_75t_L g5559 ( 
.A(n_5537),
.Y(n_5559)
);

NOR2xp33_ASAP7_75t_L g5560 ( 
.A(n_5541),
.B(n_5495),
.Y(n_5560)
);

NAND2xp5_ASAP7_75t_L g5561 ( 
.A(n_5539),
.B(n_5513),
.Y(n_5561)
);

OR2x2_ASAP7_75t_L g5562 ( 
.A(n_5545),
.B(n_5465),
.Y(n_5562)
);

INVx1_ASAP7_75t_L g5563 ( 
.A(n_5531),
.Y(n_5563)
);

OR2x2_ASAP7_75t_L g5564 ( 
.A(n_5525),
.B(n_5505),
.Y(n_5564)
);

OR2x2_ASAP7_75t_L g5565 ( 
.A(n_5526),
.B(n_5397),
.Y(n_5565)
);

NAND2xp5_ASAP7_75t_SL g5566 ( 
.A(n_5537),
.B(n_5501),
.Y(n_5566)
);

OR2x2_ASAP7_75t_L g5567 ( 
.A(n_5538),
.B(n_5494),
.Y(n_5567)
);

INVx2_ASAP7_75t_L g5568 ( 
.A(n_5534),
.Y(n_5568)
);

OAI22xp5_ASAP7_75t_L g5569 ( 
.A1(n_5557),
.A2(n_5444),
.B1(n_5484),
.B2(n_5556),
.Y(n_5569)
);

AOI32xp33_ASAP7_75t_L g5570 ( 
.A1(n_5551),
.A2(n_5476),
.A3(n_5506),
.B1(n_5488),
.B2(n_5482),
.Y(n_5570)
);

OAI32xp33_ASAP7_75t_L g5571 ( 
.A1(n_5551),
.A2(n_5425),
.A3(n_5453),
.B1(n_5378),
.B2(n_5379),
.Y(n_5571)
);

AO21x1_ASAP7_75t_L g5572 ( 
.A1(n_5558),
.A2(n_5515),
.B(n_5503),
.Y(n_5572)
);

AND2x2_ASAP7_75t_L g5573 ( 
.A(n_5549),
.B(n_5506),
.Y(n_5573)
);

INVx1_ASAP7_75t_L g5574 ( 
.A(n_5547),
.Y(n_5574)
);

BUFx2_ASAP7_75t_L g5575 ( 
.A(n_5568),
.Y(n_5575)
);

OAI22xp33_ASAP7_75t_L g5576 ( 
.A1(n_5558),
.A2(n_5472),
.B1(n_5378),
.B2(n_5379),
.Y(n_5576)
);

INVx1_ASAP7_75t_L g5577 ( 
.A(n_5546),
.Y(n_5577)
);

NOR3xp33_ASAP7_75t_L g5578 ( 
.A(n_5560),
.B(n_5543),
.C(n_5542),
.Y(n_5578)
);

INVx1_ASAP7_75t_L g5579 ( 
.A(n_5548),
.Y(n_5579)
);

NOR2x1_ASAP7_75t_L g5580 ( 
.A(n_5566),
.B(n_5492),
.Y(n_5580)
);

OAI22xp5_ASAP7_75t_L g5581 ( 
.A1(n_5553),
.A2(n_5431),
.B1(n_5384),
.B2(n_5486),
.Y(n_5581)
);

AND2x4_ASAP7_75t_L g5582 ( 
.A(n_5555),
.B(n_5559),
.Y(n_5582)
);

OR2x2_ASAP7_75t_L g5583 ( 
.A(n_5550),
.B(n_5494),
.Y(n_5583)
);

NAND2xp5_ASAP7_75t_L g5584 ( 
.A(n_5554),
.B(n_5552),
.Y(n_5584)
);

O2A1O1Ixp33_ASAP7_75t_L g5585 ( 
.A1(n_5552),
.A2(n_5503),
.B(n_5510),
.C(n_5492),
.Y(n_5585)
);

NAND2xp5_ASAP7_75t_L g5586 ( 
.A(n_5573),
.B(n_5524),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_5582),
.Y(n_5587)
);

INVx1_ASAP7_75t_SL g5588 ( 
.A(n_5583),
.Y(n_5588)
);

OR2x2_ASAP7_75t_L g5589 ( 
.A(n_5584),
.B(n_5567),
.Y(n_5589)
);

OR2x2_ASAP7_75t_L g5590 ( 
.A(n_5582),
.B(n_5561),
.Y(n_5590)
);

AND2x2_ASAP7_75t_L g5591 ( 
.A(n_5575),
.B(n_5527),
.Y(n_5591)
);

AND2x2_ASAP7_75t_SL g5592 ( 
.A(n_5578),
.B(n_5564),
.Y(n_5592)
);

OR2x2_ASAP7_75t_L g5593 ( 
.A(n_5574),
.B(n_5565),
.Y(n_5593)
);

CKINVDCx16_ASAP7_75t_R g5594 ( 
.A(n_5580),
.Y(n_5594)
);

AND2x4_ASAP7_75t_L g5595 ( 
.A(n_5577),
.B(n_5542),
.Y(n_5595)
);

INVx1_ASAP7_75t_SL g5596 ( 
.A(n_5579),
.Y(n_5596)
);

NOR2x1_ASAP7_75t_L g5597 ( 
.A(n_5585),
.B(n_5543),
.Y(n_5597)
);

AND2x2_ASAP7_75t_L g5598 ( 
.A(n_5581),
.B(n_5513),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_5590),
.Y(n_5599)
);

INVx2_ASAP7_75t_L g5600 ( 
.A(n_5591),
.Y(n_5600)
);

OAI22xp5_ASAP7_75t_L g5601 ( 
.A1(n_5594),
.A2(n_5569),
.B1(n_5489),
.B2(n_5570),
.Y(n_5601)
);

OAI322xp33_ASAP7_75t_L g5602 ( 
.A1(n_5596),
.A2(n_5576),
.A3(n_5496),
.B1(n_5498),
.B2(n_5507),
.C1(n_5508),
.C2(n_5511),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_5597),
.Y(n_5603)
);

INVx2_ASAP7_75t_SL g5604 ( 
.A(n_5587),
.Y(n_5604)
);

NOR3xp33_ASAP7_75t_L g5605 ( 
.A(n_5588),
.B(n_5562),
.C(n_5571),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_5589),
.Y(n_5606)
);

AOI22xp5_ASAP7_75t_L g5607 ( 
.A1(n_5592),
.A2(n_5572),
.B1(n_5510),
.B2(n_5512),
.Y(n_5607)
);

OAI21xp33_ASAP7_75t_L g5608 ( 
.A1(n_5586),
.A2(n_5473),
.B(n_5477),
.Y(n_5608)
);

INVxp67_ASAP7_75t_SL g5609 ( 
.A(n_5598),
.Y(n_5609)
);

NAND2xp5_ASAP7_75t_L g5610 ( 
.A(n_5595),
.B(n_5535),
.Y(n_5610)
);

INVxp67_ASAP7_75t_SL g5611 ( 
.A(n_5593),
.Y(n_5611)
);

INVx1_ASAP7_75t_SL g5612 ( 
.A(n_5595),
.Y(n_5612)
);

INVx2_ASAP7_75t_L g5613 ( 
.A(n_5591),
.Y(n_5613)
);

INVx1_ASAP7_75t_L g5614 ( 
.A(n_5609),
.Y(n_5614)
);

O2A1O1Ixp5_ASAP7_75t_L g5615 ( 
.A1(n_5603),
.A2(n_5518),
.B(n_5520),
.C(n_5563),
.Y(n_5615)
);

NAND2xp5_ASAP7_75t_L g5616 ( 
.A(n_5612),
.B(n_5514),
.Y(n_5616)
);

INVx1_ASAP7_75t_SL g5617 ( 
.A(n_5600),
.Y(n_5617)
);

INVx1_ASAP7_75t_L g5618 ( 
.A(n_5610),
.Y(n_5618)
);

AND2x4_ASAP7_75t_L g5619 ( 
.A(n_5613),
.B(n_5440),
.Y(n_5619)
);

NAND2xp5_ASAP7_75t_L g5620 ( 
.A(n_5607),
.B(n_5604),
.Y(n_5620)
);

AND2x2_ASAP7_75t_L g5621 ( 
.A(n_5611),
.B(n_5404),
.Y(n_5621)
);

INVx2_ASAP7_75t_SL g5622 ( 
.A(n_5599),
.Y(n_5622)
);

OAI21xp33_ASAP7_75t_L g5623 ( 
.A1(n_5608),
.A2(n_5392),
.B(n_5387),
.Y(n_5623)
);

AOI22xp5_ASAP7_75t_L g5624 ( 
.A1(n_5601),
.A2(n_5443),
.B1(n_5457),
.B2(n_5472),
.Y(n_5624)
);

OAI22xp5_ASAP7_75t_L g5625 ( 
.A1(n_5617),
.A2(n_5607),
.B1(n_5606),
.B2(n_5472),
.Y(n_5625)
);

NAND2xp5_ASAP7_75t_L g5626 ( 
.A(n_5621),
.B(n_5605),
.Y(n_5626)
);

NAND2xp5_ASAP7_75t_L g5627 ( 
.A(n_5619),
.B(n_5415),
.Y(n_5627)
);

NAND2x1_ASAP7_75t_L g5628 ( 
.A(n_5614),
.B(n_5443),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_5620),
.Y(n_5629)
);

NAND2xp5_ASAP7_75t_L g5630 ( 
.A(n_5622),
.B(n_5624),
.Y(n_5630)
);

AND2x2_ASAP7_75t_L g5631 ( 
.A(n_5623),
.B(n_5415),
.Y(n_5631)
);

NAND2xp5_ASAP7_75t_L g5632 ( 
.A(n_5616),
.B(n_5409),
.Y(n_5632)
);

INVx1_ASAP7_75t_L g5633 ( 
.A(n_5615),
.Y(n_5633)
);

INVx1_ASAP7_75t_SL g5634 ( 
.A(n_5618),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_5621),
.Y(n_5635)
);

HB1xp67_ASAP7_75t_L g5636 ( 
.A(n_5628),
.Y(n_5636)
);

AOI222xp33_ASAP7_75t_L g5637 ( 
.A1(n_5633),
.A2(n_5602),
.B1(n_5404),
.B2(n_5403),
.C1(n_5400),
.C2(n_5457),
.Y(n_5637)
);

AOI221xp5_ASAP7_75t_L g5638 ( 
.A1(n_5625),
.A2(n_5629),
.B1(n_5626),
.B2(n_5631),
.C(n_5635),
.Y(n_5638)
);

INVx1_ASAP7_75t_L g5639 ( 
.A(n_5627),
.Y(n_5639)
);

INVx2_ASAP7_75t_L g5640 ( 
.A(n_5632),
.Y(n_5640)
);

AOI22xp5_ASAP7_75t_L g5641 ( 
.A1(n_5634),
.A2(n_5410),
.B1(n_5408),
.B2(n_5434),
.Y(n_5641)
);

NOR2xp67_ASAP7_75t_SL g5642 ( 
.A(n_5630),
.B(n_5324),
.Y(n_5642)
);

AOI221xp5_ASAP7_75t_L g5643 ( 
.A1(n_5625),
.A2(n_5438),
.B1(n_5319),
.B2(n_5324),
.C(n_5407),
.Y(n_5643)
);

INVx2_ASAP7_75t_L g5644 ( 
.A(n_5628),
.Y(n_5644)
);

NAND3xp33_ASAP7_75t_L g5645 ( 
.A(n_5625),
.B(n_5365),
.C(n_5405),
.Y(n_5645)
);

AOI22xp33_ASAP7_75t_SL g5646 ( 
.A1(n_5631),
.A2(n_5349),
.B1(n_5319),
.B2(n_5439),
.Y(n_5646)
);

AOI21xp5_ASAP7_75t_L g5647 ( 
.A1(n_5626),
.A2(n_5410),
.B(n_5421),
.Y(n_5647)
);

AOI21xp5_ASAP7_75t_L g5648 ( 
.A1(n_5626),
.A2(n_5410),
.B(n_5435),
.Y(n_5648)
);

AOI21xp5_ASAP7_75t_L g5649 ( 
.A1(n_5626),
.A2(n_5439),
.B(n_5399),
.Y(n_5649)
);

AOI221xp5_ASAP7_75t_L g5650 ( 
.A1(n_5625),
.A2(n_5439),
.B1(n_5402),
.B2(n_5395),
.C(n_5315),
.Y(n_5650)
);

NAND3xp33_ASAP7_75t_SL g5651 ( 
.A(n_5626),
.B(n_5418),
.C(n_5344),
.Y(n_5651)
);

OA21x2_ASAP7_75t_L g5652 ( 
.A1(n_5626),
.A2(n_5417),
.B(n_5420),
.Y(n_5652)
);

INVx1_ASAP7_75t_SL g5653 ( 
.A(n_5627),
.Y(n_5653)
);

NOR2x1_ASAP7_75t_L g5654 ( 
.A(n_5625),
.B(n_5352),
.Y(n_5654)
);

NOR2xp67_ASAP7_75t_L g5655 ( 
.A(n_5636),
.B(n_352),
.Y(n_5655)
);

INVx1_ASAP7_75t_L g5656 ( 
.A(n_5644),
.Y(n_5656)
);

INVxp67_ASAP7_75t_SL g5657 ( 
.A(n_5642),
.Y(n_5657)
);

NAND2xp5_ASAP7_75t_L g5658 ( 
.A(n_5641),
.B(n_5295),
.Y(n_5658)
);

AOI221xp5_ASAP7_75t_L g5659 ( 
.A1(n_5643),
.A2(n_5420),
.B1(n_5301),
.B2(n_5300),
.C(n_5342),
.Y(n_5659)
);

AOI22xp33_ASAP7_75t_L g5660 ( 
.A1(n_5651),
.A2(n_5646),
.B1(n_5645),
.B2(n_5654),
.Y(n_5660)
);

AOI22xp33_ASAP7_75t_L g5661 ( 
.A1(n_5637),
.A2(n_5420),
.B1(n_5417),
.B2(n_5368),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5652),
.Y(n_5662)
);

NAND2xp5_ASAP7_75t_L g5663 ( 
.A(n_5647),
.B(n_5648),
.Y(n_5663)
);

NAND2xp33_ASAP7_75t_L g5664 ( 
.A(n_5653),
.B(n_5640),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_5652),
.Y(n_5665)
);

NOR2x1_ASAP7_75t_L g5666 ( 
.A(n_5639),
.B(n_5364),
.Y(n_5666)
);

NAND4xp25_ASAP7_75t_L g5667 ( 
.A(n_5638),
.B(n_5649),
.C(n_5650),
.D(n_5363),
.Y(n_5667)
);

AND2x2_ASAP7_75t_L g5668 ( 
.A(n_5641),
.B(n_5411),
.Y(n_5668)
);

AOI21xp5_ASAP7_75t_L g5669 ( 
.A1(n_5636),
.A2(n_5429),
.B(n_5426),
.Y(n_5669)
);

NAND2xp5_ASAP7_75t_L g5670 ( 
.A(n_5641),
.B(n_5413),
.Y(n_5670)
);

INVx1_ASAP7_75t_L g5671 ( 
.A(n_5636),
.Y(n_5671)
);

NAND4xp75_ASAP7_75t_L g5672 ( 
.A(n_5638),
.B(n_5361),
.C(n_5309),
.D(n_5313),
.Y(n_5672)
);

NAND3xp33_ASAP7_75t_L g5673 ( 
.A(n_5642),
.B(n_5317),
.C(n_5304),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_5636),
.Y(n_5674)
);

NAND2xp5_ASAP7_75t_L g5675 ( 
.A(n_5641),
.B(n_5398),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5636),
.Y(n_5676)
);

AOI22xp33_ASAP7_75t_SL g5677 ( 
.A1(n_5636),
.A2(n_5327),
.B1(n_5261),
.B2(n_5348),
.Y(n_5677)
);

AND2x2_ASAP7_75t_L g5678 ( 
.A(n_5641),
.B(n_5325),
.Y(n_5678)
);

NAND2xp5_ASAP7_75t_L g5679 ( 
.A(n_5641),
.B(n_5355),
.Y(n_5679)
);

AOI221x1_ASAP7_75t_L g5680 ( 
.A1(n_5644),
.A2(n_5353),
.B1(n_354),
.B2(n_352),
.C(n_353),
.Y(n_5680)
);

INVxp33_ASAP7_75t_L g5681 ( 
.A(n_5667),
.Y(n_5681)
);

NOR3xp33_ASAP7_75t_L g5682 ( 
.A(n_5664),
.B(n_354),
.C(n_356),
.Y(n_5682)
);

INVx2_ASAP7_75t_SL g5683 ( 
.A(n_5666),
.Y(n_5683)
);

AOI211xp5_ASAP7_75t_L g5684 ( 
.A1(n_5655),
.A2(n_359),
.B(n_356),
.C(n_357),
.Y(n_5684)
);

AND4x1_ASAP7_75t_L g5685 ( 
.A(n_5660),
.B(n_366),
.C(n_362),
.D(n_365),
.Y(n_5685)
);

AOI221xp5_ASAP7_75t_L g5686 ( 
.A1(n_5671),
.A2(n_5674),
.B1(n_5676),
.B2(n_5657),
.C(n_5656),
.Y(n_5686)
);

OAI211xp5_ASAP7_75t_SL g5687 ( 
.A1(n_5663),
.A2(n_369),
.B(n_367),
.C(n_368),
.Y(n_5687)
);

NOR2xp33_ASAP7_75t_L g5688 ( 
.A(n_5658),
.B(n_368),
.Y(n_5688)
);

NOR3xp33_ASAP7_75t_SL g5689 ( 
.A(n_5662),
.B(n_370),
.C(n_371),
.Y(n_5689)
);

OAI211xp5_ASAP7_75t_L g5690 ( 
.A1(n_5680),
.A2(n_373),
.B(n_371),
.C(n_372),
.Y(n_5690)
);

NAND4xp25_ASAP7_75t_L g5691 ( 
.A(n_5668),
.B(n_375),
.C(n_372),
.D(n_374),
.Y(n_5691)
);

NAND2xp5_ASAP7_75t_SL g5692 ( 
.A(n_5669),
.B(n_374),
.Y(n_5692)
);

OAI21xp5_ASAP7_75t_SL g5693 ( 
.A1(n_5670),
.A2(n_376),
.B(n_377),
.Y(n_5693)
);

NAND4xp75_ASAP7_75t_L g5694 ( 
.A(n_5665),
.B(n_378),
.C(n_376),
.D(n_377),
.Y(n_5694)
);

NAND4xp25_ASAP7_75t_SL g5695 ( 
.A(n_5661),
.B(n_382),
.C(n_378),
.D(n_379),
.Y(n_5695)
);

NOR2xp33_ASAP7_75t_L g5696 ( 
.A(n_5675),
.B(n_379),
.Y(n_5696)
);

NOR2xp67_ASAP7_75t_L g5697 ( 
.A(n_5673),
.B(n_382),
.Y(n_5697)
);

NAND2xp5_ASAP7_75t_L g5698 ( 
.A(n_5678),
.B(n_383),
.Y(n_5698)
);

AOI221xp5_ASAP7_75t_L g5699 ( 
.A1(n_5679),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.C(n_387),
.Y(n_5699)
);

NAND2xp5_ASAP7_75t_SL g5700 ( 
.A(n_5677),
.B(n_385),
.Y(n_5700)
);

NAND3xp33_ASAP7_75t_L g5701 ( 
.A(n_5659),
.B(n_387),
.C(n_388),
.Y(n_5701)
);

NOR4xp25_ASAP7_75t_L g5702 ( 
.A(n_5672),
.B(n_390),
.C(n_388),
.D(n_389),
.Y(n_5702)
);

AOI221xp5_ASAP7_75t_L g5703 ( 
.A1(n_5671),
.A2(n_390),
.B1(n_391),
.B2(n_393),
.C(n_394),
.Y(n_5703)
);

AND2x2_ASAP7_75t_L g5704 ( 
.A(n_5668),
.B(n_391),
.Y(n_5704)
);

NOR2xp33_ASAP7_75t_L g5705 ( 
.A(n_5658),
.B(n_395),
.Y(n_5705)
);

NAND2xp5_ASAP7_75t_L g5706 ( 
.A(n_5655),
.B(n_395),
.Y(n_5706)
);

NAND4xp25_ASAP7_75t_L g5707 ( 
.A(n_5660),
.B(n_398),
.C(n_396),
.D(n_397),
.Y(n_5707)
);

NOR2x1_ASAP7_75t_L g5708 ( 
.A(n_5662),
.B(n_396),
.Y(n_5708)
);

NAND3xp33_ASAP7_75t_SL g5709 ( 
.A(n_5685),
.B(n_399),
.C(n_401),
.Y(n_5709)
);

OAI321xp33_ASAP7_75t_L g5710 ( 
.A1(n_5707),
.A2(n_402),
.A3(n_403),
.B1(n_404),
.B2(n_405),
.C(n_407),
.Y(n_5710)
);

NAND4xp25_ASAP7_75t_L g5711 ( 
.A(n_5686),
.B(n_409),
.C(n_402),
.D(n_408),
.Y(n_5711)
);

NOR3x1_ASAP7_75t_L g5712 ( 
.A(n_5693),
.B(n_5701),
.C(n_5690),
.Y(n_5712)
);

AOI22xp5_ASAP7_75t_L g5713 ( 
.A1(n_5695),
.A2(n_413),
.B1(n_410),
.B2(n_411),
.Y(n_5713)
);

NOR2x1_ASAP7_75t_L g5714 ( 
.A(n_5694),
.B(n_413),
.Y(n_5714)
);

INVx2_ASAP7_75t_L g5715 ( 
.A(n_5704),
.Y(n_5715)
);

NAND5xp2_ASAP7_75t_L g5716 ( 
.A(n_5681),
.B(n_414),
.C(n_415),
.D(n_416),
.E(n_418),
.Y(n_5716)
);

O2A1O1Ixp33_ASAP7_75t_L g5717 ( 
.A1(n_5683),
.A2(n_420),
.B(n_418),
.C(n_419),
.Y(n_5717)
);

NAND4xp25_ASAP7_75t_L g5718 ( 
.A(n_5696),
.B(n_422),
.C(n_419),
.D(n_421),
.Y(n_5718)
);

INVx1_ASAP7_75t_SL g5719 ( 
.A(n_5706),
.Y(n_5719)
);

AOI21xp33_ASAP7_75t_SL g5720 ( 
.A1(n_5682),
.A2(n_422),
.B(n_423),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_5708),
.Y(n_5721)
);

AOI22xp5_ASAP7_75t_L g5722 ( 
.A1(n_5688),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_5722)
);

NOR3xp33_ASAP7_75t_L g5723 ( 
.A(n_5705),
.B(n_425),
.C(n_426),
.Y(n_5723)
);

AOI221xp5_ASAP7_75t_L g5724 ( 
.A1(n_5702),
.A2(n_426),
.B1(n_427),
.B2(n_428),
.C(n_429),
.Y(n_5724)
);

AOI211xp5_ASAP7_75t_L g5725 ( 
.A1(n_5687),
.A2(n_431),
.B(n_427),
.C(n_430),
.Y(n_5725)
);

AOI322xp5_ASAP7_75t_L g5726 ( 
.A1(n_5692),
.A2(n_430),
.A3(n_432),
.B1(n_433),
.B2(n_434),
.C1(n_435),
.C2(n_436),
.Y(n_5726)
);

AOI221xp5_ASAP7_75t_L g5727 ( 
.A1(n_5700),
.A2(n_434),
.B1(n_436),
.B2(n_437),
.C(n_438),
.Y(n_5727)
);

AOI221xp5_ASAP7_75t_L g5728 ( 
.A1(n_5698),
.A2(n_439),
.B1(n_440),
.B2(n_442),
.C(n_443),
.Y(n_5728)
);

NAND3xp33_ASAP7_75t_L g5729 ( 
.A(n_5689),
.B(n_439),
.C(n_440),
.Y(n_5729)
);

AO22x2_ASAP7_75t_L g5730 ( 
.A1(n_5684),
.A2(n_5691),
.B1(n_5697),
.B2(n_5699),
.Y(n_5730)
);

NAND4xp25_ASAP7_75t_SL g5731 ( 
.A(n_5703),
.B(n_442),
.C(n_443),
.D(n_444),
.Y(n_5731)
);

NOR4xp25_ASAP7_75t_L g5732 ( 
.A(n_5707),
.B(n_445),
.C(n_446),
.D(n_447),
.Y(n_5732)
);

AOI211x1_ASAP7_75t_L g5733 ( 
.A1(n_5685),
.A2(n_445),
.B(n_448),
.C(n_449),
.Y(n_5733)
);

AOI321xp33_ASAP7_75t_L g5734 ( 
.A1(n_5715),
.A2(n_448),
.A3(n_449),
.B1(n_450),
.B2(n_451),
.C(n_452),
.Y(n_5734)
);

CKINVDCx5p33_ASAP7_75t_R g5735 ( 
.A(n_5719),
.Y(n_5735)
);

INVxp67_ASAP7_75t_L g5736 ( 
.A(n_5716),
.Y(n_5736)
);

AOI21xp5_ASAP7_75t_L g5737 ( 
.A1(n_5709),
.A2(n_450),
.B(n_451),
.Y(n_5737)
);

OAI211xp5_ASAP7_75t_SL g5738 ( 
.A1(n_5714),
.A2(n_452),
.B(n_453),
.C(n_454),
.Y(n_5738)
);

INVx2_ASAP7_75t_SL g5739 ( 
.A(n_5721),
.Y(n_5739)
);

OAI211xp5_ASAP7_75t_L g5740 ( 
.A1(n_5727),
.A2(n_453),
.B(n_455),
.C(n_457),
.Y(n_5740)
);

OAI22xp5_ASAP7_75t_L g5741 ( 
.A1(n_5713),
.A2(n_457),
.B1(n_458),
.B2(n_459),
.Y(n_5741)
);

OAI22xp5_ASAP7_75t_L g5742 ( 
.A1(n_5729),
.A2(n_458),
.B1(n_460),
.B2(n_461),
.Y(n_5742)
);

AOI22xp5_ASAP7_75t_L g5743 ( 
.A1(n_5731),
.A2(n_462),
.B1(n_463),
.B2(n_464),
.Y(n_5743)
);

CKINVDCx16_ASAP7_75t_R g5744 ( 
.A(n_5732),
.Y(n_5744)
);

CKINVDCx6p67_ASAP7_75t_R g5745 ( 
.A(n_5733),
.Y(n_5745)
);

AOI31xp33_ASAP7_75t_L g5746 ( 
.A1(n_5725),
.A2(n_462),
.A3(n_467),
.B(n_468),
.Y(n_5746)
);

AOI221xp5_ASAP7_75t_L g5747 ( 
.A1(n_5724),
.A2(n_467),
.B1(n_468),
.B2(n_469),
.C(n_470),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_5717),
.Y(n_5748)
);

NOR2xp33_ASAP7_75t_L g5749 ( 
.A(n_5718),
.B(n_469),
.Y(n_5749)
);

NAND3xp33_ASAP7_75t_L g5750 ( 
.A(n_5723),
.B(n_471),
.C(n_472),
.Y(n_5750)
);

NAND3xp33_ASAP7_75t_L g5751 ( 
.A(n_5711),
.B(n_471),
.C(n_472),
.Y(n_5751)
);

INVx1_ASAP7_75t_SL g5752 ( 
.A(n_5722),
.Y(n_5752)
);

NOR2x1_ASAP7_75t_L g5753 ( 
.A(n_5738),
.B(n_5726),
.Y(n_5753)
);

OR2x2_ASAP7_75t_L g5754 ( 
.A(n_5744),
.B(n_5741),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_5745),
.Y(n_5755)
);

NOR2x1_ASAP7_75t_L g5756 ( 
.A(n_5750),
.B(n_5710),
.Y(n_5756)
);

NOR2x1_ASAP7_75t_L g5757 ( 
.A(n_5748),
.B(n_5720),
.Y(n_5757)
);

NOR2x1_ASAP7_75t_L g5758 ( 
.A(n_5751),
.B(n_5712),
.Y(n_5758)
);

INVx1_ASAP7_75t_L g5759 ( 
.A(n_5743),
.Y(n_5759)
);

OAI22xp33_ASAP7_75t_L g5760 ( 
.A1(n_5746),
.A2(n_5728),
.B1(n_5730),
.B2(n_476),
.Y(n_5760)
);

INVx2_ASAP7_75t_L g5761 ( 
.A(n_5739),
.Y(n_5761)
);

NOR2x1_ASAP7_75t_L g5762 ( 
.A(n_5742),
.B(n_5730),
.Y(n_5762)
);

XNOR2xp5_ASAP7_75t_L g5763 ( 
.A(n_5735),
.B(n_473),
.Y(n_5763)
);

OR2x2_ASAP7_75t_L g5764 ( 
.A(n_5736),
.B(n_474),
.Y(n_5764)
);

INVx2_ASAP7_75t_L g5765 ( 
.A(n_5752),
.Y(n_5765)
);

NOR2xp67_ASAP7_75t_L g5766 ( 
.A(n_5740),
.B(n_474),
.Y(n_5766)
);

NAND4xp75_ASAP7_75t_L g5767 ( 
.A(n_5737),
.B(n_476),
.C(n_477),
.D(n_479),
.Y(n_5767)
);

NOR3xp33_ASAP7_75t_L g5768 ( 
.A(n_5749),
.B(n_481),
.C(n_482),
.Y(n_5768)
);

NAND4xp25_ASAP7_75t_SL g5769 ( 
.A(n_5755),
.B(n_5747),
.C(n_5734),
.D(n_486),
.Y(n_5769)
);

NAND4xp25_ASAP7_75t_L g5770 ( 
.A(n_5753),
.B(n_5764),
.C(n_5758),
.D(n_5762),
.Y(n_5770)
);

OR5x1_ASAP7_75t_L g5771 ( 
.A(n_5757),
.B(n_5756),
.C(n_5760),
.D(n_5766),
.E(n_5754),
.Y(n_5771)
);

AOI22xp33_ASAP7_75t_L g5772 ( 
.A1(n_5761),
.A2(n_482),
.B1(n_485),
.B2(n_486),
.Y(n_5772)
);

OAI221xp5_ASAP7_75t_SL g5773 ( 
.A1(n_5765),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.C(n_490),
.Y(n_5773)
);

NOR2xp33_ASAP7_75t_L g5774 ( 
.A(n_5767),
.B(n_489),
.Y(n_5774)
);

NAND4xp75_ASAP7_75t_L g5775 ( 
.A(n_5759),
.B(n_491),
.C(n_492),
.D(n_493),
.Y(n_5775)
);

NOR5xp2_ASAP7_75t_L g5776 ( 
.A(n_5768),
.B(n_491),
.C(n_493),
.D(n_494),
.E(n_495),
.Y(n_5776)
);

HB1xp67_ASAP7_75t_L g5777 ( 
.A(n_5763),
.Y(n_5777)
);

NAND4xp25_ASAP7_75t_L g5778 ( 
.A(n_5755),
.B(n_494),
.C(n_495),
.D(n_497),
.Y(n_5778)
);

AND2x4_ASAP7_75t_L g5779 ( 
.A(n_5755),
.B(n_498),
.Y(n_5779)
);

NOR4xp75_ASAP7_75t_L g5780 ( 
.A(n_5767),
.B(n_499),
.C(n_500),
.D(n_501),
.Y(n_5780)
);

NAND3xp33_ASAP7_75t_SL g5781 ( 
.A(n_5755),
.B(n_499),
.C(n_500),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_5763),
.Y(n_5782)
);

NOR5xp2_ASAP7_75t_L g5783 ( 
.A(n_5755),
.B(n_502),
.C(n_504),
.D(n_507),
.E(n_508),
.Y(n_5783)
);

NAND5xp2_ASAP7_75t_L g5784 ( 
.A(n_5755),
.B(n_508),
.C(n_509),
.D(n_510),
.E(n_511),
.Y(n_5784)
);

NAND4xp25_ASAP7_75t_SL g5785 ( 
.A(n_5755),
.B(n_510),
.C(n_511),
.D(n_512),
.Y(n_5785)
);

NAND3xp33_ASAP7_75t_SL g5786 ( 
.A(n_5755),
.B(n_512),
.C(n_513),
.Y(n_5786)
);

AOI21xp5_ASAP7_75t_L g5787 ( 
.A1(n_5770),
.A2(n_513),
.B(n_515),
.Y(n_5787)
);

NAND2xp5_ASAP7_75t_L g5788 ( 
.A(n_5774),
.B(n_516),
.Y(n_5788)
);

AND2x4_ASAP7_75t_L g5789 ( 
.A(n_5780),
.B(n_516),
.Y(n_5789)
);

INVx2_ASAP7_75t_SL g5790 ( 
.A(n_5779),
.Y(n_5790)
);

HB1xp67_ASAP7_75t_L g5791 ( 
.A(n_5775),
.Y(n_5791)
);

BUFx2_ASAP7_75t_L g5792 ( 
.A(n_5779),
.Y(n_5792)
);

BUFx2_ASAP7_75t_L g5793 ( 
.A(n_5778),
.Y(n_5793)
);

INVx1_ASAP7_75t_SL g5794 ( 
.A(n_5771),
.Y(n_5794)
);

NOR2xp33_ASAP7_75t_R g5795 ( 
.A(n_5781),
.B(n_517),
.Y(n_5795)
);

AO221x1_ASAP7_75t_L g5796 ( 
.A1(n_5782),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.C(n_520),
.Y(n_5796)
);

HB1xp67_ASAP7_75t_L g5797 ( 
.A(n_5785),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_5786),
.Y(n_5798)
);

NAND2xp5_ASAP7_75t_L g5799 ( 
.A(n_5772),
.B(n_518),
.Y(n_5799)
);

INVx1_ASAP7_75t_L g5800 ( 
.A(n_5784),
.Y(n_5800)
);

OAI221xp5_ASAP7_75t_SL g5801 ( 
.A1(n_5794),
.A2(n_5777),
.B1(n_5769),
.B2(n_5776),
.C(n_5783),
.Y(n_5801)
);

HB1xp67_ASAP7_75t_L g5802 ( 
.A(n_5789),
.Y(n_5802)
);

INVx2_ASAP7_75t_SL g5803 ( 
.A(n_5796),
.Y(n_5803)
);

AOI221xp5_ASAP7_75t_L g5804 ( 
.A1(n_5787),
.A2(n_5773),
.B1(n_521),
.B2(n_522),
.C(n_523),
.Y(n_5804)
);

AOI322xp5_ASAP7_75t_L g5805 ( 
.A1(n_5789),
.A2(n_520),
.A3(n_521),
.B1(n_523),
.B2(n_524),
.C1(n_525),
.C2(n_526),
.Y(n_5805)
);

AOI22x1_ASAP7_75t_L g5806 ( 
.A1(n_5792),
.A2(n_524),
.B1(n_527),
.B2(n_528),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_5788),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_5802),
.Y(n_5808)
);

AOI22xp5_ASAP7_75t_L g5809 ( 
.A1(n_5803),
.A2(n_5800),
.B1(n_5798),
.B2(n_5790),
.Y(n_5809)
);

OAI22xp5_ASAP7_75t_L g5810 ( 
.A1(n_5801),
.A2(n_5799),
.B1(n_5797),
.B2(n_5791),
.Y(n_5810)
);

AOI22xp5_ASAP7_75t_L g5811 ( 
.A1(n_5804),
.A2(n_5793),
.B1(n_5795),
.B2(n_530),
.Y(n_5811)
);

AO22x2_ASAP7_75t_L g5812 ( 
.A1(n_5807),
.A2(n_527),
.B1(n_529),
.B2(n_531),
.Y(n_5812)
);

INVx1_ASAP7_75t_L g5813 ( 
.A(n_5806),
.Y(n_5813)
);

AOI22x1_ASAP7_75t_L g5814 ( 
.A1(n_5805),
.A2(n_531),
.B1(n_532),
.B2(n_533),
.Y(n_5814)
);

OAI322xp33_ASAP7_75t_L g5815 ( 
.A1(n_5809),
.A2(n_532),
.A3(n_536),
.B1(n_538),
.B2(n_539),
.C1(n_540),
.C2(n_541),
.Y(n_5815)
);

INVx2_ASAP7_75t_L g5816 ( 
.A(n_5812),
.Y(n_5816)
);

NAND5xp2_ASAP7_75t_L g5817 ( 
.A(n_5808),
.B(n_539),
.C(n_542),
.D(n_543),
.E(n_544),
.Y(n_5817)
);

XNOR2xp5_ASAP7_75t_L g5818 ( 
.A(n_5814),
.B(n_544),
.Y(n_5818)
);

OAI22xp5_ASAP7_75t_SL g5819 ( 
.A1(n_5813),
.A2(n_5811),
.B1(n_5810),
.B2(n_547),
.Y(n_5819)
);

OAI22xp5_ASAP7_75t_L g5820 ( 
.A1(n_5809),
.A2(n_545),
.B1(n_546),
.B2(n_547),
.Y(n_5820)
);

XNOR2xp5_ASAP7_75t_L g5821 ( 
.A(n_5818),
.B(n_545),
.Y(n_5821)
);

OAI22xp5_ASAP7_75t_SL g5822 ( 
.A1(n_5819),
.A2(n_546),
.B1(n_548),
.B2(n_549),
.Y(n_5822)
);

AOI31xp33_ASAP7_75t_L g5823 ( 
.A1(n_5816),
.A2(n_549),
.A3(n_550),
.B(n_552),
.Y(n_5823)
);

INVxp67_ASAP7_75t_SL g5824 ( 
.A(n_5820),
.Y(n_5824)
);

AND2x2_ASAP7_75t_L g5825 ( 
.A(n_5817),
.B(n_555),
.Y(n_5825)
);

AOI21xp33_ASAP7_75t_L g5826 ( 
.A1(n_5821),
.A2(n_5815),
.B(n_556),
.Y(n_5826)
);

OAI22xp5_ASAP7_75t_L g5827 ( 
.A1(n_5822),
.A2(n_5824),
.B1(n_5825),
.B2(n_5823),
.Y(n_5827)
);

INVx1_ASAP7_75t_L g5828 ( 
.A(n_5825),
.Y(n_5828)
);

OAI22xp5_ASAP7_75t_L g5829 ( 
.A1(n_5821),
.A2(n_555),
.B1(n_557),
.B2(n_560),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_5829),
.Y(n_5830)
);

AOI22xp33_ASAP7_75t_L g5831 ( 
.A1(n_5828),
.A2(n_557),
.B1(n_561),
.B2(n_562),
.Y(n_5831)
);

AOI22xp5_ASAP7_75t_L g5832 ( 
.A1(n_5827),
.A2(n_561),
.B1(n_562),
.B2(n_563),
.Y(n_5832)
);

OAI21xp33_ASAP7_75t_L g5833 ( 
.A1(n_5826),
.A2(n_563),
.B(n_565),
.Y(n_5833)
);

OAI21xp5_ASAP7_75t_L g5834 ( 
.A1(n_5827),
.A2(n_567),
.B(n_568),
.Y(n_5834)
);

OAI22xp5_ASAP7_75t_L g5835 ( 
.A1(n_5833),
.A2(n_570),
.B1(n_572),
.B2(n_573),
.Y(n_5835)
);

OR2x2_ASAP7_75t_L g5836 ( 
.A(n_5830),
.B(n_5834),
.Y(n_5836)
);

AOI22xp33_ASAP7_75t_L g5837 ( 
.A1(n_5831),
.A2(n_574),
.B1(n_575),
.B2(n_576),
.Y(n_5837)
);

AOI21xp5_ASAP7_75t_L g5838 ( 
.A1(n_5832),
.A2(n_1759),
.B(n_1757),
.Y(n_5838)
);

NAND2xp5_ASAP7_75t_L g5839 ( 
.A(n_5833),
.B(n_575),
.Y(n_5839)
);

NAND2xp5_ASAP7_75t_L g5840 ( 
.A(n_5833),
.B(n_576),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_5833),
.Y(n_5841)
);

OR2x6_ASAP7_75t_L g5842 ( 
.A(n_5830),
.B(n_577),
.Y(n_5842)
);

AO22x2_ASAP7_75t_L g5843 ( 
.A1(n_5830),
.A2(n_579),
.B1(n_580),
.B2(n_581),
.Y(n_5843)
);

AOI21xp5_ASAP7_75t_L g5844 ( 
.A1(n_5830),
.A2(n_1759),
.B(n_1757),
.Y(n_5844)
);

AOI22xp5_ASAP7_75t_L g5845 ( 
.A1(n_5835),
.A2(n_5840),
.B1(n_5839),
.B2(n_5837),
.Y(n_5845)
);

OAI22xp5_ASAP7_75t_L g5846 ( 
.A1(n_5836),
.A2(n_581),
.B1(n_582),
.B2(n_583),
.Y(n_5846)
);

AO22x2_ASAP7_75t_L g5847 ( 
.A1(n_5841),
.A2(n_583),
.B1(n_584),
.B2(n_586),
.Y(n_5847)
);

AOI22xp5_ASAP7_75t_L g5848 ( 
.A1(n_5842),
.A2(n_586),
.B1(n_588),
.B2(n_589),
.Y(n_5848)
);

AO22x1_ASAP7_75t_L g5849 ( 
.A1(n_5844),
.A2(n_588),
.B1(n_590),
.B2(n_591),
.Y(n_5849)
);

AOI22xp5_ASAP7_75t_SL g5850 ( 
.A1(n_5838),
.A2(n_593),
.B1(n_594),
.B2(n_595),
.Y(n_5850)
);

OAI22xp33_ASAP7_75t_L g5851 ( 
.A1(n_5843),
.A2(n_593),
.B1(n_594),
.B2(n_598),
.Y(n_5851)
);

AOI22xp5_ASAP7_75t_L g5852 ( 
.A1(n_5835),
.A2(n_598),
.B1(n_599),
.B2(n_600),
.Y(n_5852)
);

OAI22xp5_ASAP7_75t_L g5853 ( 
.A1(n_5837),
.A2(n_599),
.B1(n_600),
.B2(n_601),
.Y(n_5853)
);

AO22x2_ASAP7_75t_L g5854 ( 
.A1(n_5841),
.A2(n_602),
.B1(n_603),
.B2(n_605),
.Y(n_5854)
);

INVx1_ASAP7_75t_L g5855 ( 
.A(n_5845),
.Y(n_5855)
);

NOR2xp33_ASAP7_75t_L g5856 ( 
.A(n_5851),
.B(n_602),
.Y(n_5856)
);

AO21x2_ASAP7_75t_L g5857 ( 
.A1(n_5852),
.A2(n_606),
.B(n_607),
.Y(n_5857)
);

NAND3xp33_ASAP7_75t_L g5858 ( 
.A(n_5853),
.B(n_1719),
.C(n_1757),
.Y(n_5858)
);

OAI21xp5_ASAP7_75t_L g5859 ( 
.A1(n_5850),
.A2(n_608),
.B(n_610),
.Y(n_5859)
);

NAND2xp5_ASAP7_75t_L g5860 ( 
.A(n_5849),
.B(n_608),
.Y(n_5860)
);

AOI21xp5_ASAP7_75t_L g5861 ( 
.A1(n_5846),
.A2(n_1719),
.B(n_1757),
.Y(n_5861)
);

OAI21xp5_ASAP7_75t_L g5862 ( 
.A1(n_5848),
.A2(n_612),
.B(n_613),
.Y(n_5862)
);

INVx1_ASAP7_75t_L g5863 ( 
.A(n_5860),
.Y(n_5863)
);

OAI22xp33_ASAP7_75t_L g5864 ( 
.A1(n_5855),
.A2(n_5854),
.B1(n_5847),
.B2(n_615),
.Y(n_5864)
);

INVx1_ASAP7_75t_L g5865 ( 
.A(n_5856),
.Y(n_5865)
);

AOI22xp5_ASAP7_75t_L g5866 ( 
.A1(n_5857),
.A2(n_613),
.B1(n_614),
.B2(n_616),
.Y(n_5866)
);

AOI221xp5_ASAP7_75t_L g5867 ( 
.A1(n_5864),
.A2(n_5859),
.B1(n_5858),
.B2(n_5861),
.C(n_5862),
.Y(n_5867)
);

AOI221xp5_ASAP7_75t_L g5868 ( 
.A1(n_5867),
.A2(n_5865),
.B1(n_5863),
.B2(n_5866),
.C(n_622),
.Y(n_5868)
);

AOI211xp5_ASAP7_75t_L g5869 ( 
.A1(n_5868),
.A2(n_617),
.B(n_618),
.C(n_619),
.Y(n_5869)
);


endmodule