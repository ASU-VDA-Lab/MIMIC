module fake_ariane_188_n_2369 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2369);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2369;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2334;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_2332;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_347;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1856;
wire n_1733;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_253;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_308;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2275;
wire n_2183;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_L g226 ( 
.A(n_20),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_96),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_65),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_97),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_9),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_220),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_87),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_82),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_139),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_142),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_29),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_117),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_84),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_122),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_24),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_48),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_1),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_55),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_127),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_33),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_159),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_108),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_3),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_156),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_123),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_48),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_34),
.Y(n_255)
);

BUFx8_ASAP7_75t_SL g256 ( 
.A(n_216),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_109),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_67),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_99),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_188),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_60),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_124),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_7),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_205),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_38),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_114),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_145),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_177),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_99),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_27),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_15),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_154),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_126),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_185),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_37),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_42),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_40),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_21),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_74),
.Y(n_279)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_9),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_36),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_42),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_74),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_85),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_182),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_47),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_79),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_155),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_8),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_217),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_81),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_134),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_191),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_137),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_22),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_208),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_20),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_173),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_70),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_160),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_104),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_176),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_43),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_102),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_31),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_121),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_63),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_206),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_80),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_2),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_161),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_16),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_65),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_211),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_204),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_158),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_90),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_87),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_63),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_175),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_138),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_62),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_183),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_130),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_94),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_71),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_162),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_95),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_38),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_171),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_33),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_24),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_166),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_153),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_41),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_152),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_72),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_143),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_93),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_172),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_221),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_78),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_75),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_7),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_225),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_43),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_219),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_120),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_41),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_40),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_189),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_0),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_32),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_11),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_170),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_200),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_196),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_190),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_163),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_39),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_144),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_207),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_23),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_184),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_0),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_98),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_97),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_222),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_113),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_164),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_103),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_115),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_80),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_150),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_165),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_29),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_91),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_12),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_13),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_202),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_37),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_168),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_27),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_180),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_77),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_75),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_49),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_140),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_53),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_101),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_44),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_50),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_100),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_19),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_223),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_194),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_30),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_1),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_136),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_58),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_135),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_209),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_25),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_195),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_8),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_111),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_82),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_15),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_129),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_3),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_102),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_34),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_131),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_10),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_12),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_62),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_72),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_70),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_56),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_90),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_224),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_125),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_28),
.Y(n_423)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_45),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_67),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_112),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_35),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_21),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_45),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_64),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_36),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_23),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_83),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_201),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_167),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_88),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_203),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_116),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_14),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_212),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_17),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_96),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_32),
.Y(n_443)
);

BUFx8_ASAP7_75t_SL g444 ( 
.A(n_28),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_66),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_235),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_235),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_237),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_237),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_227),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_R g451 ( 
.A(n_345),
.B(n_105),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_246),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_246),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_277),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_227),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_444),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_444),
.Y(n_457)
);

INVxp33_ASAP7_75t_SL g458 ( 
.A(n_287),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_274),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_256),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_285),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_262),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_300),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_285),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_290),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_290),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_292),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_314),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_336),
.B(n_2),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_336),
.B(n_4),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_292),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_338),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_287),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_256),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_296),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_240),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_243),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_296),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_302),
.B(n_4),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_301),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_301),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_311),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_248),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_302),
.Y(n_484)
);

INVx4_ASAP7_75t_R g485 ( 
.A(n_264),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_311),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_316),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_316),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_320),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_242),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_258),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_320),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_371),
.B(n_5),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_245),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_327),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_327),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_297),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_251),
.Y(n_498)
);

INVxp33_ASAP7_75t_SL g499 ( 
.A(n_414),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_326),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_371),
.B(n_401),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_330),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_360),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_330),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_340),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_340),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_414),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_351),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_244),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_351),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_355),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_355),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_262),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_254),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_401),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_255),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_362),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_353),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_353),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_259),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_261),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_362),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_265),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_269),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_369),
.B(n_5),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_353),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_408),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_277),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_369),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g530 ( 
.A(n_226),
.B(n_6),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_270),
.Y(n_531)
);

INVxp33_ASAP7_75t_L g532 ( 
.A(n_244),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_380),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_380),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_442),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_384),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_271),
.Y(n_537)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_353),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_384),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_R g540 ( 
.A(n_345),
.B(n_106),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_275),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_276),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_399),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_279),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_282),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_399),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_284),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_289),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_291),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_295),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_402),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_299),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_306),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_280),
.B(n_6),
.Y(n_554)
);

INVxp33_ASAP7_75t_SL g555 ( 
.A(n_352),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_280),
.B(n_10),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_307),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_352),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_402),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_406),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_406),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_226),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_306),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_312),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_L g565 ( 
.A(n_226),
.B(n_11),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_483),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_562),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_SL g568 ( 
.A(n_501),
.B(n_424),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_446),
.B(n_277),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_562),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_474),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_483),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_477),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_460),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_457),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_491),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_446),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_455),
.B(n_423),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_447),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_447),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_454),
.B(n_423),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_448),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_459),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_448),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_528),
.B(n_250),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_463),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_R g587 ( 
.A(n_476),
.B(n_231),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_449),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_497),
.A2(n_424),
.B1(n_443),
.B2(n_303),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_458),
.A2(n_303),
.B1(n_309),
.B2(n_228),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_484),
.B(n_443),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_449),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_452),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_468),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_452),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_472),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_490),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_500),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_479),
.B(n_250),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_453),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_R g601 ( 
.A(n_494),
.B(n_313),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_453),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_461),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_461),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_464),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_464),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_465),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_499),
.A2(n_309),
.B1(n_342),
.B2(n_228),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_509),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_465),
.B(n_332),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_466),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_498),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_514),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_503),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_558),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_516),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_466),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_527),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_467),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_467),
.B(n_372),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_471),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_471),
.B(n_332),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_520),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_R g624 ( 
.A(n_521),
.B(n_234),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_523),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_475),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_475),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_478),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_484),
.B(n_332),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_478),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_R g631 ( 
.A(n_524),
.B(n_317),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_531),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_537),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_456),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_480),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_473),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_480),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_541),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_542),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_481),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_515),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_515),
.B(n_363),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_481),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_482),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_544),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_482),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_535),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_493),
.B(n_372),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_486),
.Y(n_649)
);

NOR2x1_ASAP7_75t_L g650 ( 
.A(n_486),
.B(n_487),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_545),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_R g652 ( 
.A(n_547),
.B(n_319),
.Y(n_652)
);

AND2x6_ASAP7_75t_L g653 ( 
.A(n_487),
.B(n_236),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_507),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_548),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_488),
.Y(n_656)
);

NAND2x1p5_ASAP7_75t_L g657 ( 
.A(n_488),
.B(n_264),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_489),
.B(n_321),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_549),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_450),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_577),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_569),
.B(n_489),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_566),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_569),
.B(n_492),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_583),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_635),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_577),
.Y(n_667)
);

INVx4_ASAP7_75t_SL g668 ( 
.A(n_653),
.Y(n_668)
);

OAI22xp33_ASAP7_75t_L g669 ( 
.A1(n_590),
.A2(n_462),
.B1(n_513),
.B2(n_532),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_569),
.B(n_492),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_657),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_566),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_579),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_569),
.B(n_495),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_572),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_579),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_599),
.B(n_518),
.Y(n_677)
);

AND2x2_ASAP7_75t_SL g678 ( 
.A(n_648),
.B(n_469),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_599),
.B(n_519),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_648),
.B(n_495),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_573),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_566),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_572),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_580),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_580),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_572),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_657),
.B(n_550),
.Y(n_687)
);

INVx8_ASAP7_75t_L g688 ( 
.A(n_610),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_576),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_584),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_584),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_566),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_657),
.B(n_552),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_602),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_641),
.B(n_526),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_641),
.B(n_538),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_649),
.B(n_557),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_635),
.Y(n_698)
);

OR2x6_ASAP7_75t_L g699 ( 
.A(n_657),
.B(n_470),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_566),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_658),
.B(n_496),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_592),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_598),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_610),
.B(n_496),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_602),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_566),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_635),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_592),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_582),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_614),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_602),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_582),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_568),
.A2(n_581),
.B1(n_585),
.B2(n_601),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_SL g714 ( 
.A(n_612),
.B(n_553),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_582),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_588),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_593),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_593),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_588),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_600),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_589),
.B(n_530),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_602),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_649),
.B(n_564),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_600),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_586),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_658),
.B(n_649),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_634),
.Y(n_727)
);

INVx5_ASAP7_75t_L g728 ( 
.A(n_653),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_588),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_603),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_618),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_610),
.B(n_502),
.Y(n_732)
);

OAI21xp33_ASAP7_75t_L g733 ( 
.A1(n_620),
.A2(n_556),
.B(n_554),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_649),
.B(n_451),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_595),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_637),
.B(n_502),
.Y(n_736)
);

AND2x6_ASAP7_75t_L g737 ( 
.A(n_650),
.B(n_504),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_595),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_603),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_637),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_637),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_637),
.B(n_540),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_605),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_605),
.Y(n_744)
);

INVx4_ASAP7_75t_SL g745 ( 
.A(n_653),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_610),
.B(n_622),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_595),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_651),
.B(n_555),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_634),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_646),
.B(n_504),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_604),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_650),
.B(n_505),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_651),
.B(n_563),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_646),
.B(n_606),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_646),
.B(n_505),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_606),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_646),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_604),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_607),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_636),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_622),
.B(n_506),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_607),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_647),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_604),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_617),
.Y(n_765)
);

OR2x6_ASAP7_75t_L g766 ( 
.A(n_589),
.B(n_565),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_622),
.B(n_506),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_617),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_619),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_619),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_621),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_587),
.B(n_525),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_621),
.B(n_508),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_620),
.B(n_508),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_611),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_626),
.B(n_510),
.Y(n_776)
);

BUFx10_ASAP7_75t_L g777 ( 
.A(n_616),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_594),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_626),
.Y(n_779)
);

INVx5_ASAP7_75t_L g780 ( 
.A(n_653),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_611),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_611),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_627),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_627),
.B(n_510),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_630),
.B(n_643),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_636),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_628),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_624),
.B(n_321),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_630),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_643),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_SL g791 ( 
.A1(n_578),
.A2(n_386),
.B1(n_485),
.B2(n_342),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_644),
.B(n_396),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_644),
.B(n_511),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_628),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_656),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_656),
.B(n_511),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_622),
.B(n_512),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_628),
.B(n_512),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_640),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_640),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_640),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_596),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_631),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_623),
.B(n_396),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_567),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_581),
.B(n_629),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_629),
.B(n_642),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_653),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_642),
.B(n_517),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_660),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_567),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_654),
.B(n_517),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_570),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_570),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_638),
.B(n_409),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_654),
.B(n_522),
.Y(n_816)
);

AND2x2_ASAP7_75t_SL g817 ( 
.A(n_597),
.B(n_229),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_591),
.B(n_522),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_591),
.B(n_529),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_653),
.Y(n_820)
);

NOR2x1p5_ASAP7_75t_L g821 ( 
.A(n_639),
.B(n_363),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_SL g822 ( 
.A1(n_817),
.A2(n_578),
.B1(n_659),
.B2(n_613),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_678),
.A2(n_608),
.B1(n_590),
.B2(n_609),
.Y(n_823)
);

INVxp67_ASAP7_75t_SL g824 ( 
.A(n_666),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_701),
.B(n_774),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_733),
.A2(n_233),
.B(n_281),
.C(n_229),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_726),
.A2(n_533),
.B(n_529),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_701),
.B(n_645),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_817),
.B(n_803),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_677),
.B(n_597),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_774),
.B(n_613),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_675),
.Y(n_832)
);

NAND3xp33_ASAP7_75t_L g833 ( 
.A(n_678),
.B(n_652),
.C(n_534),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_679),
.B(n_625),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_680),
.B(n_625),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_746),
.B(n_632),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_721),
.A2(n_608),
.B1(n_615),
.B2(n_609),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_752),
.B(n_632),
.Y(n_838)
);

INVx8_ASAP7_75t_L g839 ( 
.A(n_737),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_675),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_721),
.A2(n_615),
.B1(n_534),
.B2(n_536),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_752),
.B(n_633),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_705),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_688),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_688),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_694),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_705),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_697),
.B(n_633),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_723),
.B(n_655),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_683),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_683),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_748),
.B(n_655),
.Y(n_852)
);

OAI22xp33_ASAP7_75t_L g853 ( 
.A1(n_713),
.A2(n_699),
.B1(n_786),
.B2(n_760),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_746),
.B(n_659),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_741),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_695),
.B(n_574),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_696),
.B(n_575),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_712),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_760),
.B(n_575),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_662),
.B(n_533),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_786),
.B(n_386),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_741),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_709),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_662),
.B(n_536),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_709),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_797),
.A2(n_233),
.B(n_281),
.C(n_229),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_687),
.B(n_571),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_671),
.B(n_539),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_694),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_686),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_746),
.B(n_662),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_716),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_671),
.B(n_386),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_664),
.B(n_386),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_664),
.B(n_539),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_686),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_694),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_664),
.B(n_543),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_716),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_670),
.B(n_543),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_670),
.B(n_546),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_719),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_688),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_737),
.A2(n_699),
.B1(n_674),
.B2(n_670),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_688),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_719),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_749),
.B(n_546),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_666),
.Y(n_888)
);

AO22x1_ASAP7_75t_L g889 ( 
.A1(n_737),
.A2(n_559),
.B1(n_560),
.B2(n_551),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_729),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_674),
.B(n_551),
.Y(n_891)
);

OAI221xp5_ASAP7_75t_L g892 ( 
.A1(n_806),
.A2(n_283),
.B1(n_415),
.B2(n_416),
.C(n_392),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_674),
.B(n_559),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_729),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_704),
.B(n_560),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_704),
.B(n_561),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_704),
.B(n_561),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_738),
.Y(n_898)
);

AND2x6_ASAP7_75t_SL g899 ( 
.A(n_753),
.B(n_230),
.Y(n_899)
);

AND2x2_ASAP7_75t_SL g900 ( 
.A(n_740),
.B(n_233),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_732),
.B(n_409),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_740),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_732),
.B(n_440),
.Y(n_903)
);

NAND2xp33_ASAP7_75t_L g904 ( 
.A(n_737),
.B(n_653),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_732),
.B(n_440),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_665),
.Y(n_906)
);

BUFx12f_ASAP7_75t_L g907 ( 
.A(n_777),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_721),
.A2(n_333),
.B1(n_413),
.B2(n_306),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_687),
.B(n_693),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_761),
.B(n_281),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_737),
.A2(n_322),
.B1(n_329),
.B2(n_328),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_738),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_SL g913 ( 
.A(n_669),
.B(n_306),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_698),
.Y(n_914)
);

OAI22x1_ASAP7_75t_SL g915 ( 
.A1(n_810),
.A2(n_725),
.B1(n_778),
.B2(n_665),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_740),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_761),
.B(n_310),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_747),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_747),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_812),
.A2(n_349),
.B(n_367),
.C(n_310),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_751),
.Y(n_921)
);

NOR2xp67_ASAP7_75t_L g922 ( 
.A(n_808),
.B(n_107),
.Y(n_922)
);

INVx5_ASAP7_75t_L g923 ( 
.A(n_808),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_698),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_761),
.B(n_310),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_767),
.B(n_807),
.Y(n_926)
);

O2A1O1Ixp5_ASAP7_75t_L g927 ( 
.A1(n_742),
.A2(n_367),
.B(n_393),
.C(n_349),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_711),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_737),
.A2(n_337),
.B1(n_343),
.B2(n_335),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_767),
.B(n_349),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_767),
.B(n_230),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_707),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_762),
.B(n_367),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_785),
.A2(n_393),
.B(n_238),
.C(n_263),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_751),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_693),
.B(n_346),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_749),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_762),
.B(n_393),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_816),
.B(n_232),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_758),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_707),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_814),
.B(n_363),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_776),
.B(n_394),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_758),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_764),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_727),
.B(n_232),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_764),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_796),
.B(n_809),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_804),
.B(n_354),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_775),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_699),
.A2(n_365),
.B1(n_366),
.B2(n_441),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_775),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_721),
.A2(n_766),
.B1(n_699),
.B2(n_804),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_821),
.B(n_238),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_815),
.B(n_376),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_781),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_818),
.B(n_263),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_725),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_722),
.B(n_394),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_815),
.B(n_772),
.Y(n_960)
);

NAND2x1p5_ASAP7_75t_L g961 ( 
.A(n_820),
.B(n_236),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_781),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_819),
.B(n_278),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_722),
.B(n_394),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_722),
.B(n_278),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_794),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_711),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_757),
.B(n_283),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_681),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_757),
.B(n_286),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_794),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_801),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_757),
.B(n_286),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_799),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_712),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_801),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_801),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_712),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_712),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_777),
.B(n_377),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_R g981 ( 
.A(n_778),
.B(n_239),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_712),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_777),
.B(n_378),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_715),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_661),
.B(n_304),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_715),
.Y(n_986)
);

BUFx12f_ASAP7_75t_L g987 ( 
.A(n_766),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_715),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_715),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_766),
.A2(n_413),
.B1(n_437),
.B2(n_333),
.Y(n_990)
);

BUFx12f_ASAP7_75t_L g991 ( 
.A(n_766),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_800),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_667),
.B(n_304),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_673),
.A2(n_383),
.B(n_445),
.C(n_389),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_772),
.B(n_379),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_SL g996 ( 
.A1(n_810),
.A2(n_417),
.B1(n_385),
.B2(n_439),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_843),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_907),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_836),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_825),
.B(n_802),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_843),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_844),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_832),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_835),
.B(n_788),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_832),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_852),
.B(n_714),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_840),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_836),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_900),
.A2(n_792),
.B1(n_788),
.B2(n_742),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_907),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_840),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_830),
.B(n_792),
.Y(n_1012)
);

AND2x6_ASAP7_75t_SL g1013 ( 
.A(n_834),
.B(n_318),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_847),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_847),
.Y(n_1015)
);

INVx5_ASAP7_75t_L g1016 ( 
.A(n_923),
.Y(n_1016)
);

BUFx4f_ASAP7_75t_L g1017 ( 
.A(n_839),
.Y(n_1017)
);

NOR3xp33_ASAP7_75t_SL g1018 ( 
.A(n_906),
.B(n_387),
.C(n_381),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_848),
.B(n_676),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_R g1020 ( 
.A(n_906),
.B(n_689),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_900),
.B(n_734),
.Y(n_1021)
);

BUFx10_ASAP7_75t_L g1022 ( 
.A(n_958),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_850),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_937),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_855),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_855),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_900),
.B(n_734),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_845),
.Y(n_1028)
);

CKINVDCx8_ASAP7_75t_R g1029 ( 
.A(n_958),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_850),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_844),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_849),
.B(n_684),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_851),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_871),
.B(n_703),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_845),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_844),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_SL g1037 ( 
.A(n_856),
.B(n_397),
.C(n_391),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_851),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_870),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_926),
.A2(n_754),
.B1(n_690),
.B2(n_691),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_870),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_875),
.B(n_685),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_845),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_836),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_948),
.A2(n_708),
.B(n_702),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_969),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_862),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_853),
.A2(n_833),
.B1(n_884),
.B2(n_960),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_828),
.B(n_731),
.Y(n_1049)
);

AND2x6_ASAP7_75t_SL g1050 ( 
.A(n_859),
.B(n_318),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_915),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_R g1052 ( 
.A(n_831),
.B(n_689),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_885),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_875),
.B(n_717),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_876),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_862),
.Y(n_1056)
);

AND2x6_ASAP7_75t_L g1057 ( 
.A(n_885),
.B(n_715),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_885),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_895),
.B(n_718),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_863),
.Y(n_1060)
);

INVx5_ASAP7_75t_L g1061 ( 
.A(n_923),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_923),
.A2(n_724),
.B(n_720),
.Y(n_1062)
);

NOR3xp33_ASAP7_75t_SL g1063 ( 
.A(n_980),
.B(n_400),
.C(n_398),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_844),
.B(n_668),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_895),
.B(n_897),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_876),
.Y(n_1066)
);

INVx3_ASAP7_75t_SL g1067 ( 
.A(n_836),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_854),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_863),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_839),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_854),
.B(n_791),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_SL g1072 ( 
.A(n_983),
.B(n_405),
.C(n_403),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_897),
.B(n_730),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_897),
.B(n_739),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_865),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_SL g1076 ( 
.A(n_996),
.B(n_410),
.C(n_407),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_839),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_839),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_871),
.B(n_763),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_879),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_SL g1081 ( 
.A(n_996),
.B(n_412),
.C(n_411),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_865),
.Y(n_1082)
);

BUFx4f_ASAP7_75t_L g1083 ( 
.A(n_839),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_871),
.B(n_743),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_823),
.A2(n_805),
.B1(n_813),
.B2(n_811),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_879),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_897),
.B(n_744),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_872),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_860),
.B(n_756),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_838),
.B(n_710),
.Y(n_1090)
);

NOR3xp33_ASAP7_75t_SL g1091 ( 
.A(n_857),
.B(n_427),
.C(n_418),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_886),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_871),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_872),
.Y(n_1094)
);

AND3x1_ASAP7_75t_L g1095 ( 
.A(n_913),
.B(n_331),
.C(n_325),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_SL g1096 ( 
.A(n_951),
.B(n_430),
.C(n_429),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_915),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_SL g1098 ( 
.A(n_994),
.B(n_432),
.C(n_431),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_854),
.B(n_759),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_864),
.B(n_765),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_854),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_878),
.B(n_768),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_880),
.B(n_769),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_881),
.B(n_770),
.Y(n_1104)
);

BUFx12f_ASAP7_75t_SL g1105 ( 
.A(n_954),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_887),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_858),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_888),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_833),
.A2(n_790),
.B1(n_783),
.B2(n_771),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_888),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_887),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_891),
.B(n_779),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_893),
.B(n_789),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_931),
.B(n_795),
.Y(n_1114)
);

AND3x1_ASAP7_75t_L g1115 ( 
.A(n_913),
.B(n_331),
.C(n_325),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_981),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_883),
.B(n_710),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_858),
.Y(n_1118)
);

NAND2x2_ASAP7_75t_L g1119 ( 
.A(n_946),
.B(n_842),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_882),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_882),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_883),
.B(n_668),
.Y(n_1122)
);

INVxp67_ASAP7_75t_L g1123 ( 
.A(n_946),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_979),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_884),
.B(n_668),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_858),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_896),
.B(n_773),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_886),
.Y(n_1128)
);

NOR3xp33_ASAP7_75t_SL g1129 ( 
.A(n_867),
.B(n_436),
.C(n_344),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_979),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_931),
.B(n_805),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_979),
.Y(n_1132)
);

AND3x2_ASAP7_75t_SL g1133 ( 
.A(n_899),
.B(n_700),
.C(n_692),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_899),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_901),
.Y(n_1135)
);

AND2x6_ASAP7_75t_L g1136 ( 
.A(n_846),
.B(n_735),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_923),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_890),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_923),
.A2(n_750),
.B(n_736),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_939),
.B(n_784),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_890),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_894),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_898),
.Y(n_1143)
);

OR2x6_ASAP7_75t_L g1144 ( 
.A(n_987),
.B(n_991),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_987),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_898),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_939),
.B(n_793),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_923),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_903),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_894),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_957),
.B(n_755),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_957),
.B(n_798),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_912),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_888),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_950),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_963),
.B(n_735),
.Y(n_1156)
);

NOR3xp33_ASAP7_75t_SL g1157 ( 
.A(n_936),
.B(n_344),
.C(n_339),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_858),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_914),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_912),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_991),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_858),
.Y(n_1162)
);

BUFx12f_ASAP7_75t_L g1163 ( 
.A(n_954),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_822),
.B(n_735),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_829),
.A2(n_787),
.B1(n_782),
.B2(n_735),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_837),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_918),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_846),
.A2(n_735),
.B1(n_782),
.B2(n_787),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_918),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_919),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_967),
.Y(n_1171)
);

INVx6_ASAP7_75t_L g1172 ( 
.A(n_914),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_846),
.Y(n_1173)
);

BUFx10_ASAP7_75t_L g1174 ( 
.A(n_995),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_889),
.B(n_808),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_911),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_963),
.B(n_905),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_953),
.B(n_782),
.Y(n_1178)
);

AND3x2_ASAP7_75t_SL g1179 ( 
.A(n_889),
.B(n_700),
.C(n_692),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_914),
.Y(n_1180)
);

NAND2xp33_ASAP7_75t_SL g1181 ( 
.A(n_869),
.B(n_782),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_967),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_950),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_910),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_919),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_921),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_924),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_909),
.B(n_782),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_949),
.B(n_787),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_921),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_935),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1188),
.A2(n_826),
.B(n_927),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1019),
.A2(n_967),
.B1(n_869),
.B2(n_902),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1000),
.B(n_841),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1006),
.A2(n_1048),
.B(n_1012),
.C(n_1009),
.Y(n_1195)
);

OA21x2_ASAP7_75t_L g1196 ( 
.A1(n_1048),
.A2(n_920),
.B(n_974),
.Y(n_1196)
);

NOR3xp33_ASAP7_75t_L g1197 ( 
.A(n_1090),
.B(n_955),
.C(n_892),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1016),
.A2(n_877),
.B(n_869),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1016),
.A2(n_902),
.B(n_877),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_1040),
.A2(n_992),
.A3(n_974),
.B(n_938),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1020),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_L g1202 ( 
.A(n_1049),
.B(n_929),
.C(n_911),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_997),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_997),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1001),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1062),
.A2(n_971),
.B(n_992),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1036),
.B(n_877),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_1067),
.Y(n_1208)
);

BUFx5_ASAP7_75t_L g1209 ( 
.A(n_1136),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1139),
.A2(n_971),
.B(n_940),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1189),
.A2(n_933),
.B(n_961),
.Y(n_1211)
);

NOR2xp67_ASAP7_75t_L g1212 ( 
.A(n_1149),
.B(n_929),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1045),
.A2(n_1168),
.B(n_1077),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1009),
.A2(n_827),
.B(n_934),
.C(n_965),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1016),
.A2(n_916),
.B(n_902),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1070),
.A2(n_940),
.B(n_935),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1001),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1014),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1060),
.A2(n_1075),
.A3(n_1082),
.B(n_1069),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1176),
.B(n_861),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1070),
.A2(n_961),
.B(n_866),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1147),
.B(n_908),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1003),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1014),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1177),
.B(n_990),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1032),
.B(n_917),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1042),
.B(n_925),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1176),
.A2(n_1115),
.B1(n_1095),
.B2(n_1079),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1042),
.B(n_1054),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_999),
.Y(n_1230)
);

NOR2x1_ASAP7_75t_L g1231 ( 
.A(n_1116),
.B(n_924),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1034),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1070),
.A2(n_945),
.B(n_944),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_SL g1234 ( 
.A(n_1029),
.B(n_868),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1077),
.A2(n_945),
.B(n_944),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1106),
.B(n_954),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1140),
.A2(n_1004),
.B(n_1152),
.C(n_1151),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1054),
.B(n_930),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1077),
.A2(n_952),
.B(n_947),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1137),
.A2(n_1148),
.B(n_1158),
.Y(n_1240)
);

NOR2x1_ASAP7_75t_R g1241 ( 
.A(n_1051),
.B(n_954),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1073),
.A2(n_916),
.B1(n_824),
.B2(n_928),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1059),
.B(n_868),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_SL g1244 ( 
.A1(n_1036),
.A2(n_1109),
.B(n_1025),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1059),
.B(n_943),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1114),
.B(n_993),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_1060),
.A2(n_962),
.B(n_956),
.Y(n_1247)
);

AOI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1021),
.A2(n_964),
.B(n_959),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1027),
.A2(n_976),
.B(n_972),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1034),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1114),
.B(n_985),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1151),
.A2(n_970),
.B(n_973),
.C(n_968),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1148),
.A2(n_961),
.B(n_978),
.Y(n_1253)
);

NAND2x1_ASAP7_75t_L g1254 ( 
.A(n_1036),
.B(n_975),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1034),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1029),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1069),
.A2(n_966),
.A3(n_988),
.B(n_986),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1074),
.A2(n_1087),
.B1(n_1067),
.B2(n_1084),
.Y(n_1258)
);

AOI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1075),
.A2(n_1088),
.B(n_1082),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1109),
.A2(n_976),
.B(n_972),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_998),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1088),
.A2(n_1120),
.B(n_1094),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1111),
.B(n_942),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1015),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1016),
.A2(n_916),
.B(n_922),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1067),
.A2(n_928),
.B1(n_941),
.B2(n_932),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1148),
.A2(n_982),
.B(n_978),
.Y(n_1267)
);

NOR2x1_ASAP7_75t_L g1268 ( 
.A(n_998),
.B(n_924),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_999),
.B(n_874),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1123),
.B(n_873),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_SL g1271 ( 
.A1(n_1015),
.A2(n_977),
.B(n_982),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1158),
.A2(n_988),
.B(n_986),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1158),
.A2(n_966),
.B(n_989),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1127),
.A2(n_977),
.B(n_989),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1043),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1065),
.B(n_932),
.Y(n_1276)
);

NAND2x1_ASAP7_75t_L g1277 ( 
.A(n_1057),
.B(n_1136),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1162),
.A2(n_984),
.B(n_975),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_SL g1279 ( 
.A1(n_1025),
.A2(n_706),
.B(n_820),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1131),
.B(n_932),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1046),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1064),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1016),
.A2(n_984),
.B(n_928),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1131),
.A2(n_1026),
.B(n_1056),
.C(n_1047),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1061),
.A2(n_984),
.B(n_904),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1061),
.A2(n_787),
.B(n_706),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1124),
.B(n_787),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1026),
.A2(n_433),
.B(n_428),
.C(n_445),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1079),
.B(n_339),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1010),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1061),
.A2(n_672),
.B(n_663),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1156),
.A2(n_1100),
.B(n_1089),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1047),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1162),
.A2(n_383),
.B(n_373),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1099),
.B(n_373),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1099),
.B(n_389),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1166),
.B(n_1008),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1102),
.A2(n_820),
.B(n_653),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1166),
.B(n_390),
.Y(n_1299)
);

NOR2xp67_ASAP7_75t_L g1300 ( 
.A(n_1024),
.B(n_663),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1056),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1061),
.A2(n_672),
.B(n_663),
.Y(n_1302)
);

NAND2x1_ASAP7_75t_L g1303 ( 
.A(n_1057),
.B(n_663),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1094),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1093),
.B(n_668),
.Y(n_1305)
);

AOI211x1_ASAP7_75t_L g1306 ( 
.A1(n_1103),
.A2(n_425),
.B(n_420),
.C(n_428),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1061),
.A2(n_672),
.B(n_663),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1061),
.A2(n_682),
.B(n_672),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1008),
.B(n_390),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1181),
.A2(n_682),
.B(n_672),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1104),
.A2(n_682),
.B(n_728),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1162),
.A2(n_415),
.B(n_392),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1044),
.B(n_416),
.Y(n_1313)
);

NOR2x1_ASAP7_75t_SL g1314 ( 
.A(n_1175),
.B(n_682),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1120),
.A2(n_420),
.B(n_419),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1112),
.A2(n_780),
.B(n_728),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1121),
.A2(n_425),
.B(n_419),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1121),
.A2(n_433),
.B(n_682),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1093),
.B(n_1101),
.Y(n_1319)
);

AOI221x1_ASAP7_75t_L g1320 ( 
.A1(n_1178),
.A2(n_305),
.B1(n_248),
.B2(n_350),
.C(n_236),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1143),
.A2(n_745),
.B(n_728),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1124),
.B(n_248),
.Y(n_1322)
);

CKINVDCx6p67_ASAP7_75t_R g1323 ( 
.A(n_1010),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1003),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1143),
.A2(n_745),
.B(n_728),
.Y(n_1325)
);

INVxp67_ASAP7_75t_SL g1326 ( 
.A(n_1107),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1044),
.B(n_13),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1113),
.A2(n_780),
.B(n_728),
.Y(n_1328)
);

O2A1O1Ixp5_ASAP7_75t_L g1329 ( 
.A1(n_1124),
.A2(n_305),
.B(n_248),
.C(n_350),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1079),
.B(n_333),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1017),
.A2(n_780),
.B(n_247),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1130),
.B(n_248),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1017),
.A2(n_780),
.B(n_249),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_SL g1334 ( 
.A1(n_1175),
.A2(n_236),
.B(n_241),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1146),
.A2(n_437),
.A3(n_413),
.B(n_333),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1043),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1017),
.A2(n_780),
.B(n_253),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_SL g1338 ( 
.A1(n_1175),
.A2(n_236),
.B(n_252),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1085),
.A2(n_305),
.B(n_350),
.C(n_248),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1146),
.A2(n_745),
.B(n_437),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1153),
.A2(n_260),
.B(n_257),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1129),
.A2(n_305),
.B(n_350),
.C(n_236),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1153),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1064),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1068),
.B(n_14),
.Y(n_1345)
);

INVx5_ASAP7_75t_L g1346 ( 
.A(n_1057),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1068),
.B(n_17),
.Y(n_1347)
);

AND2x6_ASAP7_75t_L g1348 ( 
.A(n_1064),
.B(n_745),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1160),
.A2(n_413),
.B(n_437),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1160),
.A2(n_148),
.B(n_110),
.Y(n_1350)
);

AO31x2_ASAP7_75t_L g1351 ( 
.A1(n_1167),
.A2(n_305),
.A3(n_350),
.B(n_22),
.Y(n_1351)
);

NAND2xp33_ASAP7_75t_L g1352 ( 
.A(n_1136),
.B(n_305),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1135),
.B(n_18),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1083),
.A2(n_438),
.B(n_435),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1084),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1213),
.A2(n_1169),
.B(n_1167),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1203),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1204),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1213),
.A2(n_1170),
.B(n_1169),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1352),
.A2(n_1175),
.B(n_1083),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1220),
.B(n_1013),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1256),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1195),
.A2(n_1136),
.B(n_1157),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1284),
.A2(n_1339),
.B(n_1244),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1211),
.A2(n_1185),
.B(n_1170),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1346),
.Y(n_1366)
);

O2A1O1Ixp33_ASAP7_75t_SL g1367 ( 
.A1(n_1195),
.A2(n_1031),
.B(n_1002),
.C(n_1053),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1229),
.B(n_1101),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1202),
.A2(n_1084),
.B1(n_1119),
.B2(n_1096),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1211),
.A2(n_1186),
.B(n_1185),
.Y(n_1370)
);

NAND3xp33_ASAP7_75t_SL g1371 ( 
.A(n_1197),
.B(n_1052),
.C(n_1134),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1259),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1205),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1210),
.A2(n_1190),
.B(n_1186),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1217),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1261),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1262),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1346),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1197),
.A2(n_1098),
.B(n_1037),
.C(n_1091),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1297),
.B(n_1178),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1346),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1284),
.A2(n_1164),
.B(n_1190),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1223),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1262),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1346),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1267),
.A2(n_1191),
.B(n_1007),
.Y(n_1386)
);

AOI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1248),
.A2(n_1191),
.B(n_1007),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1220),
.A2(n_1228),
.B1(n_1117),
.B2(n_1269),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1299),
.A2(n_1071),
.B1(n_1134),
.B2(n_1163),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1246),
.A2(n_1081),
.B(n_1076),
.C(n_1063),
.Y(n_1390)
);

BUFx2_ASAP7_75t_R g1391 ( 
.A(n_1201),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1355),
.B(n_1013),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1355),
.B(n_1125),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1230),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1267),
.A2(n_1011),
.B(n_1005),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1330),
.A2(n_1163),
.B1(n_1105),
.B2(n_1117),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1272),
.A2(n_1011),
.B(n_1005),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1319),
.B(n_1125),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1230),
.B(n_1117),
.Y(n_1399)
);

AOI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1288),
.A2(n_1050),
.B1(n_1051),
.B2(n_1097),
.C(n_1072),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1272),
.A2(n_1030),
.B(n_1023),
.Y(n_1401)
);

OAI21xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1207),
.A2(n_1031),
.B(n_1002),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1277),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1256),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1273),
.A2(n_1030),
.B(n_1023),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1252),
.A2(n_1136),
.B(n_1154),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1319),
.B(n_1125),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1218),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1224),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1324),
.Y(n_1410)
);

AOI21xp33_ASAP7_75t_L g1411 ( 
.A1(n_1225),
.A2(n_1184),
.B(n_1165),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1216),
.A2(n_1038),
.B(n_1033),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1233),
.A2(n_1038),
.B(n_1033),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1264),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1251),
.B(n_1050),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1201),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1219),
.B(n_1180),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1348),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1219),
.B(n_1180),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1235),
.A2(n_1041),
.B(n_1039),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1290),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1245),
.A2(n_1018),
.B(n_1053),
.C(n_1173),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1239),
.A2(n_1041),
.B(n_1039),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1243),
.A2(n_1119),
.B1(n_1083),
.B2(n_1031),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1206),
.A2(n_1066),
.B(n_1055),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1194),
.B(n_1174),
.Y(n_1426)
);

INVxp67_ASAP7_75t_SL g1427 ( 
.A(n_1352),
.Y(n_1427)
);

INVx6_ASAP7_75t_L g1428 ( 
.A(n_1208),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1281),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1319),
.B(n_1028),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1262),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1289),
.B(n_1174),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1348),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1340),
.A2(n_1066),
.B(n_1055),
.Y(n_1434)
);

CKINVDCx6p67_ASAP7_75t_R g1435 ( 
.A(n_1323),
.Y(n_1435)
);

BUFx2_ASAP7_75t_SL g1436 ( 
.A(n_1209),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1348),
.Y(n_1437)
);

CKINVDCx11_ASAP7_75t_R g1438 ( 
.A(n_1290),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1293),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1236),
.B(n_1174),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1252),
.A2(n_1136),
.B(n_1154),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1237),
.B(n_1022),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1326),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1247),
.Y(n_1444)
);

INVx3_ASAP7_75t_SL g1445 ( 
.A(n_1208),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1320),
.A2(n_1086),
.B(n_1080),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1237),
.B(n_1022),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1275),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1227),
.B(n_1022),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1340),
.A2(n_1086),
.B(n_1080),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1282),
.B(n_1028),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1292),
.A2(n_1136),
.B(n_1173),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1275),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1253),
.A2(n_1128),
.B(n_1092),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1253),
.A2(n_1128),
.B(n_1092),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1193),
.A2(n_1173),
.B(n_1132),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_SL g1457 ( 
.A1(n_1271),
.A2(n_1179),
.B(n_1141),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1263),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1327),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1301),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1350),
.A2(n_1141),
.B(n_1138),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1304),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1343),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1345),
.Y(n_1464)
);

NAND2x1_ASAP7_75t_L g1465 ( 
.A(n_1279),
.B(n_1057),
.Y(n_1465)
);

AO21x2_ASAP7_75t_L g1466 ( 
.A1(n_1339),
.A2(n_1142),
.B(n_1138),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1269),
.A2(n_1097),
.B1(n_1161),
.B2(n_1145),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1219),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1219),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1350),
.A2(n_1150),
.B(n_1142),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1247),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1341),
.A2(n_1132),
.B(n_1130),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1265),
.A2(n_1118),
.B(n_1107),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1247),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1257),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1192),
.A2(n_1155),
.B(n_1150),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1257),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1348),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1260),
.A2(n_1183),
.B(n_1155),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_SL g1480 ( 
.A1(n_1314),
.A2(n_1179),
.B(n_1183),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1295),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1296),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1232),
.B(n_1250),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1234),
.B(n_1105),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1255),
.A2(n_1133),
.B1(n_1144),
.B2(n_1145),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1212),
.A2(n_1133),
.B1(n_1144),
.B2(n_1161),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1222),
.B(n_1238),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1274),
.A2(n_1179),
.B(n_1133),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1192),
.A2(n_1221),
.B(n_1240),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_SL g1490 ( 
.A1(n_1249),
.A2(n_1057),
.B(n_1107),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1221),
.A2(n_1132),
.B(n_1130),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1257),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1329),
.A2(n_1122),
.B(n_267),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1258),
.A2(n_1144),
.B1(n_1057),
.B2(n_1035),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1196),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1200),
.B(n_1108),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1200),
.B(n_1110),
.Y(n_1497)
);

NAND2x1p5_ASAP7_75t_L g1498 ( 
.A(n_1303),
.B(n_1107),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1226),
.A2(n_1172),
.B1(n_1187),
.B2(n_1159),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1318),
.A2(n_1118),
.B(n_1107),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1278),
.A2(n_1126),
.B(n_1118),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1270),
.A2(n_1144),
.B1(n_1159),
.B2(n_1187),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1309),
.Y(n_1503)
);

AOI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1322),
.A2(n_1122),
.B(n_1064),
.Y(n_1504)
);

NAND2x1p5_ASAP7_75t_L g1505 ( 
.A(n_1275),
.B(n_1118),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1196),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1196),
.Y(n_1507)
);

AOI221x1_ASAP7_75t_L g1508 ( 
.A1(n_1214),
.A2(n_1126),
.B1(n_1118),
.B2(n_1171),
.C(n_1182),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1313),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1214),
.A2(n_1122),
.B(n_266),
.Y(n_1510)
);

O2A1O1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1342),
.A2(n_1110),
.B(n_1122),
.C(n_1172),
.Y(n_1511)
);

INVx6_ASAP7_75t_L g1512 ( 
.A(n_1305),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1275),
.Y(n_1513)
);

BUFx12f_ASAP7_75t_L g1514 ( 
.A(n_1336),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1200),
.Y(n_1515)
);

INVx5_ASAP7_75t_L g1516 ( 
.A(n_1348),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1198),
.A2(n_1126),
.B(n_1182),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1282),
.B(n_1171),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1241),
.B(n_1172),
.Y(n_1519)
);

OAI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1347),
.A2(n_1058),
.B1(n_1043),
.B2(n_1182),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1315),
.A2(n_1126),
.B(n_1057),
.Y(n_1521)
);

NOR2xp67_ASAP7_75t_L g1522 ( 
.A(n_1353),
.B(n_1171),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1200),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1344),
.B(n_1043),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1344),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1280),
.B(n_1043),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1305),
.B(n_1058),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1342),
.A2(n_350),
.B(n_1058),
.Y(n_1528)
);

AO21x2_ASAP7_75t_L g1529 ( 
.A1(n_1349),
.A2(n_1126),
.B(n_1171),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1276),
.B(n_1171),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1317),
.Y(n_1531)
);

INVx4_ASAP7_75t_L g1532 ( 
.A(n_1305),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1242),
.A2(n_1058),
.B1(n_1182),
.B2(n_1078),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1294),
.A2(n_1078),
.B(n_1182),
.Y(n_1534)
);

O2A1O1Ixp33_ASAP7_75t_SL g1535 ( 
.A1(n_1207),
.A2(n_1078),
.B(n_1058),
.C(n_25),
.Y(n_1535)
);

AOI222xp33_ASAP7_75t_L g1536 ( 
.A1(n_1361),
.A2(n_1288),
.B1(n_1231),
.B2(n_1300),
.C1(n_1349),
.C2(n_1268),
.Y(n_1536)
);

BUFx4f_ASAP7_75t_L g1537 ( 
.A(n_1435),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1508),
.A2(n_1312),
.B(n_1322),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1400),
.A2(n_1306),
.B1(n_1338),
.B2(n_1334),
.C(n_1354),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1387),
.A2(n_1285),
.B(n_1283),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1376),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1357),
.Y(n_1542)
);

INVx6_ASAP7_75t_L g1543 ( 
.A(n_1514),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1416),
.Y(n_1544)
);

NAND3xp33_ASAP7_75t_L g1545 ( 
.A(n_1379),
.B(n_1332),
.C(n_1336),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1487),
.B(n_1335),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1358),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1380),
.B(n_1335),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1373),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1375),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1388),
.A2(n_1266),
.B1(n_1326),
.B2(n_1332),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1415),
.A2(n_1298),
.B1(n_1209),
.B2(n_1336),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1514),
.Y(n_1553)
);

AOI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1387),
.A2(n_1287),
.B(n_1310),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1389),
.A2(n_1209),
.B1(n_1336),
.B2(n_1287),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1380),
.B(n_1335),
.Y(n_1556)
);

OAI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1363),
.A2(n_1311),
.B1(n_1286),
.B2(n_1254),
.C(n_268),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1449),
.A2(n_1199),
.B1(n_1215),
.B2(n_1078),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1408),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1376),
.Y(n_1560)
);

AOI221xp5_ASAP7_75t_L g1561 ( 
.A1(n_1371),
.A2(n_370),
.B1(n_273),
.B2(n_288),
.C(n_293),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1392),
.A2(n_1209),
.B1(n_1078),
.B2(n_1335),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1409),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1442),
.A2(n_1316),
.B1(n_1291),
.B2(n_1302),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1368),
.B(n_18),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1394),
.B(n_1351),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1435),
.Y(n_1567)
);

O2A1O1Ixp33_ASAP7_75t_SL g1568 ( 
.A1(n_1447),
.A2(n_1209),
.B(n_1307),
.C(n_1308),
.Y(n_1568)
);

INVx4_ASAP7_75t_SL g1569 ( 
.A(n_1433),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1398),
.B(n_1351),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1481),
.A2(n_1209),
.B1(n_1328),
.B2(n_1351),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1458),
.B(n_26),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1503),
.B(n_31),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1482),
.A2(n_1321),
.B1(n_1325),
.B2(n_272),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1453),
.Y(n_1575)
);

AOI21xp33_ASAP7_75t_L g1576 ( 
.A1(n_1422),
.A2(n_1510),
.B(n_1426),
.Y(n_1576)
);

NAND2x1p5_ASAP7_75t_L g1577 ( 
.A(n_1516),
.B(n_1321),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1398),
.B(n_1325),
.Y(n_1578)
);

AOI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1390),
.A2(n_361),
.B1(n_298),
.B2(n_308),
.C(n_434),
.Y(n_1579)
);

NAND2x1p5_ASAP7_75t_L g1580 ( 
.A(n_1516),
.B(n_1331),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1427),
.A2(n_1369),
.B1(n_1432),
.B2(n_1399),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1414),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1509),
.A2(n_1488),
.B1(n_1459),
.B2(n_1464),
.Y(n_1583)
);

NAND3xp33_ASAP7_75t_L g1584 ( 
.A(n_1424),
.B(n_1486),
.C(n_1510),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1394),
.B(n_35),
.Y(n_1585)
);

A2O1A1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1528),
.A2(n_1337),
.B(n_1333),
.C(n_426),
.Y(n_1586)
);

INVxp67_ASAP7_75t_L g1587 ( 
.A(n_1443),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1488),
.A2(n_422),
.B1(n_421),
.B2(n_404),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1439),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1460),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1462),
.Y(n_1591)
);

CKINVDCx16_ASAP7_75t_R g1592 ( 
.A(n_1362),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1398),
.B(n_39),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1463),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1438),
.Y(n_1595)
);

NAND2xp33_ASAP7_75t_R g1596 ( 
.A(n_1360),
.B(n_118),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1511),
.A2(n_395),
.B(n_388),
.C(n_382),
.Y(n_1597)
);

OAI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1452),
.A2(n_375),
.B(n_374),
.Y(n_1598)
);

OAI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1396),
.A2(n_1440),
.B1(n_1467),
.B2(n_1502),
.C(n_1399),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1483),
.B(n_44),
.Y(n_1600)
);

NAND2xp33_ASAP7_75t_R g1601 ( 
.A(n_1443),
.B(n_119),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1429),
.B(n_46),
.Y(n_1602)
);

NAND2xp33_ASAP7_75t_SL g1603 ( 
.A(n_1445),
.B(n_294),
.Y(n_1603)
);

BUFx4f_ASAP7_75t_SL g1604 ( 
.A(n_1362),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1383),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1404),
.A2(n_368),
.B1(n_364),
.B2(n_359),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_1438),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1404),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1416),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1383),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1393),
.B(n_1421),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1407),
.B(n_46),
.Y(n_1612)
);

AND2x2_ASAP7_75t_SL g1613 ( 
.A(n_1433),
.B(n_1496),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1410),
.Y(n_1614)
);

OR2x6_ASAP7_75t_L g1615 ( 
.A(n_1433),
.B(n_128),
.Y(n_1615)
);

AOI21xp33_ASAP7_75t_L g1616 ( 
.A1(n_1510),
.A2(n_358),
.B(n_357),
.Y(n_1616)
);

OR2x6_ASAP7_75t_L g1617 ( 
.A(n_1433),
.B(n_132),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1483),
.B(n_47),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1417),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1488),
.A2(n_356),
.B1(n_348),
.B2(n_347),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1445),
.A2(n_341),
.B1(n_334),
.B2(n_324),
.Y(n_1621)
);

NAND2x1_ASAP7_75t_L g1622 ( 
.A(n_1403),
.B(n_215),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1532),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1417),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1393),
.B(n_49),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1484),
.A2(n_1494),
.B1(n_1485),
.B2(n_1519),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1419),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1411),
.A2(n_323),
.B1(n_315),
.B2(n_52),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1421),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1430),
.B(n_50),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1532),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_1631)
);

OAI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1419),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1468),
.Y(n_1633)
);

NAND2x1p5_ASAP7_75t_L g1634 ( 
.A(n_1516),
.B(n_214),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1469),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1382),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1475),
.Y(n_1637)
);

NAND2x1p5_ASAP7_75t_L g1638 ( 
.A(n_1516),
.B(n_213),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1469),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_SL g1640 ( 
.A1(n_1382),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1382),
.A2(n_1407),
.B1(n_1364),
.B2(n_1477),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1496),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1430),
.B(n_59),
.Y(n_1643)
);

INVx5_ASAP7_75t_SL g1644 ( 
.A(n_1433),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1430),
.B(n_60),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1532),
.Y(n_1646)
);

CKINVDCx16_ASAP7_75t_R g1647 ( 
.A(n_1448),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1448),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1407),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1428),
.A2(n_61),
.B1(n_68),
.B2(n_69),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1364),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_1651)
);

OAI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1516),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1367),
.A2(n_73),
.B(n_76),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1364),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1406),
.A2(n_83),
.B(n_84),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1428),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_1656)
);

INVx4_ASAP7_75t_SL g1657 ( 
.A(n_1428),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1451),
.B(n_86),
.Y(n_1658)
);

AOI21xp33_ASAP7_75t_L g1659 ( 
.A1(n_1497),
.A2(n_89),
.B(n_91),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1512),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1441),
.A2(n_89),
.B(n_92),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1451),
.B(n_92),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1477),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_1663)
);

OR2x6_ASAP7_75t_L g1664 ( 
.A(n_1378),
.B(n_199),
.Y(n_1664)
);

NOR3xp33_ASAP7_75t_SL g1665 ( 
.A(n_1402),
.B(n_98),
.C(n_100),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1451),
.B(n_101),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1492),
.A2(n_1497),
.B1(n_1506),
.B2(n_1512),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1530),
.B(n_133),
.Y(n_1668)
);

CKINVDCx6p67_ASAP7_75t_R g1669 ( 
.A(n_1453),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1492),
.A2(n_1506),
.B1(n_1512),
.B2(n_1507),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1512),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1372),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1489),
.A2(n_141),
.B(n_146),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1391),
.Y(n_1674)
);

OAI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1456),
.A2(n_147),
.B(n_149),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1428),
.Y(n_1676)
);

AOI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1372),
.A2(n_151),
.B1(n_157),
.B2(n_169),
.C(n_174),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_SL g1678 ( 
.A1(n_1495),
.A2(n_178),
.B1(n_179),
.B2(n_186),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1525),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1386),
.Y(n_1680)
);

AND2x6_ASAP7_75t_L g1681 ( 
.A(n_1418),
.B(n_187),
.Y(n_1681)
);

AOI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1499),
.A2(n_192),
.B1(n_193),
.B2(n_197),
.C(n_198),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1508),
.A2(n_1473),
.B(n_1517),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1386),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1495),
.A2(n_1507),
.B1(n_1515),
.B2(n_1523),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1513),
.Y(n_1686)
);

BUFx4f_ASAP7_75t_SL g1687 ( 
.A(n_1524),
.Y(n_1687)
);

A2O1A1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1522),
.A2(n_1472),
.B(n_1515),
.C(n_1523),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1466),
.A2(n_1479),
.B1(n_1527),
.B2(n_1471),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1518),
.B(n_1525),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1518),
.B(n_1527),
.Y(n_1691)
);

BUFx10_ASAP7_75t_L g1692 ( 
.A(n_1524),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1527),
.B(n_1524),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1374),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1466),
.A2(n_1479),
.B1(n_1444),
.B2(n_1474),
.Y(n_1695)
);

OAI21x1_ASAP7_75t_L g1696 ( 
.A1(n_1489),
.A2(n_1450),
.B(n_1434),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_SL g1697 ( 
.A1(n_1457),
.A2(n_1446),
.B1(n_1480),
.B2(n_1466),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1377),
.A2(n_1431),
.B1(n_1384),
.B2(n_1535),
.C(n_1457),
.Y(n_1698)
);

INVx8_ASAP7_75t_L g1699 ( 
.A(n_1418),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1479),
.A2(n_1444),
.B1(n_1471),
.B2(n_1474),
.Y(n_1700)
);

AO21x2_ASAP7_75t_L g1701 ( 
.A1(n_1480),
.A2(n_1490),
.B(n_1434),
.Y(n_1701)
);

AO21x2_ASAP7_75t_L g1702 ( 
.A1(n_1490),
.A2(n_1450),
.B(n_1470),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1377),
.A2(n_1431),
.B1(n_1384),
.B2(n_1526),
.C(n_1520),
.Y(n_1703)
);

OAI221xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1531),
.A2(n_1403),
.B1(n_1437),
.B2(n_1418),
.C(n_1478),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1381),
.Y(n_1705)
);

OAI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1437),
.A2(n_1478),
.B1(n_1381),
.B2(n_1385),
.Y(n_1706)
);

NAND2xp33_ASAP7_75t_SL g1707 ( 
.A(n_1381),
.B(n_1385),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1446),
.A2(n_1478),
.B1(n_1436),
.B2(n_1493),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1529),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1381),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1446),
.A2(n_1476),
.B1(n_1529),
.B2(n_1493),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1374),
.Y(n_1712)
);

AO21x2_ASAP7_75t_L g1713 ( 
.A1(n_1461),
.A2(n_1470),
.B(n_1529),
.Y(n_1713)
);

NOR2x1_ASAP7_75t_SL g1714 ( 
.A(n_1381),
.B(n_1385),
.Y(n_1714)
);

BUFx8_ASAP7_75t_L g1715 ( 
.A(n_1385),
.Y(n_1715)
);

INVx4_ASAP7_75t_L g1716 ( 
.A(n_1505),
.Y(n_1716)
);

CKINVDCx6p67_ASAP7_75t_R g1717 ( 
.A(n_1385),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1505),
.Y(n_1718)
);

INVx5_ASAP7_75t_L g1719 ( 
.A(n_1378),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1476),
.A2(n_1493),
.B1(n_1365),
.B2(n_1370),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1476),
.A2(n_1370),
.B1(n_1533),
.B2(n_1359),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1465),
.A2(n_1501),
.B(n_1521),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1589),
.B(n_1356),
.Y(n_1723)
);

NAND3xp33_ASAP7_75t_L g1724 ( 
.A(n_1651),
.B(n_1403),
.C(n_1465),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_SL g1725 ( 
.A1(n_1584),
.A2(n_1436),
.B1(n_1378),
.B2(n_1366),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1632),
.A2(n_1366),
.B1(n_1498),
.B2(n_1461),
.C(n_1423),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1632),
.A2(n_1454),
.B1(n_1455),
.B2(n_1405),
.Y(n_1727)
);

INVxp33_ASAP7_75t_SL g1728 ( 
.A(n_1674),
.Y(n_1728)
);

OAI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1601),
.A2(n_1631),
.B1(n_1626),
.B2(n_1652),
.Y(n_1729)
);

INVx4_ASAP7_75t_L g1730 ( 
.A(n_1676),
.Y(n_1730)
);

OAI322xp33_ASAP7_75t_L g1731 ( 
.A1(n_1652),
.A2(n_1498),
.A3(n_1366),
.B1(n_1504),
.B2(n_1425),
.C1(n_1423),
.C2(n_1412),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1675),
.A2(n_1521),
.B(n_1501),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1629),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1651),
.A2(n_1455),
.B1(n_1454),
.B2(n_1405),
.Y(n_1734)
);

OAI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1654),
.A2(n_1504),
.B1(n_1420),
.B2(n_1413),
.C(n_1412),
.Y(n_1735)
);

AO221x1_ASAP7_75t_L g1736 ( 
.A1(n_1575),
.A2(n_1534),
.B1(n_1491),
.B2(n_1500),
.C(n_1413),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1541),
.Y(n_1737)
);

AOI211xp5_ASAP7_75t_L g1738 ( 
.A1(n_1650),
.A2(n_1491),
.B(n_1534),
.C(n_1500),
.Y(n_1738)
);

OA21x2_ASAP7_75t_L g1739 ( 
.A1(n_1696),
.A2(n_1425),
.B(n_1397),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1542),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1575),
.B(n_1395),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1649),
.A2(n_1420),
.B1(n_1397),
.B2(n_1401),
.Y(n_1742)
);

AO31x2_ASAP7_75t_L g1743 ( 
.A1(n_1688),
.A2(n_1401),
.A3(n_1564),
.B(n_1683),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1547),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1649),
.A2(n_1654),
.B1(n_1663),
.B2(n_1665),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1601),
.A2(n_1612),
.B1(n_1593),
.B2(n_1596),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1640),
.A2(n_1636),
.B1(n_1663),
.B2(n_1628),
.Y(n_1747)
);

OAI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1596),
.A2(n_1599),
.B1(n_1592),
.B2(n_1655),
.Y(n_1748)
);

CKINVDCx20_ASAP7_75t_R g1749 ( 
.A(n_1604),
.Y(n_1749)
);

BUFx4f_ASAP7_75t_SL g1750 ( 
.A(n_1669),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1640),
.A2(n_1636),
.B1(n_1628),
.B2(n_1588),
.Y(n_1751)
);

CKINVDCx6p67_ASAP7_75t_R g1752 ( 
.A(n_1607),
.Y(n_1752)
);

OAI21x1_ASAP7_75t_L g1753 ( 
.A1(n_1540),
.A2(n_1554),
.B(n_1722),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1587),
.Y(n_1754)
);

NAND3xp33_ASAP7_75t_L g1755 ( 
.A(n_1665),
.B(n_1620),
.C(n_1588),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1587),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1620),
.A2(n_1546),
.B1(n_1659),
.B2(n_1583),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1661),
.A2(n_1593),
.B1(n_1612),
.B2(n_1604),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1616),
.A2(n_1572),
.B1(n_1573),
.B2(n_1576),
.C(n_1602),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1543),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1583),
.A2(n_1539),
.B1(n_1548),
.B2(n_1556),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1691),
.B(n_1565),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1608),
.A2(n_1585),
.B1(n_1658),
.B2(n_1662),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1568),
.A2(n_1653),
.B(n_1704),
.Y(n_1764)
);

BUFx12f_ASAP7_75t_L g1765 ( 
.A(n_1544),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1549),
.Y(n_1766)
);

OA21x2_ASAP7_75t_L g1767 ( 
.A1(n_1711),
.A2(n_1709),
.B(n_1689),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1570),
.A2(n_1562),
.B1(n_1678),
.B2(n_1656),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1613),
.A2(n_1681),
.B1(n_1625),
.B2(n_1615),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1550),
.Y(n_1770)
);

NAND4xp25_ASAP7_75t_L g1771 ( 
.A(n_1600),
.B(n_1618),
.C(n_1595),
.D(n_1666),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1559),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1545),
.A2(n_1645),
.B1(n_1643),
.B2(n_1551),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1693),
.B(n_1647),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1562),
.A2(n_1678),
.B1(n_1536),
.B2(n_1617),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1568),
.A2(n_1704),
.B(n_1707),
.Y(n_1776)
);

BUFx4f_ASAP7_75t_SL g1777 ( 
.A(n_1595),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1566),
.B(n_1582),
.Y(n_1778)
);

OR2x2_ASAP7_75t_SL g1779 ( 
.A(n_1543),
.B(n_1590),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_SL g1780 ( 
.A1(n_1681),
.A2(n_1617),
.B1(n_1615),
.B2(n_1581),
.Y(n_1780)
);

OAI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1537),
.A2(n_1555),
.B1(n_1597),
.B2(n_1664),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1609),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1664),
.A2(n_1615),
.B1(n_1617),
.B2(n_1687),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1537),
.A2(n_1555),
.B1(n_1664),
.B2(n_1552),
.Y(n_1784)
);

BUFx4f_ASAP7_75t_SL g1785 ( 
.A(n_1553),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1591),
.A2(n_1594),
.B1(n_1681),
.B2(n_1630),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1552),
.A2(n_1598),
.B1(n_1567),
.B2(n_1686),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1690),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1672),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1681),
.A2(n_1677),
.B1(n_1624),
.B2(n_1627),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1558),
.A2(n_1706),
.B(n_1586),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1569),
.B(n_1648),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1681),
.A2(n_1642),
.B1(n_1703),
.B2(n_1679),
.Y(n_1793)
);

AOI33xp33_ASAP7_75t_L g1794 ( 
.A1(n_1571),
.A2(n_1579),
.A3(n_1561),
.B1(n_1560),
.B2(n_1697),
.B3(n_1721),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1642),
.A2(n_1682),
.B1(n_1619),
.B2(n_1641),
.Y(n_1795)
);

AOI222xp33_ASAP7_75t_L g1796 ( 
.A1(n_1606),
.A2(n_1603),
.B1(n_1641),
.B2(n_1667),
.C1(n_1633),
.C2(n_1639),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1571),
.A2(n_1693),
.B1(n_1671),
.B2(n_1687),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1667),
.A2(n_1668),
.B1(n_1670),
.B2(n_1635),
.Y(n_1798)
);

OAI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1660),
.A2(n_1634),
.B1(n_1638),
.B2(n_1543),
.Y(n_1799)
);

OAI21xp33_ASAP7_75t_L g1800 ( 
.A1(n_1721),
.A2(n_1698),
.B(n_1621),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1605),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1610),
.B(n_1614),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_1692),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1670),
.A2(n_1660),
.B1(n_1578),
.B2(n_1638),
.Y(n_1804)
);

OAI21x1_ASAP7_75t_L g1805 ( 
.A1(n_1720),
.A2(n_1673),
.B(n_1711),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1623),
.A2(n_1646),
.B1(n_1553),
.B2(n_1574),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1578),
.A2(n_1634),
.B1(n_1700),
.B2(n_1697),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1700),
.A2(n_1644),
.B1(n_1689),
.B2(n_1692),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1623),
.A2(n_1646),
.B1(n_1574),
.B2(n_1557),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1644),
.A2(n_1685),
.B1(n_1695),
.B2(n_1637),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1718),
.B(n_1657),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1694),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1712),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1716),
.B(n_1657),
.Y(n_1814)
);

AOI211xp5_ASAP7_75t_L g1815 ( 
.A1(n_1706),
.A2(n_1709),
.B(n_1684),
.C(n_1680),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1622),
.A2(n_1708),
.B(n_1538),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1644),
.A2(n_1685),
.B1(n_1695),
.B2(n_1538),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_SL g1818 ( 
.A1(n_1699),
.A2(n_1714),
.B1(n_1715),
.B2(n_1580),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1715),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1701),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1716),
.A2(n_1717),
.B1(n_1719),
.B2(n_1720),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1708),
.A2(n_1699),
.B1(n_1569),
.B2(n_1580),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1699),
.A2(n_1705),
.B1(n_1710),
.B2(n_1719),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1713),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1705),
.A2(n_1710),
.B1(n_1577),
.B2(n_1702),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1705),
.A2(n_1710),
.B1(n_1702),
.B2(n_1713),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1563),
.B(n_1394),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1632),
.A2(n_1361),
.B1(n_1197),
.B2(n_589),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1632),
.A2(n_1361),
.B1(n_1197),
.B2(n_589),
.Y(n_1829)
);

AOI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1632),
.A2(n_1197),
.B1(n_823),
.B2(n_1361),
.C(n_830),
.Y(n_1830)
);

BUFx8_ASAP7_75t_SL g1831 ( 
.A(n_1674),
.Y(n_1831)
);

OAI222xp33_ASAP7_75t_L g1832 ( 
.A1(n_1632),
.A2(n_1166),
.B1(n_1176),
.B2(n_1228),
.C1(n_822),
.C2(n_1388),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1593),
.B(n_1006),
.Y(n_1833)
);

AOI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1632),
.A2(n_1197),
.B1(n_823),
.B2(n_1361),
.C(n_830),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1632),
.A2(n_1361),
.B1(n_1197),
.B2(n_589),
.Y(n_1835)
);

AOI33xp33_ASAP7_75t_L g1836 ( 
.A1(n_1649),
.A2(n_342),
.A3(n_228),
.B1(n_309),
.B2(n_303),
.B3(n_823),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1542),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1674),
.Y(n_1838)
);

OAI221xp5_ASAP7_75t_SL g1839 ( 
.A1(n_1651),
.A2(n_823),
.B1(n_1654),
.B2(n_830),
.C(n_834),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1632),
.A2(n_1361),
.B1(n_1197),
.B2(n_589),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1632),
.A2(n_1361),
.B1(n_1197),
.B2(n_589),
.Y(n_1841)
);

OAI221xp5_ASAP7_75t_L g1842 ( 
.A1(n_1651),
.A2(n_1006),
.B1(n_1361),
.B2(n_830),
.C(n_834),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1563),
.B(n_1394),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1649),
.A2(n_1006),
.B1(n_1361),
.B2(n_834),
.Y(n_1844)
);

OAI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1651),
.A2(n_1006),
.B1(n_1361),
.B2(n_830),
.C(n_834),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1632),
.A2(n_1361),
.B1(n_1197),
.B2(n_589),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_SL g1847 ( 
.A1(n_1652),
.A2(n_1379),
.B1(n_1632),
.B2(n_1006),
.C(n_996),
.Y(n_1847)
);

OAI211xp5_ASAP7_75t_SL g1848 ( 
.A1(n_1631),
.A2(n_852),
.B(n_1018),
.C(n_651),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1563),
.B(n_1394),
.Y(n_1849)
);

AOI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1632),
.A2(n_1197),
.B1(n_823),
.B2(n_1361),
.C(n_830),
.Y(n_1850)
);

INVxp33_ASAP7_75t_L g1851 ( 
.A(n_1575),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1691),
.B(n_1611),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1691),
.B(n_1611),
.Y(n_1853)
);

AOI222xp33_ASAP7_75t_L g1854 ( 
.A1(n_1632),
.A2(n_589),
.B1(n_1361),
.B2(n_817),
.C1(n_913),
.C2(n_823),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_SL g1855 ( 
.A1(n_1584),
.A2(n_1361),
.B1(n_913),
.B2(n_1176),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1541),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1691),
.B(n_1611),
.Y(n_1857)
);

INVx4_ASAP7_75t_L g1858 ( 
.A(n_1676),
.Y(n_1858)
);

AOI222xp33_ASAP7_75t_L g1859 ( 
.A1(n_1632),
.A2(n_589),
.B1(n_1361),
.B2(n_817),
.C1(n_913),
.C2(n_823),
.Y(n_1859)
);

AOI33xp33_ASAP7_75t_L g1860 ( 
.A1(n_1649),
.A2(n_342),
.A3(n_228),
.B1(n_309),
.B2(n_303),
.B3(n_823),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1649),
.A2(n_1006),
.B1(n_1361),
.B2(n_834),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1593),
.B(n_1006),
.Y(n_1862)
);

OAI21xp33_ASAP7_75t_L g1863 ( 
.A1(n_1651),
.A2(n_1006),
.B(n_834),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1632),
.A2(n_1361),
.B1(n_1197),
.B2(n_589),
.Y(n_1864)
);

OAI221xp5_ASAP7_75t_L g1865 ( 
.A1(n_1651),
.A2(n_1006),
.B1(n_1361),
.B2(n_830),
.C(n_834),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1632),
.A2(n_1361),
.B1(n_1197),
.B2(n_589),
.Y(n_1866)
);

OAI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1651),
.A2(n_1006),
.B1(n_1361),
.B2(n_830),
.C(n_834),
.Y(n_1867)
);

NAND2x1p5_ASAP7_75t_L g1868 ( 
.A(n_1719),
.B(n_1516),
.Y(n_1868)
);

AOI221xp5_ASAP7_75t_L g1869 ( 
.A1(n_1632),
.A2(n_1197),
.B1(n_823),
.B2(n_1361),
.C(n_830),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1601),
.A2(n_1361),
.B1(n_1006),
.B2(n_830),
.Y(n_1870)
);

OAI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1601),
.A2(n_1176),
.B1(n_1361),
.B2(n_1202),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1587),
.Y(n_1872)
);

OAI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1601),
.A2(n_1176),
.B1(n_1361),
.B2(n_1202),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1601),
.A2(n_1361),
.B1(n_1006),
.B2(n_830),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1632),
.A2(n_1361),
.B1(n_1197),
.B2(n_589),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1587),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1632),
.A2(n_1361),
.B1(n_1197),
.B2(n_589),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1593),
.B(n_1006),
.Y(n_1878)
);

AO21x2_ASAP7_75t_L g1879 ( 
.A1(n_1576),
.A2(n_1616),
.B(n_1387),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1632),
.A2(n_1197),
.B1(n_823),
.B2(n_1361),
.C(n_830),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1632),
.A2(n_1361),
.B1(n_1197),
.B2(n_589),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1672),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1542),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1754),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1852),
.B(n_1853),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1857),
.B(n_1882),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1882),
.Y(n_1887)
);

AND2x4_ASAP7_75t_L g1888 ( 
.A(n_1741),
.B(n_1826),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1741),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1756),
.B(n_1872),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1788),
.B(n_1827),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1843),
.B(n_1849),
.Y(n_1892)
);

INVxp67_ASAP7_75t_SL g1893 ( 
.A(n_1876),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1812),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1737),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1728),
.B(n_1730),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1856),
.B(n_1733),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1778),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1828),
.A2(n_1846),
.B1(n_1829),
.B2(n_1875),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1762),
.B(n_1789),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1740),
.B(n_1744),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1813),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1770),
.B(n_1772),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1801),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1733),
.B(n_1837),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1826),
.B(n_1792),
.Y(n_1906)
);

INVx3_ASAP7_75t_L g1907 ( 
.A(n_1805),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_SL g1908 ( 
.A(n_1838),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1883),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1779),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1723),
.Y(n_1911)
);

AO31x2_ASAP7_75t_L g1912 ( 
.A1(n_1742),
.A2(n_1820),
.A3(n_1824),
.B(n_1764),
.Y(n_1912)
);

INVx3_ASAP7_75t_L g1913 ( 
.A(n_1739),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1739),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1739),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1766),
.B(n_1761),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1807),
.B(n_1822),
.Y(n_1917)
);

CKINVDCx16_ASAP7_75t_R g1918 ( 
.A(n_1746),
.Y(n_1918)
);

NOR2x1_ASAP7_75t_L g1919 ( 
.A(n_1776),
.B(n_1783),
.Y(n_1919)
);

OAI211xp5_ASAP7_75t_L g1920 ( 
.A1(n_1870),
.A2(n_1874),
.B(n_1880),
.C(n_1869),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1802),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1730),
.B(n_1858),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1858),
.B(n_1749),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1774),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1767),
.B(n_1743),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1767),
.B(n_1743),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1771),
.B(n_1761),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1767),
.B(n_1743),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1816),
.B(n_1743),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_SL g1930 ( 
.A(n_1871),
.B(n_1873),
.Y(n_1930)
);

INVx3_ASAP7_75t_L g1931 ( 
.A(n_1753),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1817),
.B(n_1736),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1817),
.B(n_1815),
.Y(n_1933)
);

HB1xp67_ASAP7_75t_L g1934 ( 
.A(n_1825),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1763),
.B(n_1796),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1833),
.B(n_1862),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1798),
.B(n_1786),
.Y(n_1937)
);

INVx4_ASAP7_75t_R g1938 ( 
.A(n_1819),
.Y(n_1938)
);

AOI322xp5_ASAP7_75t_L g1939 ( 
.A1(n_1828),
.A2(n_1881),
.A3(n_1866),
.B1(n_1864),
.B2(n_1829),
.C1(n_1835),
.C2(n_1875),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1833),
.B(n_1862),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1731),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1735),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1806),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1879),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1879),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1798),
.B(n_1786),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1808),
.B(n_1795),
.Y(n_1947)
);

NOR2x1_ASAP7_75t_L g1948 ( 
.A(n_1724),
.B(n_1760),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1808),
.B(n_1797),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1727),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1878),
.B(n_1773),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1727),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1878),
.B(n_1830),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1811),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1797),
.B(n_1738),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1768),
.B(n_1734),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1821),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1768),
.B(n_1734),
.Y(n_1958)
);

BUFx2_ASAP7_75t_L g1959 ( 
.A(n_1803),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1793),
.B(n_1757),
.Y(n_1960)
);

NOR4xp25_ASAP7_75t_SL g1961 ( 
.A(n_1839),
.B(n_1865),
.C(n_1867),
.D(n_1842),
.Y(n_1961)
);

BUFx2_ASAP7_75t_L g1962 ( 
.A(n_1803),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1804),
.B(n_1810),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1804),
.B(n_1810),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1726),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1851),
.B(n_1793),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1780),
.B(n_1795),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1800),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1725),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1775),
.B(n_1769),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1732),
.Y(n_1971)
);

INVxp67_ASAP7_75t_L g1972 ( 
.A(n_1787),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1794),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1809),
.Y(n_1974)
);

INVxp67_ASAP7_75t_SL g1975 ( 
.A(n_1791),
.Y(n_1975)
);

OAI211xp5_ASAP7_75t_SL g1976 ( 
.A1(n_1939),
.A2(n_1845),
.B(n_1834),
.C(n_1850),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_SL g1977 ( 
.A1(n_1918),
.A2(n_1881),
.B1(n_1835),
.B2(n_1841),
.Y(n_1977)
);

AOI21xp33_ASAP7_75t_L g1978 ( 
.A1(n_1899),
.A2(n_1755),
.B(n_1844),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1887),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1887),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1898),
.B(n_1757),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1893),
.B(n_1759),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1902),
.Y(n_1983)
);

OAI211xp5_ASAP7_75t_L g1984 ( 
.A1(n_1939),
.A2(n_1841),
.B(n_1840),
.C(n_1864),
.Y(n_1984)
);

OA21x2_ASAP7_75t_L g1985 ( 
.A1(n_1914),
.A2(n_1775),
.B(n_1847),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1891),
.B(n_1745),
.Y(n_1986)
);

INVx5_ASAP7_75t_L g1987 ( 
.A(n_1907),
.Y(n_1987)
);

CKINVDCx16_ASAP7_75t_R g1988 ( 
.A(n_1910),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1886),
.B(n_1752),
.Y(n_1989)
);

AOI221xp5_ASAP7_75t_L g1990 ( 
.A1(n_1899),
.A2(n_1877),
.B1(n_1866),
.B2(n_1846),
.C(n_1840),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1886),
.B(n_1758),
.Y(n_1991)
);

BUFx3_ASAP7_75t_L g1992 ( 
.A(n_1959),
.Y(n_1992)
);

NAND4xp25_ASAP7_75t_L g1993 ( 
.A(n_1920),
.B(n_1877),
.C(n_1854),
.D(n_1859),
.Y(n_1993)
);

NAND2xp33_ASAP7_75t_R g1994 ( 
.A(n_1961),
.B(n_1782),
.Y(n_1994)
);

OAI221xp5_ASAP7_75t_L g1995 ( 
.A1(n_1927),
.A2(n_1863),
.B1(n_1855),
.B2(n_1751),
.C(n_1861),
.Y(n_1995)
);

BUFx3_ASAP7_75t_L g1996 ( 
.A(n_1959),
.Y(n_1996)
);

AOI221xp5_ASAP7_75t_L g1997 ( 
.A1(n_1973),
.A2(n_1729),
.B1(n_1748),
.B2(n_1751),
.C(n_1832),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1894),
.Y(n_1998)
);

AOI221xp5_ASAP7_75t_L g1999 ( 
.A1(n_1973),
.A2(n_1968),
.B1(n_1941),
.B2(n_1935),
.C(n_1965),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1900),
.B(n_1790),
.Y(n_2000)
);

BUFx2_ASAP7_75t_L g2001 ( 
.A(n_1962),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1884),
.B(n_1747),
.Y(n_2002)
);

INVxp67_ASAP7_75t_SL g2003 ( 
.A(n_1943),
.Y(n_2003)
);

AOI221xp5_ASAP7_75t_L g2004 ( 
.A1(n_1968),
.A2(n_1747),
.B1(n_1848),
.B2(n_1790),
.C(n_1784),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1915),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1892),
.B(n_1823),
.Y(n_2006)
);

OAI221xp5_ASAP7_75t_L g2007 ( 
.A1(n_1927),
.A2(n_1781),
.B1(n_1823),
.B2(n_1818),
.C(n_1860),
.Y(n_2007)
);

AOI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1960),
.A2(n_1946),
.B1(n_1937),
.B2(n_1933),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1904),
.Y(n_2009)
);

AOI22xp33_ASAP7_75t_L g2010 ( 
.A1(n_1960),
.A2(n_1799),
.B1(n_1814),
.B2(n_1777),
.Y(n_2010)
);

OR2x2_ASAP7_75t_SL g2011 ( 
.A(n_1918),
.B(n_1750),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1913),
.Y(n_2012)
);

AOI221xp5_ASAP7_75t_L g2013 ( 
.A1(n_1941),
.A2(n_1836),
.B1(n_1868),
.B2(n_1831),
.C(n_1777),
.Y(n_2013)
);

OAI221xp5_ASAP7_75t_L g2014 ( 
.A1(n_1930),
.A2(n_1750),
.B1(n_1765),
.B2(n_1785),
.C(n_1975),
.Y(n_2014)
);

AOI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1937),
.A2(n_1785),
.B1(n_1946),
.B2(n_1933),
.Y(n_2015)
);

OAI21x1_ASAP7_75t_L g2016 ( 
.A1(n_1931),
.A2(n_1913),
.B(n_1907),
.Y(n_2016)
);

OA21x2_ASAP7_75t_L g2017 ( 
.A1(n_1944),
.A2(n_1945),
.B(n_1971),
.Y(n_2017)
);

OAI211xp5_ASAP7_75t_SL g2018 ( 
.A1(n_1951),
.A2(n_1953),
.B(n_1972),
.C(n_1897),
.Y(n_2018)
);

INVxp67_ASAP7_75t_L g2019 ( 
.A(n_1895),
.Y(n_2019)
);

AND2x4_ASAP7_75t_L g2020 ( 
.A(n_1906),
.B(n_1888),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_R g2021 ( 
.A(n_1908),
.B(n_1923),
.Y(n_2021)
);

AOI22xp33_ASAP7_75t_SL g2022 ( 
.A1(n_1970),
.A2(n_1967),
.B1(n_1930),
.B2(n_1955),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1913),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1900),
.B(n_1889),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1913),
.Y(n_2025)
);

AOI22xp33_ASAP7_75t_L g2026 ( 
.A1(n_1956),
.A2(n_1958),
.B1(n_1967),
.B2(n_1970),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1890),
.B(n_1974),
.Y(n_2027)
);

OAI31xp33_ASAP7_75t_L g2028 ( 
.A1(n_1956),
.A2(n_1958),
.A3(n_1947),
.B(n_1955),
.Y(n_2028)
);

INVxp67_ASAP7_75t_SL g2029 ( 
.A(n_1934),
.Y(n_2029)
);

OAI211xp5_ASAP7_75t_SL g2030 ( 
.A1(n_1936),
.A2(n_1940),
.B(n_1905),
.C(n_1965),
.Y(n_2030)
);

BUFx2_ASAP7_75t_L g2031 ( 
.A(n_1889),
.Y(n_2031)
);

OA21x2_ASAP7_75t_L g2032 ( 
.A1(n_1944),
.A2(n_1945),
.B(n_1971),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1885),
.B(n_1890),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1885),
.B(n_1929),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_1911),
.Y(n_2035)
);

AOI221xp5_ASAP7_75t_L g2036 ( 
.A1(n_1974),
.A2(n_1942),
.B1(n_1932),
.B2(n_1950),
.C(n_1952),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1901),
.B(n_1903),
.Y(n_2037)
);

NOR2x2_ASAP7_75t_L g2038 ( 
.A(n_1938),
.B(n_1954),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1909),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1983),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_2034),
.B(n_2012),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_2035),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_2003),
.B(n_1950),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_2017),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_2034),
.B(n_1932),
.Y(n_2045)
);

HB1xp67_ASAP7_75t_L g2046 ( 
.A(n_2017),
.Y(n_2046)
);

HB1xp67_ASAP7_75t_L g2047 ( 
.A(n_2017),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_2024),
.B(n_1929),
.Y(n_2048)
);

BUFx2_ASAP7_75t_L g2049 ( 
.A(n_2038),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1979),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2025),
.B(n_1928),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2025),
.B(n_1928),
.Y(n_2052)
);

INVx4_ASAP7_75t_L g2053 ( 
.A(n_1987),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2029),
.B(n_1911),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2025),
.B(n_1925),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2024),
.B(n_1925),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1982),
.B(n_1942),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1986),
.B(n_1998),
.Y(n_2058)
);

INVx1_ASAP7_75t_SL g2059 ( 
.A(n_2001),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_1986),
.B(n_1952),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1979),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1980),
.Y(n_2062)
);

INVx2_ASAP7_75t_SL g2063 ( 
.A(n_1987),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1998),
.B(n_1901),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_2002),
.B(n_1912),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1980),
.Y(n_2066)
);

BUFx2_ASAP7_75t_L g2067 ( 
.A(n_2016),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2017),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2009),
.B(n_1912),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2033),
.B(n_1926),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2033),
.B(n_1926),
.Y(n_2071)
);

HB1xp67_ASAP7_75t_L g2072 ( 
.A(n_2032),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2032),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2023),
.B(n_1987),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_1981),
.B(n_1912),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_1981),
.B(n_1912),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2032),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2031),
.B(n_1907),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2031),
.B(n_1907),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1991),
.B(n_1957),
.Y(n_2080)
);

INVxp67_ASAP7_75t_SL g2081 ( 
.A(n_2005),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1991),
.B(n_1957),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1987),
.B(n_1912),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2023),
.B(n_1912),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_1987),
.B(n_1906),
.Y(n_2085)
);

INVx5_ASAP7_75t_L g2086 ( 
.A(n_1987),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_SL g2087 ( 
.A(n_1988),
.B(n_1948),
.Y(n_2087)
);

OR2x2_ASAP7_75t_L g2088 ( 
.A(n_2027),
.B(n_1921),
.Y(n_2088)
);

INVx4_ASAP7_75t_L g2089 ( 
.A(n_1985),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2032),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2057),
.B(n_2000),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2050),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2049),
.B(n_2001),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2049),
.B(n_1989),
.Y(n_2094)
);

OAI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_2049),
.A2(n_1995),
.B1(n_1993),
.B2(n_1947),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2050),
.Y(n_2096)
);

INVx1_ASAP7_75t_SL g2097 ( 
.A(n_2060),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2070),
.B(n_1989),
.Y(n_2098)
);

NAND4xp25_ASAP7_75t_L g2099 ( 
.A(n_2059),
.B(n_1990),
.C(n_1978),
.D(n_1993),
.Y(n_2099)
);

AND2x4_ASAP7_75t_L g2100 ( 
.A(n_2086),
.B(n_2020),
.Y(n_2100)
);

AOI22xp33_ASAP7_75t_SL g2101 ( 
.A1(n_2089),
.A2(n_1977),
.B1(n_1984),
.B2(n_1917),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2057),
.B(n_2000),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2050),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_2089),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2061),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2061),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_2087),
.A2(n_2022),
.B(n_2018),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_2086),
.B(n_2020),
.Y(n_2108)
);

OR2x2_ASAP7_75t_L g2109 ( 
.A(n_2058),
.B(n_2037),
.Y(n_2109)
);

AND2x4_ASAP7_75t_L g2110 ( 
.A(n_2086),
.B(n_2020),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_2042),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2080),
.B(n_2082),
.Y(n_2112)
);

HB1xp67_ASAP7_75t_L g2113 ( 
.A(n_2042),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2061),
.Y(n_2114)
);

NOR2xp67_ASAP7_75t_L g2115 ( 
.A(n_2086),
.B(n_2089),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_2058),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2070),
.B(n_2019),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2062),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_2043),
.B(n_1985),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_2043),
.B(n_1985),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2089),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_2087),
.B(n_1988),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2062),
.Y(n_2123)
);

INVx1_ASAP7_75t_SL g2124 ( 
.A(n_2060),
.Y(n_2124)
);

INVx2_ASAP7_75t_SL g2125 ( 
.A(n_2086),
.Y(n_2125)
);

AOI322xp5_ASAP7_75t_L g2126 ( 
.A1(n_2045),
.A2(n_2026),
.A3(n_2008),
.B1(n_1999),
.B2(n_1997),
.C1(n_2036),
.C2(n_2004),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2070),
.B(n_1992),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_2080),
.B(n_2030),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2089),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2062),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2080),
.B(n_2082),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2066),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2071),
.B(n_1992),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2082),
.B(n_2006),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2066),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2071),
.B(n_1992),
.Y(n_2136)
);

INVxp67_ASAP7_75t_L g2137 ( 
.A(n_2060),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2054),
.B(n_1985),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2066),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2089),
.Y(n_2140)
);

INVxp67_ASAP7_75t_L g2141 ( 
.A(n_2054),
.Y(n_2141)
);

NOR2xp67_ASAP7_75t_L g2142 ( 
.A(n_2086),
.B(n_2014),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2071),
.B(n_1996),
.Y(n_2143)
);

OAI21xp5_ASAP7_75t_L g2144 ( 
.A1(n_2075),
.A2(n_1976),
.B(n_1919),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2048),
.B(n_2056),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2043),
.B(n_2039),
.Y(n_2146)
);

INVx1_ASAP7_75t_SL g2147 ( 
.A(n_2059),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2040),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2040),
.Y(n_2149)
);

OAI332xp33_ASAP7_75t_L g2150 ( 
.A1(n_2095),
.A2(n_1977),
.A3(n_2076),
.B1(n_2075),
.B2(n_2065),
.B3(n_2073),
.C1(n_2090),
.C2(n_2068),
.Y(n_2150)
);

OR2x4_ASAP7_75t_L g2151 ( 
.A(n_2128),
.B(n_1896),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_2101),
.A2(n_1917),
.B1(n_1994),
.B2(n_2076),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_2099),
.B(n_2011),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2092),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2092),
.Y(n_2155)
);

INVx1_ASAP7_75t_SL g2156 ( 
.A(n_2094),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2096),
.Y(n_2157)
);

BUFx2_ASAP7_75t_L g2158 ( 
.A(n_2094),
.Y(n_2158)
);

INVx5_ASAP7_75t_L g2159 ( 
.A(n_2100),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2145),
.B(n_2056),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_2144),
.B(n_2011),
.Y(n_2161)
);

AOI221xp5_ASAP7_75t_L g2162 ( 
.A1(n_2138),
.A2(n_2076),
.B1(n_2075),
.B2(n_2065),
.C(n_2044),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2134),
.B(n_2045),
.Y(n_2163)
);

NOR2xp67_ASAP7_75t_L g2164 ( 
.A(n_2100),
.B(n_2108),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_L g2165 ( 
.A(n_2137),
.B(n_2045),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2145),
.B(n_2056),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_2111),
.Y(n_2167)
);

INVx2_ASAP7_75t_SL g2168 ( 
.A(n_2100),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2096),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2093),
.B(n_2100),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2103),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2103),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2097),
.B(n_2056),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2093),
.B(n_2048),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2108),
.B(n_2048),
.Y(n_2175)
);

INVx3_ASAP7_75t_L g2176 ( 
.A(n_2108),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2124),
.B(n_2065),
.Y(n_2177)
);

INVxp67_ASAP7_75t_L g2178 ( 
.A(n_2107),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2141),
.B(n_2116),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2105),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2091),
.B(n_2051),
.Y(n_2181)
);

INVx2_ASAP7_75t_SL g2182 ( 
.A(n_2108),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2110),
.B(n_2078),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2112),
.B(n_2088),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2102),
.B(n_2051),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2131),
.B(n_2051),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2105),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_2109),
.B(n_2088),
.Y(n_2188)
);

OR2x2_ASAP7_75t_L g2189 ( 
.A(n_2109),
.B(n_2088),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2110),
.B(n_2078),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2106),
.Y(n_2191)
);

BUFx12f_ASAP7_75t_L g2192 ( 
.A(n_2110),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2110),
.B(n_2078),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2147),
.B(n_2064),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_2098),
.B(n_1922),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2106),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2117),
.B(n_2051),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2114),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2104),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2117),
.B(n_2052),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2113),
.B(n_2052),
.Y(n_2201)
);

NOR3xp33_ASAP7_75t_L g2202 ( 
.A(n_2104),
.B(n_2013),
.C(n_2007),
.Y(n_2202)
);

AND2x4_ASAP7_75t_L g2203 ( 
.A(n_2098),
.B(n_2086),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2178),
.B(n_2126),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2158),
.Y(n_2205)
);

OAI22xp5_ASAP7_75t_L g2206 ( 
.A1(n_2152),
.A2(n_1919),
.B1(n_2122),
.B2(n_2142),
.Y(n_2206)
);

INVx2_ASAP7_75t_SL g2207 ( 
.A(n_2159),
.Y(n_2207)
);

HB1xp67_ASAP7_75t_L g2208 ( 
.A(n_2156),
.Y(n_2208)
);

NOR3xp33_ASAP7_75t_SL g2209 ( 
.A(n_2161),
.B(n_2146),
.C(n_2028),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_2202),
.A2(n_1917),
.B1(n_2120),
.B2(n_2119),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2167),
.Y(n_2211)
);

OR2x2_ASAP7_75t_L g2212 ( 
.A(n_2188),
.B(n_2119),
.Y(n_2212)
);

AOI322xp5_ASAP7_75t_L g2213 ( 
.A1(n_2153),
.A2(n_2015),
.A3(n_2047),
.B1(n_2044),
.B2(n_2072),
.C1(n_2046),
.C2(n_2073),
.Y(n_2213)
);

INVxp67_ASAP7_75t_L g2214 ( 
.A(n_2153),
.Y(n_2214)
);

AOI21xp33_ASAP7_75t_SL g2215 ( 
.A1(n_2161),
.A2(n_2125),
.B(n_2063),
.Y(n_2215)
);

INVx1_ASAP7_75t_SL g2216 ( 
.A(n_2170),
.Y(n_2216)
);

OAI22xp33_ASAP7_75t_L g2217 ( 
.A1(n_2151),
.A2(n_2120),
.B1(n_1969),
.B2(n_2086),
.Y(n_2217)
);

OR2x2_ASAP7_75t_L g2218 ( 
.A(n_2188),
.B(n_2069),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2154),
.Y(n_2219)
);

NOR2xp33_ASAP7_75t_L g2220 ( 
.A(n_2151),
.B(n_2127),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2165),
.B(n_2052),
.Y(n_2221)
);

OAI221xp5_ASAP7_75t_SL g2222 ( 
.A1(n_2162),
.A2(n_2028),
.B1(n_2083),
.B2(n_2084),
.C(n_2067),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2155),
.Y(n_2223)
);

O2A1O1Ixp33_ASAP7_75t_SL g2224 ( 
.A1(n_2179),
.A2(n_2063),
.B(n_2125),
.C(n_2021),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2165),
.B(n_2052),
.Y(n_2225)
);

AOI221xp5_ASAP7_75t_L g2226 ( 
.A1(n_2150),
.A2(n_2047),
.B1(n_2072),
.B2(n_2046),
.C(n_2077),
.Y(n_2226)
);

OAI22xp5_ASAP7_75t_L g2227 ( 
.A1(n_2195),
.A2(n_2142),
.B1(n_1961),
.B2(n_2143),
.Y(n_2227)
);

AOI221xp5_ASAP7_75t_L g2228 ( 
.A1(n_2177),
.A2(n_2077),
.B1(n_2068),
.B2(n_2073),
.C(n_2090),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2170),
.B(n_2174),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2189),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2157),
.Y(n_2231)
);

INVxp67_ASAP7_75t_L g2232 ( 
.A(n_2195),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2169),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2171),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2172),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2180),
.Y(n_2236)
);

OAI32xp33_ASAP7_75t_L g2237 ( 
.A1(n_2189),
.A2(n_2084),
.A3(n_2083),
.B1(n_2140),
.B2(n_2121),
.Y(n_2237)
);

INVxp67_ASAP7_75t_L g2238 ( 
.A(n_2194),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2187),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2191),
.Y(n_2240)
);

INVx2_ASAP7_75t_SL g2241 ( 
.A(n_2159),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2163),
.B(n_2055),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2184),
.B(n_2055),
.Y(n_2243)
);

AOI22x1_ASAP7_75t_L g2244 ( 
.A1(n_2192),
.A2(n_2140),
.B1(n_2129),
.B2(n_2121),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2196),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_2199),
.Y(n_2246)
);

AOI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_2204),
.A2(n_2083),
.B1(n_1917),
.B2(n_1949),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2212),
.Y(n_2248)
);

XOR2x2_ASAP7_75t_L g2249 ( 
.A(n_2222),
.B(n_2173),
.Y(n_2249)
);

AOI211xp5_ASAP7_75t_SL g2250 ( 
.A1(n_2224),
.A2(n_2164),
.B(n_2176),
.C(n_2115),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2232),
.B(n_2174),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2219),
.Y(n_2252)
);

AOI222xp33_ASAP7_75t_L g2253 ( 
.A1(n_2214),
.A2(n_2068),
.B1(n_2077),
.B2(n_2090),
.C1(n_2069),
.C2(n_1963),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2223),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2229),
.B(n_2175),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2230),
.B(n_2160),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2230),
.B(n_2208),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2231),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_L g2259 ( 
.A(n_2216),
.B(n_2192),
.Y(n_2259)
);

NAND2xp33_ASAP7_75t_SL g2260 ( 
.A(n_2205),
.B(n_2168),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2205),
.B(n_2160),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2233),
.Y(n_2262)
);

O2A1O1Ixp33_ASAP7_75t_L g2263 ( 
.A1(n_2209),
.A2(n_2129),
.B(n_2201),
.C(n_2067),
.Y(n_2263)
);

NOR4xp25_ASAP7_75t_L g2264 ( 
.A(n_2211),
.B(n_2199),
.C(n_2182),
.D(n_2168),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2238),
.B(n_2166),
.Y(n_2265)
);

AOI221x1_ASAP7_75t_SL g2266 ( 
.A1(n_2217),
.A2(n_2198),
.B1(n_2200),
.B2(n_2197),
.C(n_2203),
.Y(n_2266)
);

AND2x4_ASAP7_75t_L g2267 ( 
.A(n_2229),
.B(n_2159),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_2220),
.B(n_2159),
.Y(n_2268)
);

OAI22xp33_ASAP7_75t_L g2269 ( 
.A1(n_2210),
.A2(n_1969),
.B1(n_2086),
.B2(n_2053),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2234),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2220),
.B(n_2175),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2235),
.Y(n_2272)
);

BUFx2_ASAP7_75t_L g2273 ( 
.A(n_2207),
.Y(n_2273)
);

INVx3_ASAP7_75t_L g2274 ( 
.A(n_2207),
.Y(n_2274)
);

INVxp67_ASAP7_75t_L g2275 ( 
.A(n_2241),
.Y(n_2275)
);

AOI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_2227),
.A2(n_1949),
.B1(n_2085),
.B2(n_1963),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2213),
.B(n_2166),
.Y(n_2277)
);

NOR3xp33_ASAP7_75t_SL g2278 ( 
.A(n_2260),
.B(n_2217),
.C(n_2237),
.Y(n_2278)
);

NOR3xp33_ASAP7_75t_SL g2279 ( 
.A(n_2260),
.B(n_2206),
.C(n_2226),
.Y(n_2279)
);

OAI22xp33_ASAP7_75t_L g2280 ( 
.A1(n_2277),
.A2(n_2212),
.B1(n_2241),
.B2(n_2221),
.Y(n_2280)
);

NAND2x1_ASAP7_75t_L g2281 ( 
.A(n_2267),
.B(n_2176),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2257),
.Y(n_2282)
);

OR2x2_ASAP7_75t_L g2283 ( 
.A(n_2256),
.B(n_2225),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2248),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2251),
.B(n_2236),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2248),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2265),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2252),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2254),
.Y(n_2289)
);

NOR2x1_ASAP7_75t_L g2290 ( 
.A(n_2274),
.B(n_2239),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2258),
.Y(n_2291)
);

NOR4xp25_ASAP7_75t_SL g2292 ( 
.A(n_2273),
.B(n_2224),
.C(n_2215),
.D(n_2228),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2262),
.Y(n_2293)
);

INVxp67_ASAP7_75t_SL g2294 ( 
.A(n_2274),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2270),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2259),
.B(n_2275),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2255),
.B(n_2271),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2264),
.B(n_2240),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2272),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2261),
.B(n_2245),
.Y(n_2300)
);

INVxp67_ASAP7_75t_SL g2301 ( 
.A(n_2294),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2294),
.Y(n_2302)
);

AOI21xp5_ASAP7_75t_L g2303 ( 
.A1(n_2292),
.A2(n_2263),
.B(n_2249),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2284),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2297),
.B(n_2259),
.Y(n_2305)
);

OAI221xp5_ASAP7_75t_L g2306 ( 
.A1(n_2279),
.A2(n_2266),
.B1(n_2249),
.B2(n_2247),
.C(n_2276),
.Y(n_2306)
);

NAND3xp33_ASAP7_75t_SL g2307 ( 
.A(n_2298),
.B(n_2253),
.C(n_2268),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2286),
.Y(n_2308)
);

OAI22xp33_ASAP7_75t_L g2309 ( 
.A1(n_2280),
.A2(n_2269),
.B1(n_2250),
.B2(n_2159),
.Y(n_2309)
);

O2A1O1Ixp5_ASAP7_75t_SL g2310 ( 
.A1(n_2282),
.A2(n_2274),
.B(n_2176),
.C(n_2268),
.Y(n_2310)
);

AOI211xp5_ASAP7_75t_L g2311 ( 
.A1(n_2280),
.A2(n_2269),
.B(n_2296),
.C(n_2300),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2285),
.Y(n_2312)
);

OAI22xp5_ASAP7_75t_L g2313 ( 
.A1(n_2278),
.A2(n_2267),
.B1(n_2203),
.B2(n_2182),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_L g2314 ( 
.A(n_2283),
.B(n_2267),
.Y(n_2314)
);

AOI211xp5_ASAP7_75t_L g2315 ( 
.A1(n_2287),
.A2(n_2246),
.B(n_2218),
.C(n_2084),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2302),
.Y(n_2316)
);

NAND4xp25_ASAP7_75t_L g2317 ( 
.A(n_2303),
.B(n_2290),
.C(n_2295),
.D(n_2293),
.Y(n_2317)
);

AOI221x1_ASAP7_75t_L g2318 ( 
.A1(n_2307),
.A2(n_2304),
.B1(n_2308),
.B2(n_2305),
.C(n_2312),
.Y(n_2318)
);

AO221x1_ASAP7_75t_L g2319 ( 
.A1(n_2309),
.A2(n_2299),
.B1(n_2291),
.B2(n_2289),
.C(n_2288),
.Y(n_2319)
);

NAND4xp25_ASAP7_75t_L g2320 ( 
.A(n_2311),
.B(n_2279),
.C(n_2278),
.D(n_2203),
.Y(n_2320)
);

NAND4xp25_ASAP7_75t_L g2321 ( 
.A(n_2314),
.B(n_2307),
.C(n_2306),
.D(n_2313),
.Y(n_2321)
);

A2O1A1Ixp33_ASAP7_75t_L g2322 ( 
.A1(n_2301),
.A2(n_2315),
.B(n_2246),
.C(n_2281),
.Y(n_2322)
);

NOR2x1_ASAP7_75t_SL g2323 ( 
.A(n_2310),
.B(n_2183),
.Y(n_2323)
);

OAI21xp5_ASAP7_75t_SL g2324 ( 
.A1(n_2303),
.A2(n_2190),
.B(n_2183),
.Y(n_2324)
);

AOI211xp5_ASAP7_75t_L g2325 ( 
.A1(n_2303),
.A2(n_2218),
.B(n_2084),
.C(n_2243),
.Y(n_2325)
);

AOI211xp5_ASAP7_75t_L g2326 ( 
.A1(n_2303),
.A2(n_2067),
.B(n_2193),
.C(n_2190),
.Y(n_2326)
);

AOI211x1_ASAP7_75t_SL g2327 ( 
.A1(n_2307),
.A2(n_2242),
.B(n_2244),
.C(n_2181),
.Y(n_2327)
);

AOI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2307),
.A2(n_2085),
.B1(n_2185),
.B2(n_2193),
.Y(n_2328)
);

NAND3xp33_ASAP7_75t_SL g2329 ( 
.A(n_2303),
.B(n_2074),
.C(n_2136),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_2320),
.B(n_2114),
.Y(n_2330)
);

NAND4xp25_ASAP7_75t_SL g2331 ( 
.A(n_2318),
.B(n_2143),
.C(n_2136),
.D(n_2127),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2316),
.Y(n_2332)
);

AOI222xp33_ASAP7_75t_L g2333 ( 
.A1(n_2329),
.A2(n_1964),
.B1(n_2081),
.B2(n_1916),
.C1(n_2055),
.C2(n_1966),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2327),
.B(n_2186),
.Y(n_2334)
);

OAI211xp5_ASAP7_75t_L g2335 ( 
.A1(n_2317),
.A2(n_2053),
.B(n_2086),
.C(n_2063),
.Y(n_2335)
);

INVx1_ASAP7_75t_SL g2336 ( 
.A(n_2328),
.Y(n_2336)
);

OAI321xp33_ASAP7_75t_L g2337 ( 
.A1(n_2321),
.A2(n_2325),
.A3(n_2326),
.B1(n_2322),
.B2(n_2319),
.C(n_2323),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_R g2338 ( 
.A(n_2324),
.B(n_2133),
.Y(n_2338)
);

NOR2xp67_ASAP7_75t_L g2339 ( 
.A(n_2331),
.B(n_2335),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2332),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_2336),
.Y(n_2341)
);

BUFx2_ASAP7_75t_L g2342 ( 
.A(n_2338),
.Y(n_2342)
);

NOR2x1p5_ASAP7_75t_L g2343 ( 
.A(n_2334),
.B(n_2053),
.Y(n_2343)
);

NAND2x1p5_ASAP7_75t_L g2344 ( 
.A(n_2330),
.B(n_2053),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2333),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2337),
.Y(n_2346)
);

AND2x4_ASAP7_75t_L g2347 ( 
.A(n_2332),
.B(n_2133),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2347),
.B(n_2041),
.Y(n_2348)
);

OAI21xp33_ASAP7_75t_SL g2349 ( 
.A1(n_2346),
.A2(n_2339),
.B(n_2343),
.Y(n_2349)
);

NOR3xp33_ASAP7_75t_L g2350 ( 
.A(n_2341),
.B(n_2053),
.C(n_2063),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2341),
.B(n_2118),
.Y(n_2351)
);

OAI22x1_ASAP7_75t_L g2352 ( 
.A1(n_2342),
.A2(n_2340),
.B1(n_2345),
.B2(n_2347),
.Y(n_2352)
);

NAND3xp33_ASAP7_75t_SL g2353 ( 
.A(n_2340),
.B(n_2010),
.C(n_1924),
.Y(n_2353)
);

OAI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2344),
.A2(n_2149),
.B1(n_2148),
.B2(n_2139),
.Y(n_2354)
);

XOR2x2_ASAP7_75t_L g2355 ( 
.A(n_2351),
.B(n_2344),
.Y(n_2355)
);

CKINVDCx5p33_ASAP7_75t_R g2356 ( 
.A(n_2352),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2348),
.Y(n_2357)
);

INVx3_ASAP7_75t_L g2358 ( 
.A(n_2350),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2356),
.Y(n_2359)
);

AOI221xp5_ASAP7_75t_L g2360 ( 
.A1(n_2359),
.A2(n_2356),
.B1(n_2349),
.B2(n_2357),
.C(n_2358),
.Y(n_2360)
);

INVx1_ASAP7_75t_SL g2361 ( 
.A(n_2360),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2360),
.Y(n_2362)
);

AOI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_2361),
.A2(n_2355),
.B(n_2358),
.Y(n_2363)
);

AOI21xp5_ASAP7_75t_L g2364 ( 
.A1(n_2362),
.A2(n_2354),
.B(n_2353),
.Y(n_2364)
);

AOI222xp33_ASAP7_75t_L g2365 ( 
.A1(n_2363),
.A2(n_2149),
.B1(n_2148),
.B2(n_2139),
.C1(n_2135),
.C2(n_2132),
.Y(n_2365)
);

AOI22xp33_ASAP7_75t_SL g2366 ( 
.A1(n_2364),
.A2(n_2053),
.B1(n_2085),
.B2(n_2130),
.Y(n_2366)
);

AOI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_2366),
.A2(n_2135),
.B1(n_2132),
.B2(n_2130),
.Y(n_2367)
);

OAI221xp5_ASAP7_75t_R g2368 ( 
.A1(n_2367),
.A2(n_2365),
.B1(n_1938),
.B2(n_2118),
.C(n_2123),
.Y(n_2368)
);

AOI211xp5_ASAP7_75t_L g2369 ( 
.A1(n_2368),
.A2(n_2123),
.B(n_2079),
.C(n_2085),
.Y(n_2369)
);


endmodule