module fake_jpeg_22988_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_SL g10 ( 
.A(n_4),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

OR2x4_ASAP7_75t_L g14 ( 
.A(n_12),
.B(n_0),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_14),
.A2(n_10),
.B(n_9),
.Y(n_25)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_18),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_8),
.B(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_17),
.Y(n_26)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_11),
.B1(n_12),
.B2(n_3),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_19),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_18),
.B1(n_15),
.B2(n_9),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_17),
.B1(n_7),
.B2(n_3),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_28),
.B1(n_12),
.B2(n_7),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2x1_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_40),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_29),
.B(n_26),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_34),
.B(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_22),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_34),
.A3(n_31),
.B1(n_32),
.B2(n_24),
.C1(n_27),
.C2(n_5),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_42),
.Y(n_44)
);


endmodule