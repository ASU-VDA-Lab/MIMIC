module real_jpeg_30719_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_0),
.Y(n_112)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_0),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_43),
.Y(n_42)
);

AND2x4_ASAP7_75t_L g58 ( 
.A(n_1),
.B(n_59),
.Y(n_58)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_1),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_1),
.B(n_112),
.Y(n_111)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_1),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_1),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_1),
.B(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_1),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_2),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_2),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_2),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_2),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_2),
.B(n_116),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_19),
.B(n_454),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_3),
.B(n_455),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_4),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_5),
.Y(n_118)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_6),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_7),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_7),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_7),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_7),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_7),
.B(n_273),
.Y(n_272)
);

NAND2x1_ASAP7_75t_L g443 ( 
.A(n_7),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_8),
.B(n_47),
.Y(n_46)
);

NAND2x1_ASAP7_75t_L g138 ( 
.A(n_8),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_8),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_8),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_8),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_8),
.B(n_279),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_8),
.B(n_282),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_8),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_9),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_9),
.B(n_116),
.Y(n_115)
);

NAND2x1_ASAP7_75t_SL g142 ( 
.A(n_9),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_9),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_9),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g435 ( 
.A(n_9),
.B(n_105),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_10),
.Y(n_179)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_11),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_12),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_12),
.B(n_248),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_SL g320 ( 
.A(n_12),
.B(n_321),
.Y(n_320)
);

NAND2x1_ASAP7_75t_L g333 ( 
.A(n_12),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_12),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_12),
.B(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_13),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_14),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_14),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_14),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_14),
.B(n_266),
.Y(n_265)
);

AND2x4_ASAP7_75t_SL g317 ( 
.A(n_14),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_14),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_14),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_14),
.B(n_358),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_15),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_16),
.Y(n_131)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_16),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_16),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_64),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_17),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_17),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_17),
.B(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_17),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_17),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_17),
.B(n_347),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_414),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_233),
.B(n_412),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_182),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_24),
.B(n_183),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_107),
.C(n_146),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_25),
.B(n_408),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_74),
.C(n_89),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_26),
.B(n_401),
.Y(n_400)
);

OAI21x1_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_55),
.B(n_73),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_39),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_28),
.B(n_39),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_28),
.A2(n_29),
.B1(n_39),
.B2(n_40),
.Y(n_299)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_30),
.B(n_34),
.Y(n_245)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_34),
.A2(n_35),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_35),
.B(n_111),
.C(n_115),
.Y(n_202)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_38),
.Y(n_136)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_46),
.C(n_51),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_41),
.A2(n_42),
.B1(n_51),
.B2(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_41),
.B(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_44),
.Y(n_318)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_44),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_45),
.Y(n_286)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_46),
.Y(n_241)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_49),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_50),
.Y(n_255)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_51),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_54),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_54),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_54),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_55),
.B(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_68),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_58),
.B(n_63),
.C(n_68),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g398 ( 
.A(n_58),
.B(n_63),
.C(n_68),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_71),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_72),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_74),
.B(n_89),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_85),
.B2(n_86),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_84),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_78),
.B(n_82),
.C(n_86),
.Y(n_172)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_81),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_82),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_82),
.B(n_217),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_82),
.A2(n_84),
.B1(n_216),
.B2(n_217),
.Y(n_287)
);

INVx4_ASAP7_75t_SL g316 ( 
.A(n_83),
.Y(n_316)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_99),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_90),
.A2(n_92),
.B(n_95),
.Y(n_291)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_94),
.Y(n_348)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_98),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_103),
.B(n_106),
.C(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_108),
.B(n_147),
.Y(n_408)
);

XNOR2x1_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_109),
.B(n_120),
.C(n_145),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_111),
.A2(n_113),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_111),
.B(n_278),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_111),
.B(n_155),
.C(n_209),
.Y(n_446)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_112),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_113),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_118),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_132),
.B1(n_144),
.B2(n_145),
.Y(n_119)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_122),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_126),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_128),
.B(n_213),
.C(n_214),
.Y(n_212)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.C(n_140),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_150),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx4f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_136),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_141),
.B1(n_142),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_141),
.A2(n_142),
.B1(n_433),
.B2(n_434),
.Y(n_432)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_168),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_148),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_153),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_149),
.B(n_153),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.C(n_163),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_154),
.B(n_164),
.Y(n_293)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2x2_ASAP7_75t_L g206 ( 
.A(n_155),
.B(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_158),
.B(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_172),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_176),
.B1(n_180),
.B2(n_181),
.Y(n_173)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_178),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_190),
.C(n_191),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_203),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_184),
.B(n_228),
.C(n_452),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_185),
.B(n_189),
.C(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_192),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_202),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_199),
.B2(n_201),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_194),
.B(n_201),
.C(n_202),
.Y(n_448)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_199),
.B(n_443),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_228),
.B2(n_232),
.Y(n_203)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_204),
.Y(n_452)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_206),
.B(n_212),
.C(n_215),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_216),
.A2(n_217),
.B1(n_424),
.B2(n_425),
.Y(n_423)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_217),
.B(n_225),
.C(n_437),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_219),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.Y(n_220)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_221),
.Y(n_437)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.C(n_231),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_390),
.B(n_409),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_304),
.B(n_389),
.Y(n_235)
);

NOR2xp67_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_288),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_237),
.B(n_288),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_261),
.C(n_276),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_238),
.B(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_244),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_240),
.B(n_245),
.C(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_252),
.C(n_256),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g302 ( 
.A(n_247),
.B(n_252),
.C(n_256),
.Y(n_302)
);

XNOR2x1_ASAP7_75t_L g379 ( 
.A(n_247),
.B(n_256),
.Y(n_379)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_251),
.Y(n_444)
);

XNOR2x1_ASAP7_75t_L g378 ( 
.A(n_252),
.B(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_261),
.A2(n_262),
.B1(n_276),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_271),
.C(n_275),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_271),
.B1(n_272),
.B2(n_275),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_276),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_281),
.C(n_287),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_277),
.B(n_281),
.Y(n_381)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_287),
.B(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_297),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_289),
.B(n_300),
.C(n_393),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_296),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_290)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_291),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_292),
.B(n_294),
.C(n_296),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_300),
.B1(n_301),
.B2(n_303),
.Y(n_297)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_298),
.Y(n_393)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_383),
.B(n_388),
.Y(n_304)
);

OAI21x1_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_371),
.B(n_382),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_339),
.B(n_370),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_323),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_308),
.B(n_323),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_317),
.C(n_319),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_309),
.A2(n_310),
.B1(n_366),
.B2(n_367),
.Y(n_365)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_314),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_314),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_317),
.A2(n_319),
.B1(n_320),
.B2(n_368),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_317),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_318),
.Y(n_338)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_329),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_325),
.B(n_328),
.C(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_332),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_330),
.B(n_333),
.C(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_337),
.Y(n_332)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_337),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_363),
.B(n_369),
.Y(n_339)
);

AOI21xp33_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_352),
.B(n_362),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_349),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_342),
.B(n_349),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_346),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_346),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_357),
.Y(n_352)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_364),
.B(n_365),
.Y(n_369)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_374),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_374),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_380),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_376),
.B(n_378),
.C(n_380),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_384),
.B(n_387),
.Y(n_388)
);

NOR2x1_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_402),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_394),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_400),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_396),
.B(n_405),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_405),
.Y(n_406)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_397),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

AO21x1_ASAP7_75t_L g403 ( 
.A1(n_400),
.A2(n_404),
.B(n_406),
.Y(n_403)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_402),
.A2(n_410),
.B(n_411),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_407),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_403),
.B(n_407),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_453),
.Y(n_414)
);

INVxp33_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_450),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_450),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_439),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_429),
.Y(n_421)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx6_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_431),
.B1(n_436),
.B2(n_438),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_431),
.Y(n_430)
);

XOR2x2_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_435),
.Y(n_431)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_433),
.Y(n_434)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_436),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_449),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_448),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_445),
.B1(n_446),
.B2(n_447),
.Y(n_441)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_442),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);


endmodule