module real_aes_381_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_231;
wire n_547;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_0), .A2(n_193), .B1(n_408), .B2(n_409), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_1), .A2(n_80), .B1(n_273), .B2(n_279), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_2), .A2(n_194), .B1(n_418), .B2(n_422), .Y(n_481) );
AO22x2_ASAP7_75t_L g259 ( .A1(n_3), .A2(n_155), .B1(n_249), .B2(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g596 ( .A(n_3), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_4), .A2(n_91), .B1(n_323), .B2(n_359), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_5), .A2(n_159), .B1(n_516), .B2(n_517), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_6), .A2(n_129), .B1(n_373), .B2(n_374), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_7), .A2(n_191), .B1(n_387), .B2(n_389), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_8), .A2(n_47), .B1(n_557), .B2(n_558), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_9), .A2(n_101), .B1(n_263), .B2(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_10), .A2(n_214), .B1(n_419), .B2(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_11), .A2(n_78), .B1(n_262), .B2(n_270), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_12), .A2(n_49), .B1(n_421), .B2(n_422), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_13), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_14), .A2(n_40), .B1(n_389), .B2(n_514), .Y(n_513) );
AO22x2_ASAP7_75t_L g256 ( .A1(n_15), .A2(n_46), .B1(n_249), .B2(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_15), .B(n_595), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_16), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_17), .A2(n_36), .B1(n_418), .B2(n_419), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_18), .A2(n_125), .B1(n_421), .B2(n_422), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_19), .A2(n_184), .B1(n_414), .B2(n_415), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_20), .A2(n_108), .B1(n_322), .B2(n_380), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_21), .A2(n_41), .B1(n_285), .B2(n_292), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_22), .A2(n_75), .B1(n_303), .B2(n_392), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_23), .A2(n_168), .B1(n_349), .B2(n_350), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_24), .A2(n_43), .B1(n_352), .B2(n_353), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_25), .A2(n_63), .B1(n_392), .B2(n_444), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_26), .A2(n_174), .B1(n_349), .B2(n_350), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_27), .A2(n_221), .B1(n_418), .B2(n_422), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_28), .A2(n_122), .B1(n_418), .B2(n_422), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_29), .A2(n_197), .B1(n_418), .B2(n_419), .Y(n_417) );
AO22x1_ASAP7_75t_L g534 ( .A1(n_30), .A2(n_160), .B1(n_353), .B2(n_535), .Y(n_534) );
OA22x2_ASAP7_75t_L g525 ( .A1(n_31), .A2(n_526), .B1(n_527), .B2(n_548), .Y(n_525) );
INVx1_ASAP7_75t_L g548 ( .A(n_31), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_32), .A2(n_133), .B1(n_341), .B2(n_342), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_33), .A2(n_92), .B1(n_408), .B2(n_409), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_34), .A2(n_145), .B1(n_405), .B2(n_435), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_35), .A2(n_82), .B1(n_355), .B2(n_356), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_37), .A2(n_173), .B1(n_462), .B2(n_463), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_38), .A2(n_99), .B1(n_356), .B2(n_383), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_39), .A2(n_51), .B1(n_313), .B2(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_42), .A2(n_103), .B1(n_318), .B2(n_415), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_44), .A2(n_62), .B1(n_399), .B2(n_400), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_45), .A2(n_74), .B1(n_312), .B2(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_48), .A2(n_93), .B1(n_409), .B2(n_492), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_50), .A2(n_111), .B1(n_399), .B2(n_490), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_52), .A2(n_150), .B1(n_460), .B2(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_53), .A2(n_210), .B1(n_399), .B2(n_400), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_54), .A2(n_115), .B1(n_373), .B2(n_546), .Y(n_545) );
OA22x2_ASAP7_75t_L g622 ( .A1(n_55), .A2(n_623), .B1(n_624), .B2(n_647), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_55), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_56), .A2(n_81), .B1(n_344), .B2(n_345), .Y(n_343) );
INVx3_ASAP7_75t_L g249 ( .A(n_57), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_58), .A2(n_127), .B1(n_345), .B2(n_460), .Y(n_459) );
AO22x2_ASAP7_75t_L g456 ( .A1(n_59), .A2(n_457), .B1(n_473), .B2(n_474), .Y(n_456) );
INVx1_ASAP7_75t_L g473 ( .A(n_59), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_60), .A2(n_71), .B1(n_262), .B2(n_268), .Y(n_261) );
XOR2x1_ASAP7_75t_L g363 ( .A(n_61), .B(n_364), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_64), .A2(n_141), .B1(n_367), .B2(n_370), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_65), .A2(n_113), .B1(n_300), .B2(n_303), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_66), .A2(n_132), .B1(n_316), .B2(n_321), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_67), .A2(n_217), .B1(n_387), .B2(n_389), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_68), .A2(n_143), .B1(n_415), .B2(n_484), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_69), .B(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_70), .B(n_560), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_72), .A2(n_207), .B1(n_350), .B2(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g250 ( .A(n_73), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_73), .B(n_98), .Y(n_597) );
INVx2_ASAP7_75t_L g229 ( .A(n_76), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_77), .A2(n_112), .B1(n_380), .B2(n_381), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_79), .A2(n_220), .B1(n_414), .B2(n_415), .Y(n_413) );
XOR2x2_ASAP7_75t_L g498 ( .A(n_83), .B(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_84), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_85), .A2(n_105), .B1(n_367), .B2(n_553), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_86), .A2(n_96), .B1(n_385), .B2(n_422), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_87), .A2(n_177), .B1(n_352), .B2(n_353), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_88), .B(n_377), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_89), .A2(n_123), .B1(n_300), .B2(n_321), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_90), .A2(n_106), .B1(n_316), .B2(n_566), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_94), .A2(n_202), .B1(n_405), .B2(n_435), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_95), .A2(n_190), .B1(n_415), .B2(n_484), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_97), .B(n_402), .Y(n_577) );
AO22x2_ASAP7_75t_L g252 ( .A1(n_98), .A2(n_161), .B1(n_249), .B2(n_253), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_100), .A2(n_158), .B1(n_339), .B2(n_375), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_102), .B(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_104), .A2(n_186), .B1(n_287), .B2(n_367), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_107), .A2(n_185), .B1(n_399), .B2(n_400), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_109), .A2(n_179), .B1(n_370), .B2(n_371), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_110), .B(n_377), .Y(n_465) );
AO22x1_ASAP7_75t_L g532 ( .A1(n_114), .A2(n_149), .B1(n_360), .B2(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_116), .Y(n_431) );
AO22x1_ASAP7_75t_L g536 ( .A1(n_117), .A2(n_153), .B1(n_318), .B2(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g251 ( .A(n_118), .Y(n_251) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_119), .A2(n_170), .B1(n_350), .B2(n_440), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_120), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_121), .A2(n_138), .B1(n_322), .B2(n_468), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_124), .A2(n_148), .B1(n_349), .B2(n_350), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_126), .A2(n_196), .B1(n_287), .B2(n_435), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_128), .B(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_130), .A2(n_188), .B1(n_323), .B2(n_359), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g434 ( .A1(n_131), .A2(n_216), .B1(n_405), .B2(n_435), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_134), .A2(n_154), .B1(n_349), .B2(n_350), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_135), .A2(n_164), .B1(n_349), .B2(n_350), .Y(n_412) );
INVx1_ASAP7_75t_L g238 ( .A(n_136), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_137), .A2(n_211), .B1(n_375), .B2(n_506), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_139), .A2(n_147), .B1(n_511), .B2(n_512), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_140), .A2(n_187), .B1(n_328), .B2(n_383), .Y(n_563) );
XNOR2x1_ASAP7_75t_L g574 ( .A(n_142), .B(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_144), .A2(n_166), .B1(n_359), .B2(n_360), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_146), .A2(n_175), .B1(n_405), .B2(n_406), .Y(n_404) );
AOI21xp5_ASAP7_75t_SL g539 ( .A1(n_151), .A2(n_540), .B(n_541), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_152), .A2(n_212), .B1(n_325), .B2(n_328), .Y(n_324) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_156), .A2(n_204), .B1(n_506), .B2(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g423 ( .A(n_157), .Y(n_423) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_162), .A2(n_223), .B(n_232), .C(n_598), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_163), .A2(n_172), .B1(n_303), .B2(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_165), .A2(n_203), .B1(n_399), .B2(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_167), .B(n_488), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_169), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_171), .B(n_242), .Y(n_508) );
XOR2x2_ASAP7_75t_L g549 ( .A(n_176), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_178), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g592 ( .A(n_178), .Y(n_592) );
AO22x2_ASAP7_75t_L g478 ( .A1(n_180), .A2(n_479), .B1(n_495), .B2(n_496), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_180), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_181), .A2(n_600), .B1(n_614), .B2(n_615), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_181), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_182), .A2(n_205), .B1(n_408), .B2(n_493), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_183), .A2(n_213), .B1(n_279), .B2(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g226 ( .A(n_189), .Y(n_226) );
AND2x2_ASAP7_75t_R g617 ( .A(n_189), .B(n_592), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_192), .B(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_195), .A2(n_208), .B1(n_307), .B2(n_312), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_198), .B(n_242), .Y(n_241) );
INVxp67_ASAP7_75t_L g231 ( .A(n_199), .Y(n_231) );
XNOR2x1_ASAP7_75t_L g333 ( .A(n_200), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g446 ( .A(n_201), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_206), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_209), .A2(n_215), .B1(n_418), .B2(n_422), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_218), .A2(n_219), .B1(n_492), .B2(n_493), .Y(n_491) );
BUFx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2x1_ASAP7_75t_R g224 ( .A(n_225), .B(n_227), .Y(n_224) );
OR2x2_ASAP7_75t_L g653 ( .A(n_225), .B(n_228), .Y(n_653) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_226), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_451), .B1(n_587), .B2(n_588), .C(n_589), .Y(n_232) );
INVx1_ASAP7_75t_L g588 ( .A(n_233), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B1(n_362), .B2(n_450), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OAI22xp5_ASAP7_75t_SL g235 ( .A1(n_236), .A2(n_237), .B1(n_331), .B2(n_361), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
XNOR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
NOR2x1_ASAP7_75t_L g239 ( .A(n_240), .B(n_298), .Y(n_239) );
NAND4xp25_ASAP7_75t_SL g240 ( .A(n_241), .B(n_261), .C(n_272), .D(n_284), .Y(n_240) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g561 ( .A(n_243), .Y(n_561) );
INVx3_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
INVx4_ASAP7_75t_SL g337 ( .A(n_244), .Y(n_337) );
INVx3_ASAP7_75t_L g377 ( .A(n_244), .Y(n_377) );
INVx4_ASAP7_75t_SL g488 ( .A(n_244), .Y(n_488) );
INVx6_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_254), .Y(n_245) );
AND2x4_ASAP7_75t_L g270 ( .A(n_246), .B(n_271), .Y(n_270) );
AND2x4_ASAP7_75t_L g295 ( .A(n_246), .B(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g402 ( .A(n_246), .B(n_254), .Y(n_402) );
AND2x2_ASAP7_75t_L g406 ( .A(n_246), .B(n_296), .Y(n_406) );
AND2x2_ASAP7_75t_L g409 ( .A(n_246), .B(n_271), .Y(n_409) );
AND2x2_ASAP7_75t_L g435 ( .A(n_246), .B(n_296), .Y(n_435) );
AND2x2_ASAP7_75t_L g493 ( .A(n_246), .B(n_271), .Y(n_493) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_252), .Y(n_246) );
INVx2_ASAP7_75t_L g267 ( .A(n_247), .Y(n_267) );
AND2x2_ASAP7_75t_L g277 ( .A(n_247), .B(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_247), .Y(n_283) );
OAI22x1_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B1(n_250), .B2(n_251), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g253 ( .A(n_249), .Y(n_253) );
INVx2_ASAP7_75t_L g257 ( .A(n_249), .Y(n_257) );
INVx1_ASAP7_75t_L g260 ( .A(n_249), .Y(n_260) );
AND2x2_ASAP7_75t_L g266 ( .A(n_252), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g278 ( .A(n_252), .Y(n_278) );
BUFx2_ASAP7_75t_L g314 ( .A(n_252), .Y(n_314) );
AND2x4_ASAP7_75t_L g302 ( .A(n_254), .B(n_277), .Y(n_302) );
AND2x4_ASAP7_75t_L g320 ( .A(n_254), .B(n_305), .Y(n_320) );
AND2x2_ASAP7_75t_L g327 ( .A(n_254), .B(n_266), .Y(n_327) );
AND2x2_ASAP7_75t_L g414 ( .A(n_254), .B(n_277), .Y(n_414) );
AND2x6_ASAP7_75t_L g418 ( .A(n_254), .B(n_266), .Y(n_418) );
AND2x2_ASAP7_75t_L g421 ( .A(n_254), .B(n_305), .Y(n_421) );
AND2x2_ASAP7_75t_L g484 ( .A(n_254), .B(n_277), .Y(n_484) );
AND2x4_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x4_ASAP7_75t_L g265 ( .A(n_256), .B(n_258), .Y(n_265) );
AND2x2_ASAP7_75t_L g282 ( .A(n_256), .B(n_259), .Y(n_282) );
INVx1_ASAP7_75t_L g291 ( .A(n_256), .Y(n_291) );
INVxp67_ASAP7_75t_L g271 ( .A(n_258), .Y(n_271) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g290 ( .A(n_259), .B(n_291), .Y(n_290) );
BUFx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_L g370 ( .A(n_263), .Y(n_370) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
BUFx2_ASAP7_75t_L g341 ( .A(n_264), .Y(n_341) );
BUFx3_ASAP7_75t_L g462 ( .A(n_264), .Y(n_462) );
AND2x4_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x2_ASAP7_75t_L g276 ( .A(n_265), .B(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g323 ( .A(n_265), .B(n_305), .Y(n_323) );
AND2x4_ASAP7_75t_L g399 ( .A(n_265), .B(n_277), .Y(n_399) );
AND2x2_ASAP7_75t_L g408 ( .A(n_265), .B(n_266), .Y(n_408) );
AND2x2_ASAP7_75t_L g419 ( .A(n_265), .B(n_305), .Y(n_419) );
AND2x2_ASAP7_75t_L g492 ( .A(n_265), .B(n_266), .Y(n_492) );
AND2x2_ASAP7_75t_L g311 ( .A(n_266), .B(n_290), .Y(n_311) );
AND2x2_ASAP7_75t_L g349 ( .A(n_266), .B(n_290), .Y(n_349) );
AND2x2_ASAP7_75t_SL g646 ( .A(n_266), .B(n_290), .Y(n_646) );
AND2x4_ASAP7_75t_L g305 ( .A(n_267), .B(n_278), .Y(n_305) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_SL g342 ( .A(n_269), .Y(n_342) );
INVx2_ASAP7_75t_L g371 ( .A(n_269), .Y(n_371) );
INVx2_ASAP7_75t_L g463 ( .A(n_269), .Y(n_463) );
INVx2_ASAP7_75t_L g504 ( .A(n_269), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_269), .B(n_542), .Y(n_541) );
INVx6_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx6f_ASAP7_75t_SL g557 ( .A(n_275), .Y(n_557) );
BUFx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
BUFx3_ASAP7_75t_L g339 ( .A(n_276), .Y(n_339) );
INVx2_ASAP7_75t_L g507 ( .A(n_276), .Y(n_507) );
AND2x2_ASAP7_75t_L g289 ( .A(n_277), .B(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g405 ( .A(n_277), .B(n_290), .Y(n_405) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_279), .Y(n_558) );
INVx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g609 ( .A(n_280), .Y(n_609) );
INVx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx12f_ASAP7_75t_L g375 ( .A(n_281), .Y(n_375) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x4_ASAP7_75t_L g304 ( .A(n_282), .B(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g313 ( .A(n_282), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g350 ( .A(n_282), .B(n_314), .Y(n_350) );
AND2x2_ASAP7_75t_SL g400 ( .A(n_282), .B(n_283), .Y(n_400) );
AND2x4_ASAP7_75t_L g415 ( .A(n_282), .B(n_305), .Y(n_415) );
AND2x2_ASAP7_75t_SL g490 ( .A(n_282), .B(n_283), .Y(n_490) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
INVx4_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g554 ( .A(n_288), .Y(n_554) );
INVx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_289), .Y(n_344) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_289), .Y(n_460) );
AND2x4_ASAP7_75t_L g330 ( .A(n_290), .B(n_305), .Y(n_330) );
AND2x6_ASAP7_75t_L g422 ( .A(n_290), .B(n_305), .Y(n_422) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_291), .Y(n_297) );
INVx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g502 ( .A(n_294), .Y(n_502) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g346 ( .A(n_295), .Y(n_346) );
BUFx3_ASAP7_75t_L g368 ( .A(n_295), .Y(n_368) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND4xp25_ASAP7_75t_L g298 ( .A(n_299), .B(n_306), .C(n_315), .D(n_324), .Y(n_298) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g535 ( .A(n_301), .Y(n_535) );
INVx1_ASAP7_75t_SL g569 ( .A(n_301), .Y(n_569) );
INVx6_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g352 ( .A(n_302), .Y(n_352) );
BUFx3_ASAP7_75t_L g392 ( .A(n_302), .Y(n_392) );
BUFx2_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
BUFx3_ASAP7_75t_L g353 ( .A(n_304), .Y(n_353) );
BUFx3_ASAP7_75t_L g444 ( .A(n_304), .Y(n_444) );
BUFx2_ASAP7_75t_SL g517 ( .A(n_304), .Y(n_517) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_309), .Y(n_514) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_309), .Y(n_530) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g388 ( .A(n_310), .Y(n_388) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx3_ASAP7_75t_L g440 ( .A(n_311), .Y(n_440) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_311), .Y(n_470) );
BUFx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx5_ASAP7_75t_SL g390 ( .A(n_313), .Y(n_390) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_318), .Y(n_516) );
INVx4_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx3_ASAP7_75t_L g359 ( .A(n_319), .Y(n_359) );
INVx3_ASAP7_75t_SL g380 ( .A(n_319), .Y(n_380) );
INVx2_ASAP7_75t_L g468 ( .A(n_319), .Y(n_468) );
INVx8_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g567 ( .A(n_322), .Y(n_567) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g357 ( .A(n_323), .Y(n_357) );
INVx2_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
INVx3_ASAP7_75t_L g355 ( .A(n_326), .Y(n_355) );
INVx2_ASAP7_75t_SL g511 ( .A(n_326), .Y(n_511) );
INVx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g385 ( .A(n_327), .Y(n_385) );
BUFx2_ASAP7_75t_L g533 ( .A(n_327), .Y(n_533) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g360 ( .A(n_329), .Y(n_360) );
INVx2_ASAP7_75t_SL g381 ( .A(n_329), .Y(n_381) );
INVx2_ASAP7_75t_L g512 ( .A(n_329), .Y(n_512) );
INVx8_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g361 ( .A(n_331), .Y(n_361) );
BUFx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_347), .Y(n_334) );
NAND4xp25_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .C(n_340), .D(n_343), .Y(n_335) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_339), .Y(n_373) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_346), .A2(n_631), .B1(n_632), .B2(n_633), .Y(n_630) );
NAND4xp25_ASAP7_75t_L g347 ( .A(n_348), .B(n_351), .C(n_354), .D(n_358), .Y(n_347) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g537 ( .A(n_357), .Y(n_537) );
INVx1_ASAP7_75t_L g450 ( .A(n_362), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_393), .B1(n_448), .B2(n_449), .Y(n_362) );
INVx1_ASAP7_75t_SL g448 ( .A(n_363), .Y(n_448) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_378), .Y(n_364) );
NAND4xp25_ASAP7_75t_L g365 ( .A(n_366), .B(n_369), .C(n_372), .D(n_376), .Y(n_365) );
BUFx6f_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g547 ( .A(n_375), .Y(n_547) );
NAND4xp25_ASAP7_75t_L g378 ( .A(n_379), .B(n_382), .C(n_386), .D(n_391), .Y(n_378) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g449 ( .A(n_393), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_424), .B1(n_425), .B2(n_447), .Y(n_393) );
INVx3_ASAP7_75t_SL g447 ( .A(n_394), .Y(n_447) );
XOR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_423), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_410), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_403), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_398), .B(n_401), .Y(n_397) );
INVx2_ASAP7_75t_SL g430 ( .A(n_402), .Y(n_430) );
BUFx2_ASAP7_75t_L g629 ( .A(n_402), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_407), .Y(n_403) );
INVxp67_ASAP7_75t_L g636 ( .A(n_408), .Y(n_636) );
INVxp67_ASAP7_75t_L g638 ( .A(n_409), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_416), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_420), .Y(n_416) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
XOR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_446), .Y(n_426) );
NAND2x1_ASAP7_75t_L g427 ( .A(n_428), .B(n_437), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_433), .Y(n_428) );
OAI21xp5_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_431), .B(n_432), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .Y(n_433) );
NOR2x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_442), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_441), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_445), .Y(n_442) );
INVx1_ASAP7_75t_L g587 ( .A(n_451), .Y(n_587) );
XOR2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_519), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_454), .B1(n_475), .B2(n_476), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g474 ( .A(n_457), .Y(n_474) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_466), .Y(n_457) );
NAND4xp25_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .C(n_464), .D(n_465), .Y(n_458) );
BUFx6f_ASAP7_75t_SL g540 ( .A(n_460), .Y(n_540) );
INVx1_ASAP7_75t_L g632 ( .A(n_460), .Y(n_632) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .C(n_471), .D(n_472), .Y(n_466) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
XNOR2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_497), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g496 ( .A(n_479), .Y(n_496) );
NOR2xp67_ASAP7_75t_L g479 ( .A(n_480), .B(n_486), .Y(n_479) );
NAND4xp25_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .C(n_483), .D(n_485), .Y(n_480) );
NAND4xp25_ASAP7_75t_SL g486 ( .A(n_487), .B(n_489), .C(n_491), .D(n_494), .Y(n_486) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NOR2xp67_ASAP7_75t_L g499 ( .A(n_500), .B(n_509), .Y(n_499) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .C(n_505), .D(n_508), .Y(n_500) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND4xp25_ASAP7_75t_L g509 ( .A(n_510), .B(n_513), .C(n_515), .D(n_518), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B1(n_571), .B2(n_586), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_549), .B2(n_570), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NOR2xp67_ASAP7_75t_L g527 ( .A(n_528), .B(n_538), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
NOR3xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .C(n_536), .Y(n_531) );
NAND4xp25_ASAP7_75t_L g538 ( .A(n_539), .B(n_543), .C(n_544), .D(n_545), .Y(n_538) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g570 ( .A(n_549), .Y(n_570) );
NOR2x1_ASAP7_75t_L g550 ( .A(n_551), .B(n_562), .Y(n_550) );
NAND4xp25_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .C(n_556), .D(n_559), .Y(n_551) );
BUFx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND4xp25_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .C(n_565), .D(n_568), .Y(n_562) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g586 ( .A(n_571), .Y(n_586) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_581), .Y(n_575) );
NAND4xp25_ASAP7_75t_SL g576 ( .A(n_577), .B(n_578), .C(n_579), .D(n_580), .Y(n_576) );
NAND4xp25_ASAP7_75t_SL g581 ( .A(n_582), .B(n_583), .C(n_584), .D(n_585), .Y(n_581) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_591), .B(n_594), .Y(n_650) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
OAI222xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_616), .B1(n_618), .B2(n_623), .C1(n_648), .C2(n_651), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g615 ( .A(n_600), .Y(n_615) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_607), .C(n_611), .Y(n_601) );
NAND4xp25_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .C(n_605), .D(n_606), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g647 ( .A(n_624), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_639), .Y(n_624) );
NOR3xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_630), .C(n_634), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_627), .B(n_628), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B1(n_637), .B2(n_638), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_643), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
CKINVDCx6p67_ASAP7_75t_R g649 ( .A(n_650), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_652), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_653), .Y(n_652) );
endmodule