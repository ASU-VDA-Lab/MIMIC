module real_jpeg_15270_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_SL g29 ( 
.A(n_0),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_486),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_1),
.B(n_487),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_2),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_2),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_2),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_2),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_2),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_2),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_2),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_2),
.B(n_36),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_3),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_3),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_3),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_4),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_4),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_5),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_5),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_5),
.B(n_83),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_5),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_5),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_5),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_5),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_5),
.B(n_240),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_6),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_6),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_6),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_6),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_6),
.B(n_42),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_6),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_7),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_7),
.B(n_47),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_7),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_7),
.B(n_258),
.Y(n_257)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_7),
.B(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_SL g401 ( 
.A(n_7),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_7),
.B(n_407),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_8),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_8),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_8),
.B(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_8),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_8),
.B(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_8),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_8),
.B(n_455),
.Y(n_454)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_9),
.Y(n_242)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_9),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_10),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_10),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g243 ( 
.A(n_10),
.B(n_244),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g294 ( 
.A(n_10),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g357 ( 
.A(n_10),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_10),
.B(n_53),
.Y(n_394)
);

AND2x2_ASAP7_75t_SL g396 ( 
.A(n_10),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_10),
.B(n_434),
.Y(n_433)
);

INVxp33_ASAP7_75t_L g487 ( 
.A(n_11),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_12),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_12),
.Y(n_104)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_12),
.Y(n_123)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_12),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g359 ( 
.A(n_12),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_12),
.Y(n_387)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_13),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_13),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_14),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_15),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_15),
.B(n_30),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g321 ( 
.A(n_15),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_15),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_15),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_15),
.B(n_430),
.Y(n_429)
);

AND2x2_ASAP7_75t_SL g441 ( 
.A(n_15),
.B(n_442),
.Y(n_441)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_16),
.Y(n_409)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g139 ( 
.A(n_17),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_17),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_179),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_R g20 ( 
.A(n_21),
.B(n_178),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_154),
.Y(n_22)
);

NOR2x1_ASAP7_75t_R g178 ( 
.A(n_23),
.B(n_154),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_94),
.C(n_129),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_24),
.B(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_66),
.C(n_80),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_25),
.B(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.C(n_51),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_26),
.B(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_27),
.B(n_35),
.C(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_28),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_28),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_28),
.B(n_91),
.Y(n_175)
);

NAND2x1_ASAP7_75t_L g220 ( 
.A(n_28),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_29),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_31),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_33),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_33),
.A2(n_38),
.B1(n_98),
.B2(n_105),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_33),
.B(n_213),
.Y(n_414)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_34),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_34),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_35),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_41),
.B(n_45),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_41),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_35),
.A2(n_37),
.B1(n_41),
.B2(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_35),
.B(n_406),
.Y(n_405)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_36),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_37),
.B(n_406),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_38),
.B(n_98),
.C(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_39),
.B(n_51),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_50),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_41),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_41),
.B(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_41),
.A2(n_195),
.B1(n_291),
.B2(n_292),
.Y(n_350)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_44),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_45),
.B(n_194),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_50),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_50),
.A2(n_320),
.B1(n_472),
.B2(n_473),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_52),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_52),
.B(n_102),
.C(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_64),
.B2(n_65),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_60),
.B(n_65),
.C(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_67),
.B(n_80),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_74),
.B1(n_78),
.B2(n_79),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_70),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_70),
.B(n_79),
.C(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_73),
.Y(n_215)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_73),
.Y(n_267)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_74),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_74),
.A2(n_79),
.B1(n_163),
.B2(n_169),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_74),
.A2(n_79),
.B1(n_92),
.B2(n_93),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_76),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_77),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g356 ( 
.A(n_77),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_81),
.C(n_92),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_81),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.C(n_89),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_82),
.A2(n_89),
.B1(n_90),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_82),
.Y(n_204)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2x1_ASAP7_75t_L g202 ( 
.A(n_86),
.B(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_89),
.B(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_89),
.B(n_138),
.C(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_94),
.A2(n_129),
.B1(n_130),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_94),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_106),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_95),
.B(n_107),
.C(n_114),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_96),
.B(n_98),
.C(n_102),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_98),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_98),
.B(n_294),
.C(n_297),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_98),
.A2(n_105),
.B1(n_294),
.B2(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g443 ( 
.A(n_100),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_101),
.A2(n_102),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_101),
.B(n_150),
.Y(n_317)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_104),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_114),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.C(n_124),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_118),
.Y(n_296)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_120),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_120),
.B(n_175),
.C(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_120),
.A2(n_153),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2x1_ASAP7_75t_SL g151 ( 
.A(n_125),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_146),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_135),
.C(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_143),
.B(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_151),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_151),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_170),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_175),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_175),
.A2(n_176),
.B1(n_197),
.B2(n_198),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_224),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_185),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_R g185 ( 
.A(n_186),
.B(n_188),
.C(n_191),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_186),
.B(n_189),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_191),
.B(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_205),
.C(n_209),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_192),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.C(n_202),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_193),
.B(n_196),
.Y(n_309)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_201),
.Y(n_328)
);

XOR2x1_ASAP7_75t_L g308 ( 
.A(n_202),
.B(n_309),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_275)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.C(n_220),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_211),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.C(n_214),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_213),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_216),
.A2(n_220),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_216),
.Y(n_271)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_220),
.Y(n_272)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_223),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_373),
.Y(n_226)
);

A2O1A1O1Ixp25_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_310),
.B(n_363),
.C(n_364),
.D(n_372),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_229),
.B(n_365),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_280),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_230),
.B(n_280),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_273),
.Y(n_230)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_231),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_256),
.C(n_268),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_233),
.B(n_283),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.C(n_246),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_234),
.B(n_330),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_236),
.A2(n_237),
.B1(n_246),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_237),
.A2(n_238),
.B(n_243),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_246),
.Y(n_331)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.C(n_251),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_248),
.Y(n_288)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_251),
.B(n_288),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_252),
.B(n_416),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_256),
.A2(n_268),
.B1(n_269),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_261),
.C(n_265),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_261),
.Y(n_303)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_264),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_266),
.B(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_273)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_276),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_276),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_278),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_285),
.C(n_307),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_281),
.A2(n_282),
.B1(n_308),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_302),
.C(n_304),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.C(n_293),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_287),
.B(n_344),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_289),
.A2(n_290),
.B1(n_293),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_294),
.Y(n_349)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_297),
.B(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_304),
.Y(n_314)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_335),
.B(n_362),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_332),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_312),
.B(n_332),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.C(n_329),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_329),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.C(n_319),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_318),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.C(n_326),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_321),
.A2(n_326),
.B1(n_327),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_321),
.Y(n_474)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_338),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_336),
.B(n_338),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_342),
.C(n_346),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_339),
.A2(n_340),
.B1(n_483),
.B2(n_484),
.Y(n_482)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_343),
.B(n_346),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_350),
.C(n_351),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_347),
.B(n_477),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_350),
.B(n_351),
.Y(n_477)
);

MAJx2_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_357),
.C(n_360),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_352),
.A2(n_353),
.B1(n_360),
.B2(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2x1_ASAP7_75t_L g422 ( 
.A(n_357),
.B(n_423),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_360),
.Y(n_424)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_362),
.Y(n_376)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_370),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_370),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.C(n_369),
.Y(n_366)
);

NAND4xp25_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.C(n_376),
.D(n_377),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_480),
.B(n_485),
.Y(n_377)
);

AOI21x1_ASAP7_75t_SL g378 ( 
.A1(n_379),
.A2(n_468),
.B(n_479),
.Y(n_378)
);

OAI21x1_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_425),
.B(n_467),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_410),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_381),
.B(n_410),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_395),
.C(n_404),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_382),
.B(n_464),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_388),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_394),
.C(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_385),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_394),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_389),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_395),
.A2(n_404),
.B1(n_405),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_401),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_396),
.B(n_401),
.Y(n_438)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_419),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_411),
.B(n_420),
.C(n_422),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_412),
.B(n_415),
.C(n_417),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_414),
.A2(n_415),
.B1(n_417),
.B2(n_418),
.Y(n_413)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_414),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_415),
.Y(n_418)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_416),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_422),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_461),
.B(n_466),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_427),
.A2(n_448),
.B(n_460),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_437),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_428),
.B(n_437),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_433),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_433),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_436),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_441),
.C(n_444),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_444),
.B2(n_445),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_453),
.B(n_459),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_452),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_462),
.B(n_463),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_478),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_478),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_476),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_475),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_475),
.C(n_476),
.Y(n_481)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_481),
.B(n_482),
.Y(n_485)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);


endmodule