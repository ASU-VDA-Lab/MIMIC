module real_jpeg_26206_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

INVx1_ASAP7_75t_L g79 ( 
.A(n_0),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_2),
.B(n_55),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_2),
.B(n_41),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_2),
.B(n_28),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_2),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_3),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_3),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_3),
.B(n_34),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_3),
.B(n_65),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_3),
.B(n_28),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_3),
.B(n_55),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_3),
.B(n_175),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_4),
.B(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_4),
.B(n_46),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_4),
.B(n_50),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_4),
.B(n_55),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_4),
.B(n_65),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_4),
.B(n_28),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_4),
.B(n_184),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

INVx8_ASAP7_75t_SL g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_9),
.B(n_50),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_9),
.B(n_41),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_9),
.B(n_65),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_9),
.B(n_28),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_9),
.B(n_46),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_10),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_10),
.B(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_10),
.B(n_50),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_10),
.B(n_82),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_11),
.B(n_28),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_11),
.B(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_12),
.B(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_12),
.B(n_65),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_12),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_12),
.B(n_50),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_12),
.B(n_55),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_12),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_12),
.B(n_28),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_15),
.B(n_65),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_16),
.B(n_65),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_16),
.B(n_50),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_16),
.B(n_55),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_16),
.B(n_28),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_16),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_16),
.B(n_41),
.Y(n_237)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_17),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_152),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_129),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_52),
.C(n_58),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_22),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.C(n_44),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_23),
.B(n_267),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_24),
.B(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_24),
.B(n_54),
.C(n_57),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.CI(n_33),
.CON(n_24),
.SN(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_36),
.A2(n_37),
.B(n_40),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_36),
.B(n_44),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_39),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.C(n_51),
.Y(n_44)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_45),
.B(n_49),
.CI(n_51),
.CON(n_133),
.SN(n_133)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_47),
.B(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_52),
.B(n_58),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_55),
.Y(n_214)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.C(n_69),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_59),
.B(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.C(n_64),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_60),
.B(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_61),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_63),
.B(n_64),
.Y(n_256)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_95),
.B2(n_128),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_86),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_79),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_84),
.B1(n_88),
.B2(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_83),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_88),
.C(n_89),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_90),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_91),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.CI(n_94),
.CON(n_91),
.SN(n_91)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_117),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_107),
.C(n_113),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_102),
.C(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_103),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_113),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.C(n_111),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_127),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_123),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_148),
.C(n_150),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_130),
.A2(n_131),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_144),
.C(n_146),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_132),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.C(n_140),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_133),
.B(n_249),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_133),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_134),
.A2(n_135),
.B1(n_140),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_140),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.C(n_143),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_141),
.B(n_142),
.CI(n_143),
.CON(n_230),
.SN(n_230)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_144),
.B(n_146),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_148),
.B(n_150),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_269),
.C(n_270),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_259),
.C(n_260),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_242),
.C(n_243),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_224),
.C(n_225),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_186),
.C(n_197),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_171),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_166),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_159),
.B(n_166),
.C(n_171),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_161),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_167),
.B(n_169),
.C(n_170),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_178),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_179),
.C(n_180),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_185),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_181),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_185),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_196),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_191),
.B1(n_196),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_220),
.C(n_221),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_206),
.C(n_211),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_204),
.C(n_205),
.Y(n_220)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.C(n_215),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_232),
.C(n_241),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_229),
.C(n_230),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_230),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_241),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_239),
.B2(n_240),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_235),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_238),
.C(n_240),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_239),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_251),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_247),
.C(n_251),
.Y(n_259)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_255),
.C(n_257),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_254),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_255),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_268),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_265),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);


endmodule