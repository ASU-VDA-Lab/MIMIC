module fake_netlist_6_2841_n_777 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_777);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_777;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_81),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_22),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_87),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

BUFx8_ASAP7_75t_SL g168 ( 
.A(n_24),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_60),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_9),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_13),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_31),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_89),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_29),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_85),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_116),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_76),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_66),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_30),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_112),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_20),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_90),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_58),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_8),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_21),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_26),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_11),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_2),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_40),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_53),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_102),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_17),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_69),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_16),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_15),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_13),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_71),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_151),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_55),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_65),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_68),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_143),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_105),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_154),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_173),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_0),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_202),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_167),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_161),
.B(n_0),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_169),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_168),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_1),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

INVxp33_ASAP7_75t_SL g238 ( 
.A(n_162),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_163),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_161),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_160),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_164),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_182),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_165),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_166),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_176),
.B(n_1),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_201),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_210),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_192),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_170),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_227),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_172),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_174),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_175),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_217),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_225),
.B(n_211),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_219),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_221),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_217),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_224),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_229),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_236),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_231),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_246),
.B(n_193),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_236),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_228),
.B(n_2),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_246),
.A2(n_216),
.B1(n_215),
.B2(n_214),
.Y(n_287)
);

AND2x6_ASAP7_75t_L g288 ( 
.A(n_251),
.B(n_193),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_225),
.B(n_218),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_233),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_252),
.A2(n_191),
.B1(n_208),
.B2(n_206),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_237),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_235),
.B(n_193),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_222),
.B(n_177),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_223),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_238),
.B(n_180),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_240),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_223),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_247),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

BUFx8_ASAP7_75t_L g306 ( 
.A(n_234),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_226),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_258),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_258),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_226),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

NAND3x1_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_252),
.C(n_228),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_259),
.C(n_198),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_260),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_283),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_277),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_238),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_303),
.B(n_213),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_232),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_276),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_298),
.A2(n_189),
.B1(n_184),
.B2(n_203),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_262),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_183),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_232),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_266),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_186),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_188),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_197),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_199),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_303),
.B(n_213),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_277),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_270),
.B(n_213),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_213),
.Y(n_343)
);

BUFx4_ASAP7_75t_L g344 ( 
.A(n_306),
.Y(n_344)
);

NAND2x1p5_ASAP7_75t_L g345 ( 
.A(n_303),
.B(n_19),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_305),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_267),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_3),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_263),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_268),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_300),
.B(n_3),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_282),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_296),
.B(n_23),
.Y(n_353)
);

AO22x2_ASAP7_75t_L g354 ( 
.A1(n_286),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_265),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_289),
.B(n_25),
.Y(n_356)
);

AND2x2_ASAP7_75t_SL g357 ( 
.A(n_284),
.B(n_4),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_269),
.B(n_27),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_289),
.B(n_28),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_265),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_275),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_278),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_306),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_269),
.B(n_32),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_271),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_272),
.Y(n_366)
);

AND2x2_ASAP7_75t_SL g367 ( 
.A(n_303),
.B(n_5),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_278),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_275),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_303),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_261),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_288),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_304),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_373)
);

OR2x6_ASAP7_75t_L g374 ( 
.A(n_304),
.B(n_12),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_316),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_315),
.B(n_274),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_318),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_326),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_338),
.Y(n_379)
);

OAI221xp5_ASAP7_75t_L g380 ( 
.A1(n_372),
.A2(n_279),
.B1(n_292),
.B2(n_281),
.C(n_299),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_363),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_325),
.Y(n_382)
);

AO22x2_ASAP7_75t_L g383 ( 
.A1(n_370),
.A2(n_286),
.B1(n_287),
.B2(n_297),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_331),
.Y(n_384)
);

AO22x2_ASAP7_75t_L g385 ( 
.A1(n_373),
.A2(n_297),
.B1(n_270),
.B2(n_305),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_313),
.B(n_304),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

NAND2x1p5_ASAP7_75t_L g388 ( 
.A(n_315),
.B(n_356),
.Y(n_388)
);

NAND2x1p5_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_304),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_367),
.A2(n_357),
.B1(n_359),
.B2(n_372),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_347),
.B(n_274),
.Y(n_391)
);

OR2x6_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_304),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_309),
.B(n_291),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_342),
.B(n_264),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_336),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_274),
.Y(n_397)
);

AND2x6_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_264),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_322),
.B(n_277),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_323),
.B(n_280),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_362),
.Y(n_401)
);

NAND2x1_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_288),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_321),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_310),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_343),
.B(n_280),
.Y(n_405)
);

AO22x2_ASAP7_75t_L g406 ( 
.A1(n_354),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_330),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_343),
.B(n_280),
.Y(n_408)
);

INVx6_ASAP7_75t_L g409 ( 
.A(n_346),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_314),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_366),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_357),
.B(n_306),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_334),
.B(n_280),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_368),
.Y(n_415)
);

NAND2x1p5_ASAP7_75t_L g416 ( 
.A(n_367),
.B(n_320),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_361),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_361),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_374),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_319),
.B(n_292),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_369),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_374),
.B(n_285),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_332),
.B(n_285),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_334),
.B(n_280),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

AO22x2_ASAP7_75t_L g427 ( 
.A1(n_354),
.A2(n_17),
.B1(n_18),
.B2(n_261),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_337),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_324),
.Y(n_429)
);

AO22x2_ASAP7_75t_L g430 ( 
.A1(n_354),
.A2(n_18),
.B1(n_261),
.B2(n_288),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_314),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_329),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_355),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_337),
.A2(n_288),
.B1(n_282),
.B2(n_35),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_329),
.Y(n_435)
);

OAI221xp5_ASAP7_75t_L g436 ( 
.A1(n_348),
.A2(n_282),
.B1(n_288),
.B2(n_36),
.C(n_37),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_360),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_358),
.B(n_33),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_348),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_320),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_360),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_353),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_351),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_327),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_390),
.B(n_404),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_394),
.B(n_327),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_444),
.B(n_333),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_SL g449 ( 
.A(n_429),
.B(n_364),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_439),
.B(n_333),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_376),
.B(n_351),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_415),
.B(n_339),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_SL g453 ( 
.A(n_381),
.B(n_339),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_386),
.B(n_345),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_395),
.B(n_311),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_413),
.B(n_345),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_376),
.B(n_311),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_403),
.B(n_352),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_389),
.B(n_423),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_398),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_SL g461 ( 
.A(n_407),
.B(n_344),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_423),
.B(n_341),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_SL g463 ( 
.A(n_378),
.B(n_438),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_377),
.B(n_341),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_424),
.B(n_352),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_398),
.B(n_317),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_375),
.B(n_317),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_382),
.B(n_340),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_398),
.B(n_328),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_391),
.B(n_397),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_398),
.B(n_328),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_335),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_SL g473 ( 
.A(n_438),
.B(n_312),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_384),
.B(n_340),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_393),
.B(n_335),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_411),
.B(n_288),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_391),
.B(n_34),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_397),
.B(n_38),
.Y(n_478)
);

NAND2xp33_ASAP7_75t_SL g479 ( 
.A(n_441),
.B(n_39),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_388),
.B(n_41),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_414),
.B(n_42),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_379),
.B(n_43),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_401),
.B(n_44),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_416),
.B(n_45),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_420),
.B(n_392),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_425),
.B(n_46),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_421),
.B(n_47),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_440),
.B(n_48),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_399),
.B(n_49),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_SL g490 ( 
.A(n_402),
.B(n_392),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_417),
.B(n_50),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_400),
.B(n_51),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_434),
.B(n_52),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_418),
.B(n_419),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_422),
.B(n_54),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_410),
.B(n_56),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_410),
.B(n_57),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_405),
.B(n_59),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_466),
.A2(n_402),
.B(n_408),
.Y(n_499)
);

NOR4xp25_ASAP7_75t_L g500 ( 
.A(n_447),
.B(n_436),
.C(n_380),
.D(n_406),
.Y(n_500)
);

A2O1A1Ixp33_ASAP7_75t_L g501 ( 
.A1(n_445),
.A2(n_431),
.B(n_432),
.C(n_435),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_458),
.B(n_383),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_450),
.B(n_387),
.Y(n_503)
);

AOI21x1_ASAP7_75t_L g504 ( 
.A1(n_454),
.A2(n_442),
.B(n_437),
.Y(n_504)
);

CKINVDCx11_ASAP7_75t_R g505 ( 
.A(n_485),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_448),
.B(n_385),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_469),
.A2(n_426),
.B(n_412),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_452),
.Y(n_508)
);

AO21x2_ASAP7_75t_L g509 ( 
.A1(n_481),
.A2(n_396),
.B(n_433),
.Y(n_509)
);

CKINVDCx14_ASAP7_75t_R g510 ( 
.A(n_461),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_455),
.A2(n_385),
.B(n_383),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_494),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_465),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_471),
.A2(n_61),
.B(n_62),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_446),
.B(n_451),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_451),
.B(n_430),
.Y(n_516)
);

AOI31xp67_ASAP7_75t_L g517 ( 
.A1(n_486),
.A2(n_430),
.A3(n_427),
.B(n_406),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_485),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_472),
.A2(n_427),
.B(n_64),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_470),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_470),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_460),
.A2(n_63),
.B(n_67),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_491),
.A2(n_476),
.B(n_475),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_459),
.B(n_409),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_493),
.A2(n_70),
.B(n_72),
.Y(n_525)
);

NAND3xp33_ASAP7_75t_SL g526 ( 
.A(n_449),
.B(n_409),
.C(n_75),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_484),
.A2(n_74),
.B(n_77),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_467),
.A2(n_78),
.B(n_79),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_490),
.A2(n_80),
.B(n_82),
.Y(n_529)
);

AO32x2_ASAP7_75t_L g530 ( 
.A1(n_456),
.A2(n_159),
.A3(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_530)
);

OAI22x1_ASAP7_75t_L g531 ( 
.A1(n_482),
.A2(n_83),
.B1(n_91),
.B2(n_92),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_473),
.B(n_93),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_457),
.A2(n_94),
.B(n_95),
.Y(n_533)
);

AO31x2_ASAP7_75t_L g534 ( 
.A1(n_498),
.A2(n_96),
.A3(n_97),
.B(n_98),
.Y(n_534)
);

NAND3x1_ASAP7_75t_L g535 ( 
.A(n_453),
.B(n_99),
.C(n_100),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_462),
.B(n_101),
.Y(n_536)
);

INVx8_ASAP7_75t_L g537 ( 
.A(n_463),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_483),
.Y(n_538)
);

AOI21x1_ASAP7_75t_L g539 ( 
.A1(n_468),
.A2(n_103),
.B(n_104),
.Y(n_539)
);

O2A1O1Ixp5_ASAP7_75t_L g540 ( 
.A1(n_487),
.A2(n_106),
.B(n_107),
.C(n_109),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_479),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_477),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_537),
.B(n_480),
.Y(n_543)
);

OAI21x1_ASAP7_75t_L g544 ( 
.A1(n_499),
.A2(n_489),
.B(n_492),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_506),
.B(n_464),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_515),
.B(n_478),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_508),
.B(n_474),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_511),
.B(n_488),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_513),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_518),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_507),
.A2(n_497),
.B(n_496),
.Y(n_551)
);

AO32x2_ASAP7_75t_L g552 ( 
.A1(n_541),
.A2(n_495),
.A3(n_115),
.B1(n_118),
.B2(n_120),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_502),
.A2(n_516),
.B1(n_519),
.B2(n_532),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_504),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_538),
.B(n_114),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_520),
.A2(n_121),
.B1(n_123),
.B2(n_126),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g557 ( 
.A1(n_523),
.A2(n_528),
.B(n_514),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_512),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_500),
.A2(n_127),
.B(n_129),
.Y(n_559)
);

NAND2x1p5_ASAP7_75t_L g560 ( 
.A(n_520),
.B(n_130),
.Y(n_560)
);

AO21x2_ASAP7_75t_L g561 ( 
.A1(n_509),
.A2(n_131),
.B(n_132),
.Y(n_561)
);

AO21x2_ASAP7_75t_L g562 ( 
.A1(n_501),
.A2(n_527),
.B(n_529),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_521),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_539),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_503),
.A2(n_133),
.B(n_134),
.Y(n_565)
);

O2A1O1Ixp33_ASAP7_75t_SL g566 ( 
.A1(n_542),
.A2(n_135),
.B(n_136),
.C(n_138),
.Y(n_566)
);

OA21x2_ASAP7_75t_L g567 ( 
.A1(n_540),
.A2(n_140),
.B(n_142),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_524),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_521),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_569)
);

AOI31xp67_ASAP7_75t_L g570 ( 
.A1(n_536),
.A2(n_150),
.A3(n_153),
.B(n_155),
.Y(n_570)
);

NAND2x1p5_ASAP7_75t_L g571 ( 
.A(n_521),
.B(n_156),
.Y(n_571)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_522),
.A2(n_157),
.B(n_525),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_534),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_517),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_541),
.A2(n_537),
.B1(n_535),
.B2(n_510),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_533),
.A2(n_526),
.B(n_534),
.Y(n_576)
);

OA21x2_ASAP7_75t_L g577 ( 
.A1(n_530),
.A2(n_534),
.B(n_531),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_505),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_530),
.B(n_511),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_530),
.B(n_428),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_513),
.Y(n_581)
);

NAND3xp33_ASAP7_75t_L g582 ( 
.A(n_508),
.B(n_447),
.C(n_394),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_550),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_549),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_568),
.B(n_582),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_558),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_580),
.B(n_579),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_581),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_574),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_545),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_563),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_554),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_573),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_554),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_543),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_547),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_578),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_563),
.Y(n_598)
);

OAI21xp33_ASAP7_75t_SL g599 ( 
.A1(n_559),
.A2(n_546),
.B(n_565),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_571),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_573),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_577),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_571),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_564),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_562),
.A2(n_546),
.B(n_572),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_560),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_553),
.B(n_548),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_548),
.B(n_555),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_575),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_577),
.Y(n_610)
);

OR2x6_ASAP7_75t_L g611 ( 
.A(n_543),
.B(n_557),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_579),
.B(n_552),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_560),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_543),
.B(n_572),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_552),
.B(n_577),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g616 ( 
.A1(n_557),
.A2(n_544),
.B(n_551),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_564),
.Y(n_617)
);

AOI21x1_ASAP7_75t_L g618 ( 
.A1(n_576),
.A2(n_544),
.B(n_551),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_564),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_561),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_561),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_561),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_578),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_543),
.A2(n_562),
.B1(n_556),
.B2(n_569),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_562),
.B(n_576),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_570),
.Y(n_626)
);

CKINVDCx11_ASAP7_75t_R g627 ( 
.A(n_566),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_566),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_567),
.Y(n_629)
);

OR2x2_ASAP7_75t_SL g630 ( 
.A(n_567),
.B(n_582),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_558),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_583),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_608),
.B(n_609),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_590),
.B(n_596),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_595),
.B(n_600),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_R g636 ( 
.A(n_597),
.B(n_585),
.Y(n_636)
);

OR2x6_ASAP7_75t_L g637 ( 
.A(n_595),
.B(n_603),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_584),
.Y(n_638)
);

OR2x6_ASAP7_75t_L g639 ( 
.A(n_595),
.B(n_606),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_607),
.B(n_586),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_613),
.B(n_599),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_631),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_614),
.B(n_611),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_614),
.B(n_624),
.Y(n_644)
);

BUFx10_ASAP7_75t_L g645 ( 
.A(n_597),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_623),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_588),
.B(n_614),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_R g648 ( 
.A(n_611),
.B(n_587),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_611),
.B(n_591),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_628),
.B(n_598),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_592),
.B(n_594),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_592),
.B(n_594),
.Y(n_652)
);

XOR2xp5_ASAP7_75t_L g653 ( 
.A(n_605),
.B(n_619),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_R g654 ( 
.A(n_611),
.B(n_602),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_604),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_R g656 ( 
.A(n_627),
.B(n_589),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_604),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_612),
.B(n_619),
.Y(n_658)
);

CKINVDCx12_ASAP7_75t_R g659 ( 
.A(n_617),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_617),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_593),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_612),
.B(n_627),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_630),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_R g664 ( 
.A(n_618),
.B(n_593),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_SL g665 ( 
.A(n_625),
.B(n_621),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_601),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_601),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_630),
.Y(n_668)
);

BUFx10_ASAP7_75t_L g669 ( 
.A(n_626),
.Y(n_669)
);

INVxp67_ASAP7_75t_SL g670 ( 
.A(n_666),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_658),
.B(n_615),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_647),
.B(n_615),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_643),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_667),
.Y(n_674)
);

AND2x2_ASAP7_75t_SL g675 ( 
.A(n_662),
.B(n_621),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_663),
.B(n_610),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_668),
.B(n_610),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_638),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_643),
.B(n_620),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_646),
.B(n_618),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_661),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_640),
.B(n_622),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_651),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_649),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_653),
.B(n_629),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_649),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_642),
.B(n_629),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_632),
.B(n_616),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_655),
.B(n_616),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_633),
.B(n_634),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_644),
.A2(n_641),
.B1(n_656),
.B2(n_635),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_652),
.Y(n_692)
);

AND2x2_ASAP7_75t_SL g693 ( 
.A(n_654),
.B(n_648),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_674),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_673),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_676),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_690),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_688),
.B(n_665),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_674),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_678),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_672),
.B(n_664),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_672),
.B(n_669),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_676),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_678),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_671),
.B(n_669),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_671),
.B(n_650),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_SL g707 ( 
.A1(n_691),
.A2(n_636),
.B(n_635),
.Y(n_707)
);

NAND3xp33_ASAP7_75t_SL g708 ( 
.A(n_680),
.B(n_657),
.C(n_660),
.Y(n_708)
);

AND2x2_ASAP7_75t_SL g709 ( 
.A(n_693),
.B(n_659),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_681),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_697),
.B(n_690),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_700),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_702),
.B(n_695),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_694),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_704),
.Y(n_715)
);

NOR2x1p5_ASAP7_75t_L g716 ( 
.A(n_708),
.B(n_673),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_694),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_698),
.B(n_685),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_699),
.Y(n_719)
);

NAND2x1p5_ASAP7_75t_L g720 ( 
.A(n_709),
.B(n_693),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_696),
.B(n_688),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_714),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_713),
.B(n_701),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_720),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_718),
.B(n_703),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_718),
.B(n_710),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_L g727 ( 
.A1(n_720),
.A2(n_707),
.B1(n_684),
.B2(n_673),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_711),
.B(n_685),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_724),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_722),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_726),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_725),
.Y(n_732)
);

AOI33xp33_ASAP7_75t_L g733 ( 
.A1(n_732),
.A2(n_727),
.A3(n_715),
.B1(n_712),
.B2(n_706),
.B3(n_681),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_729),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_731),
.A2(n_724),
.B(n_709),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_729),
.A2(n_716),
.B1(n_693),
.B2(n_728),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_734),
.B(n_645),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_733),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_735),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_738),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_737),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_739),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_738),
.Y(n_743)
);

NOR3x1_ASAP7_75t_SL g744 ( 
.A(n_740),
.B(n_645),
.C(n_736),
.Y(n_744)
);

NAND3x1_ASAP7_75t_SL g745 ( 
.A(n_742),
.B(n_723),
.C(n_701),
.Y(n_745)
);

NOR4xp25_ASAP7_75t_L g746 ( 
.A(n_743),
.B(n_730),
.C(n_698),
.D(n_721),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_SL g747 ( 
.A(n_741),
.B(n_730),
.C(n_695),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_740),
.A2(n_675),
.B1(n_713),
.B2(n_673),
.Y(n_748)
);

OAI211xp5_ASAP7_75t_SL g749 ( 
.A1(n_740),
.A2(n_717),
.B(n_686),
.C(n_682),
.Y(n_749)
);

OAI221xp5_ASAP7_75t_SL g750 ( 
.A1(n_746),
.A2(n_744),
.B1(n_748),
.B2(n_745),
.C(n_747),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_749),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_746),
.B(n_719),
.Y(n_752)
);

AOI221xp5_ASAP7_75t_L g753 ( 
.A1(n_746),
.A2(n_692),
.B1(n_706),
.B2(n_705),
.C(n_683),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_745),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_751),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_754),
.Y(n_756)
);

OAI211xp5_ASAP7_75t_L g757 ( 
.A1(n_750),
.A2(n_684),
.B(n_686),
.C(n_705),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_752),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_757),
.B(n_756),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_758),
.B(n_753),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_755),
.B(n_702),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_761),
.Y(n_762)
);

XOR2x1_ASAP7_75t_L g763 ( 
.A(n_759),
.B(n_677),
.Y(n_763)
);

NAND4xp75_ASAP7_75t_L g764 ( 
.A(n_760),
.B(n_675),
.C(n_677),
.D(n_687),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_762),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_763),
.B(n_684),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_764),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_763),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_767),
.A2(n_637),
.B1(n_686),
.B2(n_639),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_768),
.A2(n_682),
.B(n_675),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_769),
.A2(n_765),
.B1(n_766),
.B2(n_686),
.Y(n_771)
);

AOI31xp33_ASAP7_75t_L g772 ( 
.A1(n_770),
.A2(n_670),
.A3(n_683),
.B(n_692),
.Y(n_772)
);

NAND4xp25_ASAP7_75t_L g773 ( 
.A(n_771),
.B(n_679),
.C(n_689),
.D(n_687),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_773),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_774),
.Y(n_775)
);

OAI221xp5_ASAP7_75t_R g776 ( 
.A1(n_775),
.A2(n_772),
.B1(n_637),
.B2(n_639),
.C(n_670),
.Y(n_776)
);

AOI211xp5_ASAP7_75t_L g777 ( 
.A1(n_776),
.A2(n_699),
.B(n_679),
.C(n_689),
.Y(n_777)
);


endmodule