module fake_ariane_2039_n_857 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_857);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_857;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_779;
wire n_731;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_852;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_130),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_31),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_156),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_113),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_41),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_39),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_76),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_81),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_147),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_33),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_50),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_109),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_32),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_35),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_44),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_30),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_133),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_122),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_7),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_4),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_64),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_123),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_124),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_79),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_144),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_97),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_150),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_95),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_98),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_14),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_145),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_80),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_157),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_84),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_126),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_92),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_111),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_117),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_18),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_49),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_6),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_27),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_110),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_17),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_151),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_138),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_114),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_12),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_104),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_20),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_57),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_38),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_24),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_6),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_55),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_119),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_1),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_70),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_85),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

BUFx8_ASAP7_75t_SL g239 ( 
.A(n_179),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_0),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_214),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_218),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

BUFx8_ASAP7_75t_SL g247 ( 
.A(n_231),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_166),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

CKINVDCx6p67_ASAP7_75t_R g250 ( 
.A(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_2),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_171),
.B(n_3),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_173),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_181),
.Y(n_257)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_222),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_189),
.B(n_5),
.Y(n_261)
);

AND2x4_ASAP7_75t_L g262 ( 
.A(n_204),
.B(n_217),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_204),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_184),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_208),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_193),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_208),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_7),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_194),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_208),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_196),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_198),
.B(n_8),
.Y(n_272)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_208),
.Y(n_273)
);

BUFx8_ASAP7_75t_SL g274 ( 
.A(n_227),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_167),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_200),
.Y(n_276)
);

BUFx8_ASAP7_75t_L g277 ( 
.A(n_227),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_195),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_201),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_168),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_202),
.B(n_8),
.Y(n_281)
);

OAI21x1_ASAP7_75t_L g282 ( 
.A1(n_212),
.A2(n_88),
.B(n_164),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_169),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_177),
.A2(n_178),
.B1(n_221),
.B2(n_183),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_R g286 ( 
.A(n_244),
.B(n_246),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_239),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_239),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_223),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_245),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_264),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_264),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_248),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_238),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_247),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_275),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_250),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_243),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_245),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_182),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_274),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_285),
.B(n_228),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_R g307 ( 
.A(n_259),
.B(n_235),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_251),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_249),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_274),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_269),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g312 ( 
.A(n_252),
.B(n_229),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_R g313 ( 
.A(n_266),
.B(n_233),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_R g314 ( 
.A(n_280),
.B(n_170),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_253),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_284),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_253),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_280),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_172),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_280),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_277),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_277),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_279),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_278),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_242),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_278),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_278),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_R g329 ( 
.A(n_263),
.B(n_174),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_278),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_279),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_283),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_253),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_SL g334 ( 
.A(n_268),
.B(n_232),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_283),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_256),
.B(n_175),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_283),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_311),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

NAND2x1_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_262),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_309),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_302),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_291),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_281),
.Y(n_344)
);

BUFx6f_ASAP7_75t_SL g345 ( 
.A(n_321),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_293),
.B(n_263),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_291),
.B(n_262),
.Y(n_348)
);

CKINVDCx11_ASAP7_75t_R g349 ( 
.A(n_290),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_294),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_300),
.B(n_254),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_324),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_292),
.B(n_257),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_292),
.B(n_276),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_325),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_327),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_328),
.Y(n_357)
);

OR2x6_ASAP7_75t_L g358 ( 
.A(n_296),
.B(n_237),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_315),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_317),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_330),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_300),
.B(n_254),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_308),
.B(n_241),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_331),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_312),
.B(n_283),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_312),
.B(n_332),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_312),
.B(n_261),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_307),
.B(n_261),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_335),
.Y(n_370)
);

NOR3xp33_ASAP7_75t_L g371 ( 
.A(n_301),
.B(n_237),
.C(n_260),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

NOR3xp33_ASAP7_75t_L g373 ( 
.A(n_308),
.B(n_260),
.C(n_272),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_289),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_312),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_241),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_303),
.B(n_272),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_336),
.Y(n_378)
);

NOR3xp33_ASAP7_75t_L g379 ( 
.A(n_295),
.B(n_282),
.C(n_180),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_336),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_240),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_297),
.B(n_298),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_326),
.B(n_299),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_320),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_304),
.B(n_176),
.Y(n_385)
);

NAND3xp33_ASAP7_75t_L g386 ( 
.A(n_334),
.B(n_187),
.C(n_186),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_306),
.B(n_240),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_319),
.B(n_240),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_313),
.B(n_188),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_329),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_322),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_310),
.B(n_240),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_314),
.B(n_192),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_287),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_286),
.B(n_258),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_288),
.Y(n_396)
);

AND2x6_ASAP7_75t_SL g397 ( 
.A(n_290),
.B(n_9),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_291),
.B(n_273),
.Y(n_398)
);

A2O1A1Ixp33_ASAP7_75t_L g399 ( 
.A1(n_334),
.A2(n_219),
.B(n_199),
.C(n_203),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_316),
.B(n_197),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_309),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_309),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_309),
.Y(n_403)
);

BUFx6f_ASAP7_75t_SL g404 ( 
.A(n_321),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_334),
.A2(n_224),
.B1(n_207),
.B2(n_209),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_312),
.B(n_205),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_312),
.B(n_211),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_291),
.B(n_258),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_291),
.B(n_258),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_346),
.B(n_9),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_213),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_380),
.B(n_220),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_364),
.B(n_10),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_347),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_377),
.B(n_226),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_373),
.A2(n_270),
.B1(n_267),
.B2(n_265),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_341),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_349),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_368),
.A2(n_270),
.B1(n_267),
.B2(n_265),
.Y(n_420)
);

XOR2x2_ASAP7_75t_L g421 ( 
.A(n_371),
.B(n_10),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_350),
.A2(n_270),
.B1(n_267),
.B2(n_265),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_344),
.B(n_253),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_358),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_374),
.B(n_11),
.Y(n_425)
);

NOR3xp33_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_13),
.C(n_14),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_395),
.B(n_265),
.Y(n_427)
);

NAND3xp33_ASAP7_75t_L g428 ( 
.A(n_368),
.B(n_270),
.C(n_267),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_338),
.B(n_15),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_339),
.B(n_383),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_403),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_375),
.B(n_258),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_343),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_359),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_392),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_343),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_361),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_395),
.B(n_348),
.Y(n_440)
);

AO22x1_ASAP7_75t_L g441 ( 
.A1(n_382),
.A2(n_273),
.B1(n_15),
.B2(n_19),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_352),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_401),
.Y(n_443)
);

NOR2x1_ASAP7_75t_L g444 ( 
.A(n_390),
.B(n_273),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_353),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_354),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_408),
.A2(n_409),
.B(n_398),
.Y(n_447)
);

BUFx4f_ASAP7_75t_L g448 ( 
.A(n_394),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_360),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_375),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_406),
.A2(n_273),
.B1(n_21),
.B2(n_22),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_375),
.B(n_16),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_365),
.B(n_23),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_370),
.B(n_25),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_360),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_348),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_408),
.Y(n_458)
);

NOR3xp33_ASAP7_75t_SL g459 ( 
.A(n_400),
.B(n_26),
.C(n_28),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_379),
.A2(n_29),
.B1(n_34),
.B2(n_36),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_340),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_372),
.B(n_165),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_376),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_406),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_407),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_345),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_366),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_366),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_369),
.B(n_47),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_355),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_409),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_367),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_356),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_357),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_362),
.B(n_163),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_351),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_384),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_367),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_363),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_407),
.B(n_48),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_387),
.B(n_51),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_358),
.B(n_345),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_405),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_421),
.A2(n_358),
.B1(n_386),
.B2(n_389),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_R g485 ( 
.A(n_466),
.B(n_385),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_R g486 ( 
.A(n_419),
.B(n_385),
.Y(n_486)
);

O2A1O1Ixp33_ASAP7_75t_L g487 ( 
.A1(n_424),
.A2(n_399),
.B(n_393),
.C(n_381),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_451),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_447),
.A2(n_440),
.B(n_458),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_432),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_451),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_416),
.A2(n_381),
.B1(n_388),
.B2(n_404),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_448),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_442),
.Y(n_494)
);

OAI21xp33_ASAP7_75t_L g495 ( 
.A1(n_425),
.A2(n_404),
.B(n_397),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_468),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_412),
.Y(n_497)
);

A2O1A1Ixp33_ASAP7_75t_SL g498 ( 
.A1(n_411),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_415),
.Y(n_499)
);

O2A1O1Ixp33_ASAP7_75t_L g500 ( 
.A1(n_424),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_468),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_436),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_448),
.B(n_60),
.Y(n_504)
);

OAI22x1_ASAP7_75t_L g505 ( 
.A1(n_414),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_463),
.B(n_65),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_414),
.A2(n_455),
.B1(n_473),
.B2(n_470),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_482),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_416),
.B(n_445),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_437),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_471),
.Y(n_511)
);

OR2x6_ASAP7_75t_L g512 ( 
.A(n_482),
.B(n_66),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_443),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_423),
.A2(n_67),
.B(n_68),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_439),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_446),
.B(n_69),
.Y(n_516)
);

BUFx4f_ASAP7_75t_L g517 ( 
.A(n_482),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_410),
.B(n_71),
.Y(n_518)
);

BUFx12f_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_455),
.Y(n_520)
);

NAND2x1p5_ASAP7_75t_L g521 ( 
.A(n_461),
.B(n_72),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_R g522 ( 
.A(n_476),
.B(n_73),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_435),
.Y(n_523)
);

O2A1O1Ixp33_ASAP7_75t_L g524 ( 
.A1(n_413),
.A2(n_74),
.B(n_75),
.C(n_77),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_449),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_474),
.B(n_78),
.Y(n_526)
);

A2O1A1Ixp33_ASAP7_75t_L g527 ( 
.A1(n_469),
.A2(n_82),
.B(n_83),
.C(n_86),
.Y(n_527)
);

A2O1A1Ixp33_ASAP7_75t_L g528 ( 
.A1(n_462),
.A2(n_87),
.B(n_89),
.C(n_90),
.Y(n_528)
);

BUFx8_ASAP7_75t_SL g529 ( 
.A(n_477),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_479),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_472),
.A2(n_96),
.B(n_99),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_413),
.B(n_160),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_438),
.A2(n_100),
.B(n_101),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_429),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_450),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_418),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_478),
.B(n_467),
.Y(n_537)
);

O2A1O1Ixp33_ASAP7_75t_L g538 ( 
.A1(n_426),
.A2(n_102),
.B(n_103),
.C(n_105),
.Y(n_538)
);

AO21x1_ASAP7_75t_L g539 ( 
.A1(n_480),
.A2(n_159),
.B(n_107),
.Y(n_539)
);

OAI22x1_ASAP7_75t_L g540 ( 
.A1(n_417),
.A2(n_106),
.B1(n_108),
.B2(n_112),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_431),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_494),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_490),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_511),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_501),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_497),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_517),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_489),
.A2(n_481),
.B(n_427),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_499),
.Y(n_549)
);

AO21x2_ASAP7_75t_L g550 ( 
.A1(n_516),
.A2(n_481),
.B(n_428),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_520),
.B(n_441),
.Y(n_551)
);

AO21x2_ASAP7_75t_L g552 ( 
.A1(n_532),
.A2(n_428),
.B(n_475),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_513),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_531),
.A2(n_456),
.B(n_453),
.Y(n_554)
);

NAND2x1p5_ASAP7_75t_L g555 ( 
.A(n_491),
.B(n_478),
.Y(n_555)
);

BUFx4f_ASAP7_75t_SL g556 ( 
.A(n_519),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_493),
.B(n_433),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_491),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_511),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_491),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_503),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_510),
.Y(n_562)
);

INVx6_ASAP7_75t_L g563 ( 
.A(n_520),
.Y(n_563)
);

OAI21x1_ASAP7_75t_L g564 ( 
.A1(n_514),
.A2(n_452),
.B(n_465),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_533),
.A2(n_452),
.B(n_465),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_517),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g567 ( 
.A1(n_526),
.A2(n_444),
.B(n_464),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_509),
.B(n_454),
.Y(n_568)
);

NAND2x1p5_ASAP7_75t_L g569 ( 
.A(n_488),
.B(n_434),
.Y(n_569)
);

AO21x2_ASAP7_75t_L g570 ( 
.A1(n_492),
.A2(n_420),
.B(n_417),
.Y(n_570)
);

INVx8_ASAP7_75t_L g571 ( 
.A(n_512),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_529),
.Y(n_572)
);

AOI22x1_ASAP7_75t_L g573 ( 
.A1(n_523),
.A2(n_459),
.B1(n_460),
.B2(n_420),
.Y(n_573)
);

BUFx2_ASAP7_75t_SL g574 ( 
.A(n_506),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_537),
.B(n_422),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_515),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_485),
.Y(n_577)
);

BUFx12f_ASAP7_75t_L g578 ( 
.A(n_508),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_535),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_536),
.Y(n_580)
);

INVx5_ASAP7_75t_SL g581 ( 
.A(n_512),
.Y(n_581)
);

AO21x2_ASAP7_75t_L g582 ( 
.A1(n_498),
.A2(n_115),
.B(n_116),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_486),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_534),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_541),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_521),
.A2(n_118),
.B(n_120),
.Y(n_586)
);

BUFx5_ASAP7_75t_L g587 ( 
.A(n_539),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_525),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_483),
.B(n_121),
.Y(n_589)
);

CKINVDCx8_ASAP7_75t_R g590 ( 
.A(n_535),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_525),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_507),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_592),
.B(n_496),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_544),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_559),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_545),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_542),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_563),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_553),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_547),
.B(n_488),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_574),
.A2(n_484),
.B1(n_495),
.B2(n_505),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_546),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_561),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_545),
.B(n_496),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_549),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_548),
.A2(n_554),
.B(n_564),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_568),
.A2(n_528),
.B(n_518),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_543),
.Y(n_608)
);

NAND2x1p5_ASAP7_75t_L g609 ( 
.A(n_547),
.B(n_502),
.Y(n_609)
);

AO21x2_ASAP7_75t_L g610 ( 
.A1(n_550),
.A2(n_487),
.B(n_504),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_563),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_580),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_568),
.B(n_502),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_562),
.A2(n_500),
.B1(n_538),
.B2(n_527),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_562),
.B(n_522),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_590),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_558),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_585),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_576),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_588),
.Y(n_620)
);

NAND2x1p5_ASAP7_75t_L g621 ( 
.A(n_579),
.B(n_535),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_591),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_583),
.Y(n_623)
);

BUFx8_ASAP7_75t_SL g624 ( 
.A(n_572),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_557),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_584),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_557),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_583),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_586),
.Y(n_629)
);

INVx6_ASAP7_75t_L g630 ( 
.A(n_563),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_571),
.A2(n_540),
.B1(n_530),
.B2(n_524),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_577),
.B(n_158),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_555),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_558),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_577),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_558),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_555),
.Y(n_637)
);

CKINVDCx6p67_ASAP7_75t_R g638 ( 
.A(n_572),
.Y(n_638)
);

AND2x4_ASAP7_75t_SL g639 ( 
.A(n_638),
.B(n_566),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_608),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_R g641 ( 
.A(n_623),
.B(n_556),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_608),
.B(n_581),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_599),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_638),
.Y(n_644)
);

AO31x2_ASAP7_75t_L g645 ( 
.A1(n_629),
.A2(n_589),
.A3(n_575),
.B(n_587),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_601),
.A2(n_551),
.B1(n_581),
.B2(n_573),
.Y(n_646)
);

AND2x2_ASAP7_75t_SL g647 ( 
.A(n_631),
.B(n_581),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_599),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_R g649 ( 
.A(n_623),
.B(n_551),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_597),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_624),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_603),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_612),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_626),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_616),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_594),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_596),
.B(n_571),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_602),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_594),
.B(n_595),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_613),
.B(n_571),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_616),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_618),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_R g663 ( 
.A(n_628),
.B(n_556),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_595),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_602),
.Y(n_665)
);

AO31x2_ASAP7_75t_L g666 ( 
.A1(n_629),
.A2(n_589),
.A3(n_575),
.B(n_587),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_604),
.B(n_579),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_605),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_620),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_635),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_620),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_605),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_R g673 ( 
.A(n_628),
.B(n_578),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_619),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_619),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_617),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_630),
.B(n_551),
.Y(n_677)
);

OR2x6_ASAP7_75t_L g678 ( 
.A(n_630),
.B(n_560),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_622),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_613),
.B(n_560),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_593),
.B(n_560),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_598),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_598),
.B(n_570),
.Y(n_683)
);

AOI221xp5_ASAP7_75t_L g684 ( 
.A1(n_614),
.A2(n_607),
.B1(n_593),
.B2(n_615),
.C(n_627),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_600),
.B(n_570),
.Y(n_685)
);

NOR3xp33_ASAP7_75t_SL g686 ( 
.A(n_624),
.B(n_582),
.C(n_587),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_625),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_633),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_600),
.B(n_569),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_606),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_637),
.B(n_569),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_600),
.B(n_125),
.Y(n_692)
);

AOI222xp33_ASAP7_75t_L g693 ( 
.A1(n_632),
.A2(n_565),
.B1(n_567),
.B2(n_587),
.C1(n_552),
.C2(n_550),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_656),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_647),
.A2(n_609),
.B1(n_630),
.B2(n_598),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_656),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_650),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_669),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_654),
.B(n_670),
.Y(n_699)
);

AOI221xp5_ASAP7_75t_SL g700 ( 
.A1(n_646),
.A2(n_617),
.B1(n_634),
.B2(n_636),
.C(n_609),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_679),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_669),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_671),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_671),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_652),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_680),
.B(n_610),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_685),
.B(n_610),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_664),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_681),
.B(n_610),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_665),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_640),
.B(n_636),
.Y(n_711)
);

AOI33xp33_ASAP7_75t_L g712 ( 
.A1(n_684),
.A2(n_630),
.A3(n_582),
.B1(n_587),
.B2(n_552),
.B3(n_134),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_653),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_662),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_683),
.B(n_606),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_672),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_683),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_675),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_659),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_677),
.B(n_617),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_676),
.B(n_617),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_658),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_660),
.B(n_617),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_644),
.A2(n_611),
.B1(n_634),
.B2(n_636),
.Y(n_724)
);

INVxp67_ASAP7_75t_SL g725 ( 
.A(n_667),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_643),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_642),
.B(n_634),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_668),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_688),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_648),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_674),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_645),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_677),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_657),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_661),
.Y(n_735)
);

NAND3xp33_ASAP7_75t_SL g736 ( 
.A(n_641),
.B(n_611),
.C(n_621),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_729),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_725),
.B(n_689),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_699),
.B(n_661),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_715),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_694),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_697),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_701),
.B(n_655),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_694),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_712),
.B(n_693),
.C(n_686),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_705),
.Y(n_746)
);

AND2x4_ASAP7_75t_SL g747 ( 
.A(n_720),
.B(n_661),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_734),
.B(n_692),
.Y(n_748)
);

NAND3xp33_ASAP7_75t_L g749 ( 
.A(n_712),
.B(n_649),
.C(n_691),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_717),
.B(n_690),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_727),
.B(n_639),
.Y(n_751)
);

OA211x2_ASAP7_75t_L g752 ( 
.A1(n_736),
.A2(n_711),
.B(n_700),
.C(n_724),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_713),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_717),
.B(n_690),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_696),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_706),
.B(n_645),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_714),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_723),
.B(n_687),
.Y(n_758)
);

AND2x2_ASAP7_75t_SL g759 ( 
.A(n_733),
.B(n_682),
.Y(n_759)
);

NOR2xp67_ASAP7_75t_L g760 ( 
.A(n_717),
.B(n_707),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_706),
.B(n_666),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_735),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_708),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_727),
.B(n_651),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_723),
.B(n_682),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_708),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_696),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_737),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_740),
.B(n_709),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_740),
.B(n_709),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_746),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_741),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_737),
.B(n_707),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_746),
.B(n_698),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_741),
.Y(n_775)
);

AOI211xp5_ASAP7_75t_SL g776 ( 
.A1(n_740),
.A2(n_715),
.B(n_695),
.C(n_721),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_762),
.B(n_721),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_760),
.B(n_735),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_744),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_750),
.B(n_719),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_764),
.B(n_704),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_742),
.B(n_753),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_757),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_761),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_744),
.Y(n_785)
);

NAND2x1_ASAP7_75t_L g786 ( 
.A(n_750),
.B(n_704),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_767),
.B(n_698),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_745),
.A2(n_720),
.B1(n_733),
.B2(n_678),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_763),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_766),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_768),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_777),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_770),
.B(n_750),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_773),
.B(n_738),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_773),
.B(n_768),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_788),
.A2(n_749),
.B1(n_752),
.B2(n_759),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_771),
.Y(n_797)
);

INVx1_ASAP7_75t_SL g798 ( 
.A(n_781),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_774),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_769),
.B(n_748),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_772),
.Y(n_801)
);

OAI31xp33_ASAP7_75t_L g802 ( 
.A1(n_776),
.A2(n_756),
.A3(n_743),
.B(n_758),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_774),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_778),
.B(n_759),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_782),
.Y(n_805)
);

OAI21xp33_ASAP7_75t_SL g806 ( 
.A1(n_802),
.A2(n_782),
.B(n_784),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_796),
.A2(n_739),
.B(n_784),
.C(n_783),
.Y(n_807)
);

NAND4xp25_ASAP7_75t_L g808 ( 
.A(n_795),
.B(n_791),
.C(n_797),
.D(n_805),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_SL g809 ( 
.A1(n_798),
.A2(n_756),
.B1(n_770),
.B2(n_778),
.Y(n_809)
);

OAI22xp33_ASAP7_75t_L g810 ( 
.A1(n_794),
.A2(n_786),
.B1(n_733),
.B2(n_790),
.Y(n_810)
);

OAI21xp33_ASAP7_75t_L g811 ( 
.A1(n_799),
.A2(n_780),
.B(n_765),
.Y(n_811)
);

AOI32xp33_ASAP7_75t_L g812 ( 
.A1(n_806),
.A2(n_803),
.A3(n_792),
.B1(n_804),
.B2(n_780),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_808),
.B(n_800),
.Y(n_813)
);

NAND2x1p5_ASAP7_75t_L g814 ( 
.A(n_809),
.B(n_804),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_807),
.A2(n_793),
.B(n_789),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_810),
.A2(n_787),
.B(n_793),
.Y(n_816)
);

AO21x1_ASAP7_75t_SL g817 ( 
.A1(n_811),
.A2(n_787),
.B(n_663),
.Y(n_817)
);

NOR3x1_ASAP7_75t_L g818 ( 
.A(n_813),
.B(n_673),
.C(n_751),
.Y(n_818)
);

OAI21xp33_ASAP7_75t_L g819 ( 
.A1(n_812),
.A2(n_754),
.B(n_801),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_SL g820 ( 
.A(n_815),
.B(n_726),
.C(n_754),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_814),
.B(n_754),
.Y(n_821)
);

AOI211xp5_ASAP7_75t_L g822 ( 
.A1(n_816),
.A2(n_733),
.B(n_720),
.C(n_801),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_821),
.Y(n_823)
);

OA22x2_ASAP7_75t_L g824 ( 
.A1(n_819),
.A2(n_817),
.B1(n_747),
.B2(n_772),
.Y(n_824)
);

NAND4xp75_ASAP7_75t_L g825 ( 
.A(n_824),
.B(n_818),
.C(n_820),
.D(n_822),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_823),
.B(n_747),
.Y(n_826)
);

AOI221xp5_ASAP7_75t_L g827 ( 
.A1(n_823),
.A2(n_785),
.B1(n_779),
.B2(n_775),
.C(n_755),
.Y(n_827)
);

AO22x2_ASAP7_75t_L g828 ( 
.A1(n_825),
.A2(n_611),
.B1(n_755),
.B2(n_732),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_826),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_827),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_825),
.A2(n_730),
.B1(n_678),
.B2(n_732),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_826),
.B(n_703),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_829),
.B(n_127),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_R g834 ( 
.A(n_830),
.B(n_128),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_832),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_831),
.B(n_702),
.Y(n_836)
);

NAND4xp75_ASAP7_75t_L g837 ( 
.A(n_828),
.B(n_703),
.C(n_702),
.D(n_710),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_835),
.B(n_129),
.Y(n_838)
);

OA21x2_ASAP7_75t_L g839 ( 
.A1(n_833),
.A2(n_718),
.B(n_716),
.Y(n_839)
);

OAI211xp5_ASAP7_75t_SL g840 ( 
.A1(n_834),
.A2(n_131),
.B(n_136),
.C(n_137),
.Y(n_840)
);

NOR2x1_ASAP7_75t_L g841 ( 
.A(n_837),
.B(n_139),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_838),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_839),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_841),
.Y(n_844)
);

OAI22xp33_ASAP7_75t_L g845 ( 
.A1(n_840),
.A2(n_836),
.B1(n_716),
.B2(n_710),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_838),
.Y(n_846)
);

OAI22xp33_ASAP7_75t_L g847 ( 
.A1(n_844),
.A2(n_846),
.B1(n_842),
.B2(n_843),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_845),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_842),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_842),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_849),
.Y(n_851)
);

OAI22x1_ASAP7_75t_SL g852 ( 
.A1(n_850),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_851),
.B(n_848),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_853),
.B(n_847),
.C(n_852),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_854),
.A2(n_621),
.B1(n_718),
.B2(n_722),
.Y(n_855)
);

OR2x6_ASAP7_75t_L g856 ( 
.A(n_855),
.B(n_621),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_856),
.A2(n_731),
.B1(n_728),
.B2(n_722),
.Y(n_857)
);


endmodule