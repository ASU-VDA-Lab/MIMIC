module fake_jpeg_27458_n_225 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_118;
wire n_128;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_50),
.Y(n_71)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_32),
.Y(n_70)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_29),
.Y(n_49)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_0),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_24),
.B1(n_48),
.B2(n_41),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_60),
.B1(n_67),
.B2(n_77),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_24),
.B1(n_34),
.B2(n_28),
.Y(n_60)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_68),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_24),
.B1(n_32),
.B2(n_23),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_26),
.B1(n_20),
.B2(n_35),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_30),
.B1(n_25),
.B2(n_27),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_75),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_23),
.Y(n_73)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

CKINVDCx6p67_ASAP7_75t_R g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_25),
.B1(n_30),
.B2(n_18),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_79),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_46),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_84),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_27),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_15),
.C(n_14),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_44),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_95),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_45),
.B1(n_62),
.B2(n_28),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_93),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_98),
.Y(n_127)
);

OR2x2_ASAP7_75t_SL g98 ( 
.A(n_54),
.B(n_35),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_63),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_99),
.Y(n_130)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g112 ( 
.A(n_100),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_22),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_53),
.A2(n_29),
.A3(n_49),
.B1(n_26),
.B2(n_28),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_62),
.B1(n_45),
.B2(n_56),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_75),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_57),
.B(n_47),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_55),
.Y(n_120)
);

OAI22x1_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_34),
.B1(n_29),
.B2(n_61),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_114),
.B1(n_129),
.B2(n_94),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_64),
.B(n_56),
.C(n_53),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_83),
.B(n_80),
.Y(n_145)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_123),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_128),
.B1(n_88),
.B2(n_105),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_34),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_22),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_81),
.A2(n_22),
.B1(n_29),
.B2(n_3),
.Y(n_128)
);

OAI22x1_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_79),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_140),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_143),
.B1(n_108),
.B2(n_131),
.Y(n_158)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_137),
.Y(n_154)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_98),
.B(n_96),
.Y(n_138)
);

OA21x2_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_129),
.B(n_121),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_106),
.B1(n_89),
.B2(n_82),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_109),
.B1(n_126),
.B2(n_110),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_107),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_130),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_142),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_130),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_150),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_146),
.B(n_113),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_83),
.B(n_90),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_103),
.C(n_90),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_122),
.C(n_111),
.Y(n_156)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_120),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_80),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_153),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_166),
.C(n_167),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_140),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_168),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_110),
.B1(n_128),
.B2(n_131),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_123),
.C(n_125),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_113),
.C(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_136),
.B(n_152),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_169),
.B(n_171),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_145),
.B(n_132),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_112),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_159),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_178),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_176),
.A2(n_162),
.B1(n_160),
.B2(n_165),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_163),
.B(n_141),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_15),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_133),
.C(n_132),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_184),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_150),
.B(n_139),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_169),
.B(n_146),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_143),
.C(n_134),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_167),
.C(n_161),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_192),
.C(n_173),
.Y(n_201)
);

OAI31xp33_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_160),
.A3(n_162),
.B(n_164),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_SL g203 ( 
.A1(n_193),
.A2(n_184),
.B(n_182),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_163),
.B1(n_154),
.B2(n_171),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_180),
.C(n_10),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_155),
.B1(n_149),
.B2(n_135),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_186),
.B1(n_149),
.B2(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_189),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_188),
.A2(n_177),
.B1(n_187),
.B2(n_176),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_205),
.Y(n_212)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_198),
.B(n_194),
.Y(n_210)
);

INVxp33_ASAP7_75t_SL g204 ( 
.A(n_193),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_206),
.B(n_196),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_180),
.C(n_173),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_189),
.C(n_191),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_208),
.C(n_80),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_210),
.A2(n_198),
.B1(n_203),
.B2(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_214),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_137),
.A3(n_112),
.B1(n_12),
.B2(n_6),
.C1(n_7),
.C2(n_2),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_217),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_100),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_209),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_207),
.C(n_212),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_222),
.B(n_219),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_218),
.A2(n_208),
.B1(n_5),
.B2(n_6),
.Y(n_222)
);

AOI222xp33_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.C1(n_80),
.C2(n_141),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_224),
.Y(n_225)
);


endmodule