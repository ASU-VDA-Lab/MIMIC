module fake_jpeg_20684_n_277 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

AND2x4_ASAP7_75t_SL g36 ( 
.A(n_22),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_28),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_20),
.B1(n_17),
.B2(n_25),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_44),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_17),
.B1(n_25),
.B2(n_26),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_40),
.B1(n_23),
.B2(n_29),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_17),
.B1(n_25),
.B2(n_18),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_26),
.B1(n_21),
.B2(n_31),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_26),
.B1(n_24),
.B2(n_31),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_16),
.B1(n_21),
.B2(n_33),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_62),
.B1(n_40),
.B2(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_43),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_34),
.A2(n_16),
.B1(n_33),
.B2(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_73),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_24),
.B1(n_32),
.B2(n_23),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_38),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_74),
.B(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_85),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_82),
.B1(n_84),
.B2(n_19),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_78),
.B(n_86),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_29),
.B(n_23),
.C(n_43),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_43),
.B(n_35),
.C(n_63),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_27),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_46),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_38),
.B1(n_42),
.B2(n_19),
.Y(n_84)
);

CKINVDCx6p67_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_89),
.Y(n_111)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_29),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_98),
.Y(n_118)
);

OR2x4_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_79),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_78),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_28),
.Y(n_98)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_51),
.B1(n_46),
.B2(n_48),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_43),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_106),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_56),
.B1(n_52),
.B2(n_58),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_104),
.A2(n_110),
.B1(n_85),
.B2(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_83),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_30),
.C(n_28),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_84),
.C(n_69),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_42),
.B1(n_63),
.B2(n_30),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_114),
.B1(n_115),
.B2(n_99),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_27),
.B(n_1),
.C(n_2),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_75),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_122),
.B(n_135),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_81),
.Y(n_123)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_124),
.B(n_100),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_4),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_87),
.B1(n_65),
.B2(n_76),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_131),
.B1(n_112),
.B2(n_114),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_64),
.C(n_80),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_98),
.C(n_108),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_130),
.B(n_0),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_82),
.B1(n_85),
.B2(n_80),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_72),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_111),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_113),
.B(n_9),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_137),
.A2(n_102),
.B1(n_106),
.B2(n_91),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_72),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_138),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_27),
.B1(n_8),
.B2(n_10),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_113),
.B(n_115),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_160),
.B(n_162),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_157),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_152),
.B1(n_153),
.B2(n_133),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_92),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_155),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_163),
.B1(n_131),
.B2(n_123),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_151),
.A2(n_154),
.B(n_156),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_107),
.B1(n_101),
.B2(n_100),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_109),
.B1(n_2),
.B2(n_3),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_109),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_109),
.C(n_7),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_0),
.B(n_2),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_2),
.B(n_3),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_139),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_11),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_177),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_145),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_170),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_171),
.A2(n_181),
.B1(n_153),
.B2(n_158),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_187),
.B1(n_163),
.B2(n_142),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_123),
.B(n_124),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_189),
.B(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_142),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_117),
.Y(n_179)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_122),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_127),
.B1(n_121),
.B2(n_136),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_118),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_186),
.C(n_165),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_135),
.B(n_140),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_166),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_139),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_129),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_146),
.A2(n_139),
.B1(n_5),
.B2(n_6),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_181),
.C(n_175),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_194),
.C(n_197),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_172),
.C(n_186),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_184),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_195),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_147),
.C(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_167),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_201),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_157),
.C(n_141),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_210),
.C(n_168),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_205),
.B(n_189),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_173),
.B1(n_187),
.B2(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_209),
.A2(n_171),
.B1(n_174),
.B2(n_169),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_216),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_218),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_199),
.A2(n_174),
.B1(n_185),
.B2(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

BUFx12_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_201),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_192),
.Y(n_231)
);

AOI221xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_169),
.B1(n_183),
.B2(n_160),
.C(n_162),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_226),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_188),
.C(n_155),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_203),
.C(n_210),
.Y(n_227)
);

AOI221xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_164),
.B1(n_178),
.B2(n_150),
.C(n_177),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_231),
.C(n_219),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_202),
.B(n_199),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_229),
.B(n_234),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_197),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_237),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_236),
.B(n_214),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_195),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_211),
.B(n_164),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_238),
.B(n_225),
.CI(n_213),
.CON(n_244),
.SN(n_244)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_191),
.B1(n_200),
.B2(n_193),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_216),
.B1(n_222),
.B2(n_215),
.Y(n_245)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_230),
.A2(n_221),
.B1(n_217),
.B2(n_191),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_244),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_218),
.Y(n_243)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_212),
.B1(n_198),
.B2(n_215),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_248),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_238),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_257),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_233),
.C(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_254),
.B(n_248),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_245),
.A2(n_232),
.B(n_214),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_246),
.A2(n_235),
.B(n_207),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_262),
.C(n_263),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_244),
.C(n_240),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_244),
.C(n_246),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_251),
.B(n_218),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_11),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_265),
.A2(n_253),
.A3(n_249),
.B1(n_252),
.B2(n_256),
.C1(n_258),
.C2(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_267),
.Y(n_271)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_261),
.A3(n_259),
.B1(n_255),
.B2(n_198),
.C1(n_247),
.C2(n_178),
.Y(n_267)
);

AOI31xp67_ASAP7_75t_SL g268 ( 
.A1(n_263),
.A2(n_11),
.A3(n_13),
.B(n_12),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_12),
.C(n_14),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_272),
.B(n_271),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.C(n_4),
.Y(n_276)
);

AOI321xp33_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_270),
.A3(n_10),
.B1(n_13),
.B2(n_5),
.C(n_6),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_5),
.Y(n_277)
);


endmodule