module fake_jpeg_4460_n_176 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_22),
.Y(n_46)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

HAxp5_ASAP7_75t_SL g37 ( 
.A(n_14),
.B(n_7),
.CON(n_37),
.SN(n_37)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_17),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_28),
.A2(n_13),
.B1(n_26),
.B2(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_50),
.B1(n_20),
.B2(n_19),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_13),
.B1(n_18),
.B2(n_14),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_13),
.B1(n_23),
.B2(n_14),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_27),
.B1(n_25),
.B2(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_24),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_68),
.B1(n_25),
.B2(n_20),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_64),
.C(n_61),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_57),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_60),
.B(n_27),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_33),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_18),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_19),
.B1(n_20),
.B2(n_25),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_18),
.B1(n_21),
.B2(n_27),
.Y(n_68)
);

INVxp33_ASAP7_75t_SL g69 ( 
.A(n_54),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_78),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_80),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_40),
.B(n_33),
.C(n_29),
.D(n_42),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_76),
.C(n_19),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_40),
.A3(n_42),
.B1(n_39),
.B2(n_38),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_48),
.B1(n_53),
.B2(n_44),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_41),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_88),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_93),
.B1(n_87),
.B2(n_92),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_39),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_96),
.B(n_85),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_44),
.B(n_66),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_66),
.B(n_38),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_41),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_59),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_100),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_115),
.B1(n_116),
.B2(n_95),
.Y(n_124)
);

AO22x1_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_74),
.B1(n_76),
.B2(n_73),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_114),
.B(n_96),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_108),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_111),
.Y(n_120)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_79),
.B1(n_38),
.B2(n_15),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_117),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_47),
.B1(n_62),
.B2(n_16),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_62),
.B1(n_24),
.B2(n_16),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_91),
.C(n_94),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_122),
.C(n_113),
.Y(n_137)
);

AO221x1_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_75),
.B1(n_65),
.B2(n_92),
.C(n_15),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_124),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_126),
.A2(n_114),
.B(n_110),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_90),
.A3(n_98),
.B1(n_89),
.B2(n_86),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_131),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_75),
.Y(n_131)
);

OA21x2_ASAP7_75t_SL g132 ( 
.A1(n_127),
.A2(n_103),
.B(n_108),
.Y(n_132)
);

AOI31xp67_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_122),
.A3(n_119),
.B(n_128),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_142),
.B(n_123),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_90),
.B1(n_107),
.B2(n_104),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_134),
.A2(n_143),
.B1(n_15),
.B2(n_125),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_139),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_38),
.C(n_65),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_65),
.C(n_15),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_129),
.Y(n_145)
);

AOI21x1_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_65),
.B(n_15),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_24),
.B1(n_15),
.B2(n_22),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_151),
.B1(n_150),
.B2(n_22),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_147),
.B(n_151),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_124),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_146),
.A2(n_149),
.B(n_152),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_134),
.B1(n_143),
.B2(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_0),
.B(n_1),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_139),
.C(n_137),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_0),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_152),
.A2(n_136),
.B(n_135),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_158),
.B(n_160),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_157),
.B(n_159),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_147),
.A2(n_141),
.B(n_1),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_22),
.C(n_0),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_9),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_155),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_162),
.A2(n_163),
.B(n_166),
.C(n_10),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_158),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_165),
.C(n_160),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_10),
.B(n_11),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_9),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_10),
.B(n_11),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_173),
.C(n_170),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_12),
.C(n_167),
.Y(n_175)
);


endmodule