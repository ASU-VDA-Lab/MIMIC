module fake_jpeg_28680_n_363 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_363);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_363;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_50),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g128 ( 
.A(n_51),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_61),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_25),
.B(n_8),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_64),
.B(n_68),
.Y(n_114)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_25),
.B(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_74),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_26),
.B(n_15),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g141 ( 
.A(n_76),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_80),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_SL g79 ( 
.A(n_30),
.B(n_14),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_81),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_24),
.B(n_13),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_87),
.Y(n_125)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_86),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_26),
.B(n_13),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_89),
.Y(n_132)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_91),
.Y(n_127)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_93),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_27),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_47),
.C(n_35),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_96),
.A2(n_27),
.B(n_1),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_34),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_99),
.B(n_100),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_34),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_105),
.B(n_119),
.Y(n_190)
);

CKINVDCx11_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_109),
.B(n_123),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_17),
.B1(n_29),
.B2(n_47),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_110),
.A2(n_115),
.B1(n_118),
.B2(n_148),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_29),
.B1(n_38),
.B2(n_40),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_48),
.A2(n_40),
.B1(n_38),
.B2(n_35),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_55),
.B(n_44),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_50),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_46),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_138),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_86),
.B(n_44),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_140),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_93),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_90),
.A2(n_46),
.B1(n_43),
.B2(n_33),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_52),
.B(n_43),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_149),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_58),
.A2(n_33),
.B1(n_45),
.B2(n_28),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_60),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_69),
.B(n_34),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_100),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_103),
.A2(n_88),
.B1(n_84),
.B2(n_78),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_151),
.A2(n_161),
.B1(n_165),
.B2(n_168),
.Y(n_226)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_137),
.A2(n_75),
.B1(n_73),
.B2(n_72),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_155),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_103),
.A2(n_45),
.B1(n_28),
.B2(n_19),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_156),
.A2(n_180),
.B1(n_182),
.B2(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_99),
.A2(n_19),
.B1(n_11),
.B2(n_9),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_185),
.Y(n_202)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_27),
.B1(n_9),
.B2(n_2),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_167),
.Y(n_225)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_0),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_112),
.C(n_98),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_170),
.B(n_128),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_27),
.B(n_1),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_107),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_174),
.B(n_183),
.Y(n_233)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_184),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_132),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_126),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_126),
.A2(n_133),
.B1(n_145),
.B2(n_135),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_114),
.B(n_3),
.Y(n_183)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_96),
.B(n_4),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_189),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_121),
.B(n_5),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_134),
.B(n_5),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_156),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_104),
.A2(n_5),
.B1(n_129),
.B2(n_111),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_192),
.A2(n_143),
.B1(n_131),
.B2(n_141),
.Y(n_231)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_97),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_194),
.Y(n_229)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_144),
.A2(n_101),
.B1(n_132),
.B2(n_95),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_136),
.A3(n_101),
.B1(n_116),
.B2(n_98),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_127),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_196),
.B(n_95),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_133),
.A2(n_145),
.B1(n_102),
.B2(n_135),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_147),
.B(n_191),
.C(n_195),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_227),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_141),
.B(n_147),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_204),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_200),
.B(n_201),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_175),
.B(n_130),
.Y(n_201)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_174),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_212),
.Y(n_242)
);

AOI32xp33_ASAP7_75t_L g212 ( 
.A1(n_176),
.A2(n_181),
.A3(n_159),
.B1(n_163),
.B2(n_169),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_228),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_166),
.A2(n_104),
.B1(n_129),
.B2(n_116),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_195),
.A2(n_102),
.B1(n_124),
.B2(n_117),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_222),
.A2(n_231),
.B1(n_167),
.B2(n_195),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_124),
.C(n_141),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_169),
.Y(n_246)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_238),
.Y(n_263)
);

INVx11_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_247),
.Y(n_268)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_245),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_248),
.B1(n_254),
.B2(n_255),
.Y(n_267)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_246),
.B(n_228),
.Y(n_271)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_216),
.A2(n_185),
.B1(n_157),
.B2(n_155),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_166),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_258),
.Y(n_274)
);

AND2x2_ASAP7_75t_SL g250 ( 
.A(n_202),
.B(n_170),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_200),
.B(n_190),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_253),
.B(n_260),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_216),
.A2(n_187),
.B1(n_168),
.B2(n_184),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_199),
.A2(n_179),
.B1(n_153),
.B2(n_158),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_198),
.A2(n_178),
.B1(n_173),
.B2(n_162),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_261),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_212),
.A2(n_164),
.B1(n_188),
.B2(n_193),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_171),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_214),
.A2(n_116),
.B1(n_177),
.B2(n_152),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_201),
.B(n_128),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_214),
.A2(n_194),
.B1(n_143),
.B2(n_131),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_128),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_258),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_237),
.A2(n_230),
.B1(n_227),
.B2(n_220),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_264),
.A2(n_265),
.B1(n_281),
.B2(n_255),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_230),
.B1(n_204),
.B2(n_220),
.Y(n_265)
);

OAI32xp33_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_226),
.A3(n_217),
.B1(n_232),
.B2(n_233),
.Y(n_266)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_219),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_270),
.A2(n_278),
.B(n_283),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_272),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_252),
.B(n_246),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_240),
.A2(n_229),
.B(n_208),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_240),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_279),
.A2(n_256),
.B1(n_236),
.B2(n_257),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_262),
.A2(n_210),
.B1(n_211),
.B2(n_218),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_251),
.B(n_215),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_259),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_239),
.A2(n_223),
.B(n_218),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_251),
.B(n_225),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_252),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_284),
.C(n_280),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_289),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_300),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_279),
.A2(n_239),
.B1(n_250),
.B2(n_242),
.Y(n_289)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_263),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_278),
.A2(n_239),
.B(n_250),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_302),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_265),
.A2(n_234),
.B1(n_235),
.B2(n_261),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_298),
.Y(n_316)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_283),
.A2(n_239),
.B1(n_243),
.B2(n_245),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_301),
.A2(n_303),
.B(n_263),
.Y(n_317)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_270),
.A2(n_247),
.B(n_238),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_275),
.B(n_213),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_285),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_286),
.B(n_271),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_308),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_270),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_310),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_274),
.Y(n_310)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_311),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_274),
.C(n_264),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_312),
.B(n_313),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_296),
.C(n_303),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_266),
.C(n_281),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_288),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_317),
.A2(n_294),
.B(n_298),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_306),
.A2(n_291),
.B1(n_287),
.B2(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_314),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_326),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_325),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_319),
.A2(n_291),
.B1(n_294),
.B2(n_267),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_327),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_315),
.B(n_316),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_295),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_318),
.A2(n_293),
.B1(n_290),
.B2(n_267),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_330),
.A2(n_312),
.B1(n_309),
.B2(n_277),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_282),
.Y(n_334)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_304),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_324),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_337),
.B(n_320),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_325),
.A2(n_277),
.B(n_275),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_338),
.A2(n_327),
.B(n_323),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_307),
.C(n_308),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_340),
.B(n_321),
.C(n_329),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_341),
.B(n_337),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_329),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_335),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_347),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_345),
.A2(n_338),
.B(n_335),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_333),
.A2(n_326),
.B(n_302),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_346),
.A2(n_340),
.B(n_339),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_351),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_350),
.A2(n_352),
.B(n_345),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_349),
.A2(n_344),
.B1(n_332),
.B2(n_339),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_353),
.B(n_355),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_354),
.A2(n_332),
.B1(n_343),
.B2(n_350),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_357),
.B(n_321),
.Y(n_359)
);

AOI31xp33_ASAP7_75t_L g358 ( 
.A1(n_356),
.A2(n_300),
.A3(n_341),
.B(n_276),
.Y(n_358)
);

NAND3xp33_ASAP7_75t_L g360 ( 
.A(n_358),
.B(n_359),
.C(n_276),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_360),
.A2(n_268),
.B1(n_241),
.B2(n_213),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_213),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_362),
.B(n_310),
.Y(n_363)
);


endmodule