module fake_netlist_1_9207_n_710 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_710);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_710;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_466;
wire n_302;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_57), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_50), .Y(n_83) );
HB1xp67_ASAP7_75t_L g84 ( .A(n_67), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_18), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_33), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_55), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_21), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_45), .Y(n_89) );
CKINVDCx14_ASAP7_75t_R g90 ( .A(n_2), .Y(n_90) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_78), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_53), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_47), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_74), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_72), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_62), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_70), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_0), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_2), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_68), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_80), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_81), .B(n_56), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_6), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_41), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_22), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_35), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_8), .B(n_7), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_49), .Y(n_108) );
INVx3_ASAP7_75t_L g109 ( .A(n_61), .Y(n_109) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_28), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_30), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_26), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_51), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_59), .Y(n_114) );
INVxp33_ASAP7_75t_L g115 ( .A(n_16), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_58), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_16), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_29), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_11), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_77), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_64), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_27), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_75), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_69), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_79), .Y(n_125) );
INVxp67_ASAP7_75t_SL g126 ( .A(n_5), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_32), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_48), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_24), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_31), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_39), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_90), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_109), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_109), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_98), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_87), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_84), .B(n_0), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_91), .B(n_1), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_131), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_96), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_98), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_98), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_115), .B(n_1), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_94), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_110), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_82), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_86), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_109), .B(n_3), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_109), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_85), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_122), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_122), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_104), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_122), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_82), .Y(n_155) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_83), .A2(n_34), .B(n_73), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_106), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_83), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_85), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_89), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_89), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_93), .Y(n_162) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_93), .A2(n_25), .B(n_71), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_95), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_123), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_95), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_88), .Y(n_167) );
INVxp67_ASAP7_75t_SL g168 ( .A(n_117), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_97), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g170 ( .A(n_97), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_117), .B(n_3), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_100), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_100), .B(n_4), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_101), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_101), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_105), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_147), .Y(n_179) );
NAND3xp33_ASAP7_75t_L g180 ( .A(n_150), .B(n_88), .C(n_92), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_133), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_167), .B(n_92), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_133), .Y(n_184) );
NOR2xp33_ASAP7_75t_SL g185 ( .A(n_170), .B(n_125), .Y(n_185) );
INVxp67_ASAP7_75t_L g186 ( .A(n_143), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_168), .B(n_125), .Y(n_187) );
BUFx6f_ASAP7_75t_SL g188 ( .A(n_155), .Y(n_188) );
AO22x2_ASAP7_75t_L g189 ( .A1(n_148), .A2(n_130), .B1(n_129), .B2(n_128), .Y(n_189) );
INVx4_ASAP7_75t_SL g190 ( .A(n_133), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_173), .A2(n_99), .B1(n_103), .B2(n_119), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_168), .B(n_130), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_140), .B(n_129), .Y(n_193) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_153), .Y(n_194) );
AO22x2_ASAP7_75t_L g195 ( .A1(n_173), .A2(n_128), .B1(n_127), .B2(n_114), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_133), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_134), .Y(n_197) );
INVxp67_ASAP7_75t_L g198 ( .A(n_143), .Y(n_198) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_150), .B(n_173), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_134), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_133), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_133), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_161), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_145), .B(n_127), .Y(n_206) );
OR2x2_ASAP7_75t_L g207 ( .A(n_170), .B(n_126), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_149), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_171), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_146), .B(n_124), .Y(n_210) );
NAND2x1p5_ASAP7_75t_L g211 ( .A(n_171), .B(n_124), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_155), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_149), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_161), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_146), .B(n_113), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_171), .B(n_113), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_149), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_164), .B(n_105), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_161), .Y(n_219) );
OAI221xp5_ASAP7_75t_L g220 ( .A1(n_137), .A2(n_107), .B1(n_112), .B2(n_118), .C(n_121), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_139), .Y(n_221) );
NAND3xp33_ASAP7_75t_L g222 ( .A(n_137), .B(n_120), .C(n_116), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_136), .Y(n_223) );
OAI21xp33_ASAP7_75t_L g224 ( .A1(n_164), .A2(n_120), .B(n_116), .Y(n_224) );
BUFx3_ASAP7_75t_L g225 ( .A(n_165), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_161), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_161), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_176), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_161), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_161), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_176), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_166), .B(n_114), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_176), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_176), .Y(n_234) );
INVx1_ASAP7_75t_SL g235 ( .A(n_144), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_166), .B(n_111), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_155), .A2(n_111), .B1(n_108), .B2(n_102), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_176), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_172), .B(n_108), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_176), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_158), .Y(n_241) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_132), .Y(n_242) );
INVx4_ASAP7_75t_L g243 ( .A(n_188), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_183), .B(n_175), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_177), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_201), .B(n_175), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_201), .B(n_172), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_201), .B(n_138), .Y(n_248) );
NOR3xp33_ASAP7_75t_SL g249 ( .A(n_221), .B(n_159), .C(n_141), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_177), .Y(n_250) );
INVxp67_ASAP7_75t_L g251 ( .A(n_235), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_178), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_185), .A2(n_160), .B1(n_174), .B2(n_169), .Y(n_253) );
INVxp67_ASAP7_75t_L g254 ( .A(n_179), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_186), .B(n_160), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_197), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_200), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_209), .A2(n_160), .B(n_174), .C(n_169), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_207), .B(n_174), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_178), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_178), .B(n_169), .Y(n_261) );
OR2x6_ASAP7_75t_L g262 ( .A(n_211), .B(n_163), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_221), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_181), .Y(n_264) );
INVx4_ASAP7_75t_L g265 ( .A(n_188), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_197), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_202), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_202), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_181), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_181), .Y(n_270) );
NOR2xp33_ASAP7_75t_R g271 ( .A(n_223), .B(n_188), .Y(n_271) );
INVx5_ASAP7_75t_L g272 ( .A(n_212), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_211), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_212), .B(n_176), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_211), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_208), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_223), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_189), .Y(n_278) );
NAND2x1p5_ASAP7_75t_L g279 ( .A(n_225), .B(n_162), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_198), .B(n_162), .Y(n_280) );
NOR2xp33_ASAP7_75t_R g281 ( .A(n_225), .B(n_135), .Y(n_281) );
INVxp67_ASAP7_75t_L g282 ( .A(n_194), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_199), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_216), .B(n_162), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_187), .B(n_163), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_189), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_189), .A2(n_158), .B1(n_152), .B2(n_151), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_208), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_189), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_195), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_213), .Y(n_291) );
INVxp67_ASAP7_75t_SL g292 ( .A(n_212), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_207), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_187), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_213), .Y(n_295) );
AO22x1_ASAP7_75t_L g296 ( .A1(n_242), .A2(n_158), .B1(n_135), .B2(n_141), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_192), .B(n_142), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_217), .Y(n_298) );
BUFx4f_ASAP7_75t_L g299 ( .A(n_187), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_217), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g301 ( .A1(n_216), .A2(n_154), .B(n_152), .C(n_151), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_200), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_195), .Y(n_303) );
NOR2xp33_ASAP7_75t_R g304 ( .A(n_193), .B(n_206), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_192), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_191), .Y(n_306) );
NAND2xp33_ASAP7_75t_R g307 ( .A(n_192), .B(n_156), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_195), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_210), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_190), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_190), .Y(n_311) );
BUFx8_ASAP7_75t_L g312 ( .A(n_210), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_218), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_286), .A2(n_195), .B1(n_210), .B2(n_215), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_276), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_276), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_290), .A2(n_215), .B1(n_222), .B2(n_220), .Y(n_317) );
AOI22xp33_ASAP7_75t_SL g318 ( .A1(n_312), .A2(n_313), .B1(n_281), .B2(n_271), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_312), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_312), .Y(n_320) );
INVx5_ASAP7_75t_L g321 ( .A(n_243), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_261), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_285), .A2(n_215), .B(n_232), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
CKINVDCx16_ASAP7_75t_R g325 ( .A(n_271), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_285), .A2(n_236), .B(n_156), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_301), .A2(n_224), .B(n_241), .C(n_239), .Y(n_327) );
NAND2x1p5_ASAP7_75t_L g328 ( .A(n_273), .B(n_239), .Y(n_328) );
INVx2_ASAP7_75t_SL g329 ( .A(n_275), .Y(n_329) );
AND3x1_ASAP7_75t_SL g330 ( .A(n_293), .B(n_142), .C(n_5), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_272), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_246), .B(n_218), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_278), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_308), .A2(n_180), .B1(n_237), .B2(n_151), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_285), .A2(n_262), .B(n_244), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_291), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_309), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_269), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_289), .A2(n_152), .B1(n_154), .B2(n_228), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g340 ( .A(n_249), .B(n_251), .C(n_263), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_246), .B(n_154), .Y(n_341) );
NOR2x1_ASAP7_75t_L g342 ( .A(n_259), .B(n_228), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_262), .A2(n_156), .B(n_204), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_246), .B(n_190), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_291), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_254), .B(n_4), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_262), .A2(n_156), .B(n_204), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_247), .B(n_163), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_306), .A2(n_219), .B1(n_238), .B2(n_227), .C(n_229), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_245), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_247), .B(n_156), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_247), .B(n_190), .Y(n_352) );
NAND2x2_ASAP7_75t_L g353 ( .A(n_263), .B(n_6), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_303), .A2(n_203), .B1(n_196), .B2(n_184), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_313), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_299), .A2(n_203), .B1(n_196), .B2(n_184), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_299), .A2(n_182), .B1(n_238), .B2(n_227), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_269), .B(n_7), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_244), .B(n_8), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_272), .B(n_182), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_272), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_283), .B(n_9), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_279), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_248), .A2(n_182), .B1(n_229), .B2(n_219), .Y(n_364) );
NOR2x1_ASAP7_75t_L g365 ( .A(n_248), .B(n_230), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_279), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_294), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_255), .B(n_9), .Y(n_368) );
INVx4_ASAP7_75t_L g369 ( .A(n_243), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_293), .Y(n_370) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_319), .B(n_243), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_350), .Y(n_372) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_314), .A2(n_305), .B1(n_277), .B2(n_282), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_329), .B(n_252), .Y(n_374) );
BUFx4f_ASAP7_75t_SL g375 ( .A(n_319), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_328), .Y(n_376) );
NAND3xp33_ASAP7_75t_SL g377 ( .A(n_318), .B(n_304), .C(n_287), .Y(n_377) );
INVxp67_ASAP7_75t_L g378 ( .A(n_370), .Y(n_378) );
INVx4_ASAP7_75t_L g379 ( .A(n_321), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_328), .B(n_284), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_324), .B(n_265), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_358), .A2(n_248), .B1(n_304), .B2(n_260), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_367), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_328), .B(n_280), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_322), .B(n_284), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_355), .A2(n_265), .B1(n_297), .B2(n_253), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_368), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_350), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_368), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_329), .B(n_245), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_358), .A2(n_270), .B1(n_264), .B2(n_300), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_331), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_332), .B(n_250), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_324), .A2(n_265), .B1(n_307), .B2(n_250), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_358), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_370), .A2(n_296), .B1(n_258), .B2(n_301), .C(n_295), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_320), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_320), .B(n_256), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g399 ( .A1(n_317), .A2(n_292), .B(n_307), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_337), .A2(n_266), .B1(n_256), .B2(n_267), .Y(n_400) );
NAND2xp33_ASAP7_75t_R g401 ( .A(n_362), .B(n_298), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_362), .B(n_298), .Y(n_402) );
AO31x2_ASAP7_75t_L g403 ( .A1(n_326), .A2(n_268), .A3(n_266), .B(n_288), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_315), .Y(n_404) );
OR2x6_ASAP7_75t_L g405 ( .A(n_335), .B(n_267), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_315), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_380), .B(n_268), .Y(n_407) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_401), .A2(n_359), .B(n_327), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_382), .A2(n_323), .B1(n_366), .B2(n_363), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_388), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
INVxp33_ASAP7_75t_L g412 ( .A(n_397), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_380), .B(n_288), .Y(n_413) );
OA21x2_ASAP7_75t_L g414 ( .A1(n_399), .A2(n_347), .B(n_343), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_402), .B(n_337), .Y(n_415) );
OAI211xp5_ASAP7_75t_SL g416 ( .A1(n_378), .A2(n_340), .B(n_346), .C(n_365), .Y(n_416) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_396), .B(n_351), .C(n_348), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_376), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_377), .A2(n_353), .B1(n_334), .B2(n_333), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_373), .A2(n_353), .B1(n_333), .B2(n_348), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_390), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_385), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_372), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_402), .A2(n_330), .B1(n_325), .B2(n_363), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_388), .Y(n_425) );
OAI211xp5_ASAP7_75t_L g426 ( .A1(n_384), .A2(n_369), .B(n_341), .C(n_321), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_379), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_385), .B(n_345), .Y(n_428) );
OAI21xp33_ASAP7_75t_SL g429 ( .A1(n_405), .A2(n_351), .B(n_366), .Y(n_429) );
OAI22xp33_ASAP7_75t_SL g430 ( .A1(n_405), .A2(n_369), .B1(n_321), .B2(n_336), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_379), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_387), .A2(n_336), .B1(n_345), .B2(n_369), .Y(n_432) );
OAI21x1_ASAP7_75t_L g433 ( .A1(n_389), .A2(n_360), .B(n_342), .Y(n_433) );
AOI222xp33_ASAP7_75t_L g434 ( .A1(n_375), .A2(n_338), .B1(n_349), .B2(n_321), .C1(n_339), .C2(n_316), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_391), .A2(n_316), .B1(n_336), .B2(n_345), .Y(n_435) );
OAI22xp33_ASAP7_75t_L g436 ( .A1(n_395), .A2(n_321), .B1(n_331), .B2(n_361), .Y(n_436) );
AOI222xp33_ASAP7_75t_L g437 ( .A1(n_422), .A2(n_383), .B1(n_397), .B2(n_386), .C1(n_393), .C2(n_398), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_420), .A2(n_400), .B1(n_405), .B2(n_371), .C(n_381), .Y(n_438) );
AOI21xp33_ASAP7_75t_L g439 ( .A1(n_424), .A2(n_405), .B(n_394), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_410), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_423), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_427), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_424), .A2(n_390), .B1(n_372), .B2(n_398), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_410), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_410), .Y(n_445) );
BUFx3_ASAP7_75t_L g446 ( .A(n_427), .Y(n_446) );
OR2x6_ASAP7_75t_L g447 ( .A(n_411), .B(n_379), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_407), .B(n_406), .Y(n_448) );
OAI221xp5_ASAP7_75t_SL g449 ( .A1(n_419), .A2(n_393), .B1(n_364), .B2(n_404), .C(n_406), .Y(n_449) );
AND4x1_ASAP7_75t_L g450 ( .A(n_434), .B(n_404), .C(n_11), .D(n_12), .Y(n_450) );
INVx2_ASAP7_75t_SL g451 ( .A(n_427), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_425), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_422), .A2(n_398), .B1(n_374), .B2(n_392), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_425), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_407), .B(n_392), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_423), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_425), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_431), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_413), .A2(n_374), .B1(n_331), .B2(n_361), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_421), .A2(n_374), .B1(n_331), .B2(n_354), .Y(n_460) );
BUFx2_ASAP7_75t_L g461 ( .A(n_429), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_431), .Y(n_462) );
AO21x1_ASAP7_75t_SL g463 ( .A1(n_429), .A2(n_344), .B(n_403), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_421), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_413), .B(n_403), .Y(n_465) );
NAND2xp33_ASAP7_75t_SL g466 ( .A(n_412), .B(n_331), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_430), .A2(n_360), .B(n_274), .Y(n_467) );
OAI21x1_ASAP7_75t_L g468 ( .A1(n_414), .A2(n_433), .B(n_435), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_415), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_433), .Y(n_470) );
OA222x2_ASAP7_75t_L g471 ( .A1(n_431), .A2(n_403), .B1(n_12), .B2(n_13), .C1(n_14), .C2(n_15), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_433), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_430), .A2(n_274), .B(n_356), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_441), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_442), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_465), .B(n_418), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_441), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_452), .Y(n_478) );
OAI31xp33_ASAP7_75t_L g479 ( .A1(n_443), .A2(n_426), .A3(n_411), .B(n_409), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_456), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_437), .A2(n_434), .B1(n_416), .B2(n_409), .Y(n_481) );
AOI21xp33_ASAP7_75t_L g482 ( .A1(n_438), .A2(n_408), .B(n_436), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_461), .B(n_403), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_465), .B(n_418), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_452), .Y(n_485) );
OR2x6_ASAP7_75t_L g486 ( .A(n_461), .B(n_426), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_456), .B(n_428), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_452), .Y(n_488) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_468), .A2(n_408), .B(n_417), .Y(n_489) );
NOR3xp33_ASAP7_75t_SL g490 ( .A(n_462), .B(n_416), .C(n_417), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g491 ( .A1(n_469), .A2(n_428), .B1(n_415), .B2(n_435), .C(n_436), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_440), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_440), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_457), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_457), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_444), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_458), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_462), .Y(n_498) );
NAND2xp33_ASAP7_75t_L g499 ( .A(n_451), .B(n_432), .Y(n_499) );
BUFx2_ASAP7_75t_L g500 ( .A(n_442), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_459), .A2(n_414), .B1(n_352), .B2(n_403), .Y(n_501) );
AOI33xp33_ASAP7_75t_L g502 ( .A1(n_464), .A2(n_230), .A3(n_214), .B1(n_205), .B2(n_231), .B3(n_233), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_444), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_448), .B(n_414), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_445), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_448), .B(n_414), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_464), .B(n_414), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_445), .Y(n_508) );
INVx3_ASAP7_75t_L g509 ( .A(n_458), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_439), .A2(n_352), .B1(n_272), .B2(n_226), .Y(n_510) );
BUFx3_ASAP7_75t_L g511 ( .A(n_442), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_454), .B(n_10), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_454), .B(n_10), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_470), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_470), .B(n_60), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_455), .B(n_13), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_467), .A2(n_311), .B(n_310), .Y(n_517) );
AOI221xp5_ASAP7_75t_L g518 ( .A1(n_449), .A2(n_234), .B1(n_226), .B2(n_240), .C(n_231), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_458), .B(n_14), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_446), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_451), .B(n_15), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_446), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_446), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_458), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_500), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_476), .B(n_455), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_498), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_478), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_474), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_483), .B(n_472), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_504), .B(n_472), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_478), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_504), .B(n_463), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_476), .B(n_450), .Y(n_534) );
NOR3xp33_ASAP7_75t_SL g535 ( .A(n_479), .B(n_466), .C(n_453), .Y(n_535) );
AND2x2_ASAP7_75t_SL g536 ( .A(n_500), .B(n_450), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_506), .B(n_463), .Y(n_537) );
BUFx2_ASAP7_75t_L g538 ( .A(n_475), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_498), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_478), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_477), .Y(n_541) );
AND2x2_ASAP7_75t_SL g542 ( .A(n_483), .B(n_471), .Y(n_542) );
NAND5xp2_ASAP7_75t_SL g543 ( .A(n_481), .B(n_471), .C(n_459), .D(n_473), .E(n_447), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_485), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_516), .B(n_17), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_484), .B(n_447), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_523), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_523), .Y(n_548) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_482), .A2(n_491), .B(n_501), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_485), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_484), .B(n_447), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_485), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_475), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_520), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_507), .B(n_447), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_480), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_488), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_475), .Y(n_558) );
AOI21xp33_ASAP7_75t_SL g559 ( .A1(n_479), .A2(n_447), .B(n_18), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_522), .Y(n_560) );
NAND4xp25_ASAP7_75t_L g561 ( .A(n_491), .B(n_460), .C(n_357), .D(n_17), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_487), .B(n_19), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_490), .B(n_234), .C(n_226), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_488), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_488), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_494), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_483), .B(n_19), .Y(n_567) );
NAND4xp25_ASAP7_75t_SL g568 ( .A(n_516), .B(n_20), .C(n_23), .D(n_36), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_495), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_483), .B(n_37), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_507), .B(n_240), .Y(n_571) );
INVx2_ASAP7_75t_SL g572 ( .A(n_511), .Y(n_572) );
AOI211x1_ASAP7_75t_L g573 ( .A1(n_487), .A2(n_38), .B(n_40), .C(n_42), .Y(n_573) );
OAI221xp5_ASAP7_75t_L g574 ( .A1(n_482), .A2(n_233), .B1(n_214), .B2(n_205), .C(n_226), .Y(n_574) );
AND2x4_ASAP7_75t_SL g575 ( .A(n_486), .B(n_311), .Y(n_575) );
NAND2xp33_ASAP7_75t_SL g576 ( .A(n_521), .B(n_43), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_495), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_512), .B(n_234), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_514), .Y(n_579) );
OAI21xp5_ASAP7_75t_SL g580 ( .A1(n_559), .A2(n_518), .B(n_519), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_536), .A2(n_486), .B1(n_499), .B2(n_501), .Y(n_581) );
INVx2_ASAP7_75t_SL g582 ( .A(n_539), .Y(n_582) );
OAI221xp5_ASAP7_75t_L g583 ( .A1(n_545), .A2(n_486), .B1(n_518), .B2(n_519), .C(n_510), .Y(n_583) );
NAND4xp25_ASAP7_75t_L g584 ( .A(n_561), .B(n_511), .C(n_512), .D(n_513), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_539), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_543), .A2(n_514), .B1(n_513), .B2(n_524), .C(n_505), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_525), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_529), .Y(n_588) );
AND3x1_ASAP7_75t_L g589 ( .A(n_535), .B(n_509), .C(n_497), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_529), .Y(n_590) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_576), .A2(n_486), .B(n_524), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_527), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_534), .A2(n_486), .B1(n_511), .B2(n_524), .Y(n_593) );
AOI21xp33_ASAP7_75t_L g594 ( .A1(n_542), .A2(n_489), .B(n_497), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_525), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_536), .A2(n_497), .B1(n_509), .B2(n_505), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_547), .Y(n_597) );
AOI21xp5_ASAP7_75t_SL g598 ( .A1(n_568), .A2(n_515), .B(n_503), .Y(n_598) );
NOR3xp33_ASAP7_75t_L g599 ( .A(n_562), .B(n_502), .C(n_509), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_533), .B(n_497), .Y(n_600) );
AOI322xp5_ASAP7_75t_L g601 ( .A1(n_542), .A2(n_496), .A3(n_515), .B1(n_509), .B2(n_508), .C1(n_493), .C2(n_492), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_541), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_577), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_577), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_533), .B(n_496), .Y(n_605) );
XOR2x2_ASAP7_75t_L g606 ( .A(n_526), .B(n_515), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_576), .A2(n_515), .B1(n_489), .B2(n_508), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_567), .A2(n_508), .B(n_493), .Y(n_608) );
AO22x1_ASAP7_75t_L g609 ( .A1(n_567), .A2(n_493), .B1(n_492), .B2(n_489), .Y(n_609) );
NOR2x1p5_ASAP7_75t_L g610 ( .A(n_537), .B(n_489), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_537), .B(n_517), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_531), .B(n_517), .Y(n_612) );
NAND2x1p5_ASAP7_75t_L g613 ( .A(n_570), .B(n_538), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_573), .A2(n_182), .B1(n_234), .B2(n_226), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_560), .B(n_44), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_554), .B(n_46), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_556), .Y(n_617) );
NOR3xp33_ASAP7_75t_SL g618 ( .A(n_543), .B(n_52), .C(n_54), .Y(n_618) );
NAND3xp33_ASAP7_75t_SL g619 ( .A(n_570), .B(n_63), .C(n_65), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_551), .B(n_66), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_566), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_549), .A2(n_310), .B1(n_302), .B2(n_257), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_548), .B(n_76), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_549), .A2(n_257), .B1(n_302), .B2(n_546), .Y(n_624) );
OAI211xp5_ASAP7_75t_SL g625 ( .A1(n_553), .A2(n_558), .B(n_555), .C(n_569), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_555), .A2(n_575), .B1(n_549), .B2(n_538), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_588), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_591), .A2(n_572), .B(n_575), .Y(n_628) );
INVx2_ASAP7_75t_SL g629 ( .A(n_605), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_585), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_617), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_587), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_L g633 ( .A1(n_591), .A2(n_572), .B(n_530), .C(n_579), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_605), .B(n_530), .Y(n_634) );
NOR3xp33_ASAP7_75t_SL g635 ( .A(n_584), .B(n_563), .C(n_578), .Y(n_635) );
CKINVDCx20_ASAP7_75t_L g636 ( .A(n_582), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_597), .B(n_579), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_597), .B(n_530), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_621), .Y(n_639) );
NAND2xp33_ASAP7_75t_R g640 ( .A(n_618), .B(n_528), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_600), .B(n_528), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_590), .Y(n_642) );
INVx1_ASAP7_75t_SL g643 ( .A(n_592), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g644 ( .A(n_616), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_611), .B(n_532), .Y(n_645) );
AOI21xp33_ASAP7_75t_L g646 ( .A1(n_626), .A2(n_571), .B(n_540), .Y(n_646) );
NAND2x1_ASAP7_75t_SL g647 ( .A(n_607), .B(n_532), .Y(n_647) );
XNOR2xp5_ASAP7_75t_L g648 ( .A(n_606), .B(n_571), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_584), .B(n_544), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_583), .A2(n_544), .B1(n_550), .B2(n_552), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_602), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_603), .Y(n_652) );
INVx2_ASAP7_75t_SL g653 ( .A(n_613), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_613), .B(n_550), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_604), .Y(n_655) );
OAI21xp33_ASAP7_75t_SL g656 ( .A1(n_601), .A2(n_552), .B(n_557), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_586), .B(n_557), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_595), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_633), .A2(n_598), .B(n_625), .Y(n_659) );
NAND2xp33_ASAP7_75t_SL g660 ( .A(n_635), .B(n_626), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_649), .B(n_612), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_637), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_656), .B(n_594), .C(n_581), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_631), .Y(n_664) );
NOR3x1_ASAP7_75t_L g665 ( .A(n_657), .B(n_596), .C(n_653), .Y(n_665) );
AOI21xp33_ASAP7_75t_SL g666 ( .A1(n_650), .A2(n_593), .B(n_614), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_635), .A2(n_580), .B(n_619), .Y(n_667) );
NOR2x1_ASAP7_75t_SL g668 ( .A(n_629), .B(n_580), .Y(n_668) );
OAI21x1_ASAP7_75t_L g669 ( .A1(n_647), .A2(n_610), .B(n_589), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_650), .A2(n_608), .B(n_609), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_649), .B(n_624), .Y(n_671) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_632), .Y(n_672) );
NOR2x1_ASAP7_75t_L g673 ( .A(n_643), .B(n_615), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_627), .Y(n_674) );
XNOR2xp5_ASAP7_75t_L g675 ( .A(n_630), .B(n_620), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_646), .B(n_599), .Y(n_676) );
OAI21xp33_ASAP7_75t_L g677 ( .A1(n_638), .A2(n_623), .B(n_622), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_645), .B(n_564), .Y(n_678) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_672), .Y(n_679) );
NOR2xp33_ASAP7_75t_R g680 ( .A(n_660), .B(n_644), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_668), .B(n_634), .Y(n_681) );
AOI21xp33_ASAP7_75t_L g682 ( .A1(n_667), .A2(n_640), .B(n_648), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_664), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_661), .B(n_658), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_672), .B(n_641), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_674), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_660), .A2(n_639), .B1(n_632), .B2(n_655), .C(n_652), .Y(n_687) );
AOI221x1_ASAP7_75t_L g688 ( .A1(n_659), .A2(n_628), .B1(n_636), .B2(n_642), .C(n_651), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_676), .A2(n_640), .B1(n_644), .B2(n_654), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g690 ( .A1(n_676), .A2(n_565), .B(n_574), .C(n_666), .Y(n_690) );
OAI221xp5_ASAP7_75t_L g691 ( .A1(n_663), .A2(n_565), .B1(n_671), .B2(n_670), .C(n_673), .Y(n_691) );
INVxp67_ASAP7_75t_L g692 ( .A(n_675), .Y(n_692) );
XNOR2xp5_ASAP7_75t_L g693 ( .A(n_662), .B(n_678), .Y(n_693) );
NAND4xp25_ASAP7_75t_L g694 ( .A(n_665), .B(n_677), .C(n_674), .D(n_669), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_669), .A2(n_660), .B1(n_676), .B2(n_671), .Y(n_695) );
AOI21xp33_ASAP7_75t_SL g696 ( .A1(n_676), .A2(n_667), .B(n_663), .Y(n_696) );
NAND4xp75_ASAP7_75t_L g697 ( .A(n_688), .B(n_695), .C(n_682), .D(n_689), .Y(n_697) );
BUFx6f_ASAP7_75t_L g698 ( .A(n_681), .Y(n_698) );
NAND4xp25_ASAP7_75t_L g699 ( .A(n_696), .B(n_682), .C(n_694), .D(n_691), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_679), .Y(n_700) );
BUFx4f_ASAP7_75t_L g701 ( .A(n_681), .Y(n_701) );
NAND4xp75_ASAP7_75t_L g702 ( .A(n_697), .B(n_687), .C(n_680), .D(n_684), .Y(n_702) );
XOR2xp5_ASAP7_75t_L g703 ( .A(n_699), .B(n_693), .Y(n_703) );
OR2x6_ASAP7_75t_L g704 ( .A(n_698), .B(n_692), .Y(n_704) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_704), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_703), .B(n_700), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_705), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_706), .Y(n_708) );
AOI322xp5_ASAP7_75t_L g709 ( .A1(n_707), .A2(n_702), .A3(n_698), .B1(n_685), .B2(n_701), .C1(n_686), .C2(n_683), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_709), .A2(n_708), .B(n_690), .Y(n_710) );
endmodule