module fake_netlist_1_7967_n_1356 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1356);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1356;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_298;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g290 ( .A(n_25), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_6), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_109), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_193), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_288), .B(n_69), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_167), .Y(n_295) );
INVxp33_ASAP7_75t_L g296 ( .A(n_243), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_88), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_68), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_41), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_49), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_251), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_225), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_62), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_107), .Y(n_304) );
INVxp67_ASAP7_75t_SL g305 ( .A(n_121), .Y(n_305) );
CKINVDCx16_ASAP7_75t_R g306 ( .A(n_44), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_210), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_142), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_42), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_230), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_33), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_56), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_117), .Y(n_313) );
INVxp67_ASAP7_75t_L g314 ( .A(n_214), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_259), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_240), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_38), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_5), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_247), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g320 ( .A(n_275), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_27), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_285), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_101), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_13), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_131), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_197), .Y(n_326) );
INVxp67_ASAP7_75t_SL g327 ( .A(n_11), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_153), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_192), .Y(n_329) );
INVxp67_ASAP7_75t_L g330 ( .A(n_66), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_94), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_43), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_129), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_208), .Y(n_334) );
INVxp67_ASAP7_75t_L g335 ( .A(n_218), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_204), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_93), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_191), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_143), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_38), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_4), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_11), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_54), .Y(n_343) );
INVxp33_ASAP7_75t_L g344 ( .A(n_65), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_289), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_60), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_227), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_163), .Y(n_348) );
INVxp67_ASAP7_75t_L g349 ( .A(n_154), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_62), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_226), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_166), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_110), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_217), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_31), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_186), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_28), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_73), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_48), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_0), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_125), .Y(n_361) );
INVxp67_ASAP7_75t_L g362 ( .A(n_253), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_222), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_30), .Y(n_364) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_6), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_123), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_59), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_43), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_70), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_231), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_23), .Y(n_371) );
CKINVDCx16_ASAP7_75t_R g372 ( .A(n_281), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_263), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_103), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_60), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_75), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_207), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_178), .Y(n_378) );
INVxp33_ASAP7_75t_SL g379 ( .A(n_250), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_237), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_120), .Y(n_381) );
NOR2xp33_ASAP7_75t_R g382 ( .A(n_257), .B(n_82), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_16), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_245), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_104), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_63), .Y(n_386) );
CKINVDCx16_ASAP7_75t_R g387 ( .A(n_180), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_224), .Y(n_388) );
CKINVDCx16_ASAP7_75t_R g389 ( .A(n_132), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_156), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_4), .Y(n_391) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_238), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_258), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_13), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_61), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_7), .Y(n_396) );
INVxp33_ASAP7_75t_SL g397 ( .A(n_176), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_198), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_213), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_277), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_9), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_99), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_187), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_45), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_170), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_216), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_172), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_146), .Y(n_408) );
CKINVDCx16_ASAP7_75t_R g409 ( .A(n_200), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_232), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_147), .Y(n_411) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_113), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_202), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_236), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_173), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_115), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_32), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_279), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_185), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_44), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_83), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_29), .Y(n_422) );
INVxp33_ASAP7_75t_L g423 ( .A(n_219), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_203), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_215), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_49), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_133), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_76), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_28), .Y(n_429) );
BUFx10_ASAP7_75t_L g430 ( .A(n_21), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_5), .Y(n_431) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_169), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_221), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_375), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_291), .B(n_0), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_296), .B(n_1), .Y(n_436) );
CKINVDCx16_ASAP7_75t_R g437 ( .A(n_372), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_319), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_301), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_300), .B(n_1), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_319), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_301), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_322), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_291), .B(n_2), .Y(n_444) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_301), .Y(n_445) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_322), .A2(n_2), .B(n_3), .Y(n_446) );
NAND2xp33_ASAP7_75t_SL g447 ( .A(n_344), .B(n_3), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_301), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_375), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_396), .B(n_7), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_301), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_323), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_296), .B(n_8), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_375), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_423), .B(n_8), .Y(n_455) );
OR2x6_ASAP7_75t_L g456 ( .A(n_300), .B(n_342), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_308), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_308), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_342), .B(n_9), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_344), .B(n_10), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_413), .B(n_10), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_308), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_323), .Y(n_463) );
AND2x2_ASAP7_75t_SL g464 ( .A(n_326), .B(n_89), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_326), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_308), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_445), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_445), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_456), .B(n_423), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_437), .B(n_314), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_445), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_437), .B(n_387), .Y(n_472) );
INVx5_ASAP7_75t_L g473 ( .A(n_445), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_456), .Y(n_474) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_445), .Y(n_475) );
INVx1_ASAP7_75t_SL g476 ( .A(n_456), .Y(n_476) );
BUFx2_ASAP7_75t_L g477 ( .A(n_456), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_435), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_445), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_456), .B(n_422), .Y(n_480) );
NAND2x1p5_ASAP7_75t_L g481 ( .A(n_464), .B(n_292), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_456), .B(n_422), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_438), .A2(n_429), .B1(n_428), .B2(n_298), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_456), .Y(n_484) );
INVx4_ASAP7_75t_SL g485 ( .A(n_435), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_435), .B(n_396), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_435), .B(n_431), .Y(n_487) );
INVx5_ASAP7_75t_L g488 ( .A(n_445), .Y(n_488) );
INVx5_ASAP7_75t_L g489 ( .A(n_445), .Y(n_489) );
INVx4_ASAP7_75t_L g490 ( .A(n_435), .Y(n_490) );
INVx2_ASAP7_75t_SL g491 ( .A(n_438), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_451), .Y(n_492) );
INVx4_ASAP7_75t_L g493 ( .A(n_435), .Y(n_493) );
BUFx4f_ASAP7_75t_L g494 ( .A(n_464), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_451), .Y(n_495) );
INVx3_ASAP7_75t_L g496 ( .A(n_444), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_438), .B(n_334), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_444), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_444), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_444), .Y(n_500) );
INVx3_ASAP7_75t_L g501 ( .A(n_444), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_441), .B(n_334), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_451), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_444), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_450), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_451), .Y(n_506) );
AND2x6_ASAP7_75t_L g507 ( .A(n_450), .B(n_315), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_441), .B(n_389), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_460), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_450), .B(n_431), .Y(n_510) );
OAI221xp5_ASAP7_75t_L g511 ( .A1(n_447), .A2(n_365), .B1(n_327), .B2(n_429), .C(n_428), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_476), .B(n_464), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_477), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_485), .Y(n_514) );
OR2x6_ASAP7_75t_L g515 ( .A(n_477), .B(n_440), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_485), .Y(n_516) );
INVx3_ASAP7_75t_L g517 ( .A(n_490), .Y(n_517) );
BUFx3_ASAP7_75t_L g518 ( .A(n_507), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_490), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_480), .B(n_450), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_509), .B(n_453), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_484), .B(n_440), .Y(n_522) );
BUFx3_ASAP7_75t_L g523 ( .A(n_507), .Y(n_523) );
INVx5_ASAP7_75t_L g524 ( .A(n_507), .Y(n_524) );
BUFx12f_ASAP7_75t_L g525 ( .A(n_480), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_485), .Y(n_526) );
INVx3_ASAP7_75t_L g527 ( .A(n_490), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_484), .B(n_459), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_485), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_490), .Y(n_530) );
AND2x2_ASAP7_75t_SL g531 ( .A(n_494), .B(n_464), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_480), .B(n_450), .Y(n_532) );
BUFx12f_ASAP7_75t_L g533 ( .A(n_480), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_469), .B(n_453), .Y(n_534) );
BUFx2_ASAP7_75t_L g535 ( .A(n_480), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_485), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_493), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_470), .B(n_461), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_485), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_494), .A2(n_450), .B1(n_447), .B2(n_455), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_493), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_493), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_496), .Y(n_543) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_499), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_494), .A2(n_443), .B(n_452), .C(n_441), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_482), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_496), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_496), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_482), .B(n_459), .Y(n_549) );
INVx5_ASAP7_75t_L g550 ( .A(n_507), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_493), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_496), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_494), .A2(n_446), .B1(n_452), .B2(n_443), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_469), .B(n_455), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_501), .Y(n_555) );
OR2x2_ASAP7_75t_SL g556 ( .A(n_476), .B(n_306), .Y(n_556) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_499), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_501), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_481), .A2(n_443), .B1(n_463), .B2(n_452), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_501), .Y(n_560) );
OAI22xp33_ASAP7_75t_L g561 ( .A1(n_474), .A2(n_460), .B1(n_461), .B2(n_318), .Y(n_561) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_499), .Y(n_562) );
CKINVDCx14_ASAP7_75t_R g563 ( .A(n_482), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_501), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_491), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_491), .B(n_463), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_491), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_478), .Y(n_568) );
AND3x1_ASAP7_75t_SL g569 ( .A(n_511), .B(n_303), .C(n_290), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_478), .Y(n_570) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_507), .Y(n_571) );
INVx3_ASAP7_75t_L g572 ( .A(n_486), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_508), .B(n_379), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_472), .B(n_379), .Y(n_574) );
INVx4_ASAP7_75t_L g575 ( .A(n_482), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_498), .A2(n_465), .B(n_463), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_482), .B(n_465), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_507), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_507), .B(n_465), .Y(n_579) );
INVx5_ASAP7_75t_L g580 ( .A(n_507), .Y(n_580) );
NAND2x1p5_ASAP7_75t_L g581 ( .A(n_498), .B(n_446), .Y(n_581) );
INVx2_ASAP7_75t_SL g582 ( .A(n_507), .Y(n_582) );
BUFx8_ASAP7_75t_L g583 ( .A(n_486), .Y(n_583) );
INVx5_ASAP7_75t_L g584 ( .A(n_486), .Y(n_584) );
INVx4_ASAP7_75t_L g585 ( .A(n_486), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_474), .Y(n_586) );
BUFx4f_ASAP7_75t_L g587 ( .A(n_481), .Y(n_587) );
INVx3_ASAP7_75t_L g588 ( .A(n_486), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_487), .B(n_436), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_500), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_487), .B(n_409), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_483), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_487), .B(n_436), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_481), .A2(n_446), .B1(n_397), .B2(n_320), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_500), .Y(n_595) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_487), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_481), .B(n_430), .Y(n_597) );
O2A1O1Ixp5_ASAP7_75t_L g598 ( .A1(n_534), .A2(n_497), .B(n_502), .C(n_504), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_585), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_522), .B(n_483), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_575), .B(n_487), .Y(n_601) );
INVx6_ASAP7_75t_L g602 ( .A(n_583), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_531), .A2(n_320), .B1(n_378), .B2(n_297), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_517), .Y(n_604) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_571), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_592), .A2(n_511), .B1(n_505), .B2(n_504), .Y(n_606) );
NAND2x1p5_ASAP7_75t_L g607 ( .A(n_575), .B(n_510), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_517), .Y(n_608) );
AND2x4_ASAP7_75t_L g609 ( .A(n_575), .B(n_510), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_583), .Y(n_610) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_571), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_522), .B(n_311), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_585), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_531), .A2(n_505), .B1(n_502), .B2(n_497), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_528), .B(n_311), .Y(n_615) );
INVx3_ASAP7_75t_L g616 ( .A(n_596), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_554), .A2(n_510), .B(n_446), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_538), .B(n_510), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_592), .A2(n_378), .B1(n_388), .B2(n_297), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_597), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_517), .Y(n_621) );
INVx3_ASAP7_75t_L g622 ( .A(n_596), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_549), .B(n_510), .Y(n_623) );
INVx5_ASAP7_75t_L g624 ( .A(n_571), .Y(n_624) );
INVx6_ASAP7_75t_SL g625 ( .A(n_589), .Y(n_625) );
BUFx2_ASAP7_75t_L g626 ( .A(n_583), .Y(n_626) );
INVx3_ASAP7_75t_L g627 ( .A(n_596), .Y(n_627) );
AOI21x1_ASAP7_75t_L g628 ( .A1(n_579), .A2(n_471), .B(n_467), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_519), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_596), .Y(n_630) );
INVx6_ASAP7_75t_L g631 ( .A(n_583), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_566), .A2(n_446), .B(n_294), .Y(n_632) );
AOI21xp5_ASAP7_75t_SL g633 ( .A1(n_518), .A2(n_446), .B(n_392), .Y(n_633) );
OR2x6_ASAP7_75t_L g634 ( .A(n_525), .B(n_309), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_577), .B(n_388), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_585), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_561), .A2(n_332), .B1(n_340), .B2(n_317), .C(n_312), .Y(n_637) );
AND2x6_ASAP7_75t_L g638 ( .A(n_518), .B(n_315), .Y(n_638) );
BUFx2_ASAP7_75t_L g639 ( .A(n_525), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g640 ( .A1(n_531), .A2(n_318), .B1(n_360), .B2(n_341), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_528), .B(n_324), .Y(n_641) );
CKINVDCx5p33_ASAP7_75t_R g642 ( .A(n_533), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_519), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g644 ( .A(n_533), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_519), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_563), .A2(n_369), .B1(n_324), .B2(n_360), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_596), .Y(n_647) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_571), .Y(n_648) );
OR2x6_ASAP7_75t_L g649 ( .A(n_515), .B(n_343), .Y(n_649) );
BUFx3_ASAP7_75t_L g650 ( .A(n_584), .Y(n_650) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_571), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_535), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_544), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_572), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_527), .Y(n_655) );
INVx4_ASAP7_75t_L g656 ( .A(n_524), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_572), .Y(n_657) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_540), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_597), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_549), .B(n_369), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_535), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_515), .Y(n_662) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_523), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_559), .A2(n_341), .B1(n_401), .B2(n_376), .Y(n_664) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_546), .Y(n_665) );
BUFx2_ASAP7_75t_L g666 ( .A(n_515), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_527), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_527), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_530), .Y(n_669) );
BUFx2_ASAP7_75t_SL g670 ( .A(n_524), .Y(n_670) );
BUFx3_ASAP7_75t_L g671 ( .A(n_584), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_572), .Y(n_672) );
AND2x4_ASAP7_75t_L g673 ( .A(n_577), .B(n_346), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_588), .Y(n_674) );
INVx2_ASAP7_75t_SL g675 ( .A(n_589), .Y(n_675) );
BUFx8_ASAP7_75t_SL g676 ( .A(n_515), .Y(n_676) );
BUFx2_ASAP7_75t_L g677 ( .A(n_515), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_540), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_588), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_588), .A2(n_397), .B1(n_355), .B2(n_357), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_530), .Y(n_681) );
INVx2_ASAP7_75t_SL g682 ( .A(n_589), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_513), .B(n_376), .Y(n_683) );
INVx1_ASAP7_75t_SL g684 ( .A(n_513), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_512), .A2(n_401), .B1(n_321), .B2(n_359), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_576), .A2(n_412), .B(n_305), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_559), .B(n_350), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_543), .A2(n_432), .B(n_295), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_584), .Y(n_689) );
AND2x4_ASAP7_75t_L g690 ( .A(n_589), .B(n_358), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_584), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_530), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_584), .Y(n_693) );
AO22x1_ASAP7_75t_L g694 ( .A1(n_520), .A2(n_325), .B1(n_351), .B2(n_304), .Y(n_694) );
BUFx3_ASAP7_75t_L g695 ( .A(n_584), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_537), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_520), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_543), .A2(n_302), .B(n_293), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_586), .A2(n_299), .B1(n_330), .B2(n_325), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_520), .Y(n_700) );
BUFx6f_ASAP7_75t_L g701 ( .A(n_523), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_520), .B(n_364), .Y(n_702) );
BUFx6f_ASAP7_75t_L g703 ( .A(n_524), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_532), .Y(n_704) );
BUFx12f_ASAP7_75t_L g705 ( .A(n_556), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_556), .B(n_367), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_547), .A2(n_310), .B(n_307), .Y(n_707) );
AND2x6_ASAP7_75t_L g708 ( .A(n_532), .B(n_514), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_532), .A2(n_371), .B1(n_383), .B2(n_368), .Y(n_709) );
BUFx8_ASAP7_75t_L g710 ( .A(n_532), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_521), .B(n_386), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_568), .B(n_391), .Y(n_712) );
AND2x4_ASAP7_75t_L g713 ( .A(n_524), .B(n_394), .Y(n_713) );
NOR2xp33_ASAP7_75t_SL g714 ( .A(n_587), .B(n_304), .Y(n_714) );
BUFx12f_ASAP7_75t_L g715 ( .A(n_524), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_568), .B(n_395), .Y(n_716) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_524), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_593), .Y(n_718) );
NOR2xp33_ASAP7_75t_SL g719 ( .A(n_587), .B(n_351), .Y(n_719) );
INVxp67_ASAP7_75t_L g720 ( .A(n_586), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_635), .B(n_574), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_607), .Y(n_722) );
BUFx12f_ASAP7_75t_L g723 ( .A(n_642), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_607), .Y(n_724) );
AND2x4_ASAP7_75t_L g725 ( .A(n_649), .B(n_550), .Y(n_725) );
O2A1O1Ixp5_ASAP7_75t_L g726 ( .A1(n_598), .A2(n_545), .B(n_587), .C(n_591), .Y(n_726) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_619), .A2(n_594), .B1(n_550), .B2(n_580), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_612), .B(n_573), .Y(n_728) );
OAI22xp33_ASAP7_75t_SL g729 ( .A1(n_649), .A2(n_594), .B1(n_417), .B2(n_420), .Y(n_729) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_605), .Y(n_730) );
NAND2x1p5_ASAP7_75t_L g731 ( .A(n_626), .B(n_550), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_702), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_615), .A2(n_600), .B1(n_640), .B2(n_658), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_640), .A2(n_542), .B1(n_537), .B2(n_541), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_702), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_678), .A2(n_542), .B1(n_537), .B2(n_541), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g737 ( .A(n_676), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_664), .B(n_570), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_601), .Y(n_739) );
INVx4_ASAP7_75t_SL g740 ( .A(n_602), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_712), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_683), .A2(n_542), .B1(n_551), .B2(n_570), .Y(n_742) );
OR2x2_ASAP7_75t_L g743 ( .A(n_664), .B(n_590), .Y(n_743) );
BUFx2_ASAP7_75t_L g744 ( .A(n_649), .Y(n_744) );
OAI21x1_ASAP7_75t_L g745 ( .A1(n_628), .A2(n_581), .B(n_590), .Y(n_745) );
AO32x2_ASAP7_75t_L g746 ( .A1(n_614), .A2(n_582), .A3(n_578), .B1(n_553), .B2(n_569), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_601), .Y(n_747) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_605), .Y(n_748) );
INVx6_ASAP7_75t_L g749 ( .A(n_710), .Y(n_749) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_644), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_641), .B(n_430), .Y(n_751) );
AND2x4_ASAP7_75t_L g752 ( .A(n_610), .B(n_550), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_712), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g754 ( .A(n_634), .Y(n_754) );
BUFx3_ASAP7_75t_L g755 ( .A(n_602), .Y(n_755) );
CKINVDCx12_ASAP7_75t_R g756 ( .A(n_634), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_716), .Y(n_757) );
INVx5_ASAP7_75t_L g758 ( .A(n_602), .Y(n_758) );
INVx2_ASAP7_75t_SL g759 ( .A(n_631), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_716), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_635), .A2(n_551), .B1(n_595), .B2(n_557), .Y(n_761) );
NOR2x1_ASAP7_75t_SL g762 ( .A(n_634), .B(n_550), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_614), .A2(n_595), .B1(n_581), .B2(n_550), .Y(n_763) );
BUFx6f_ASAP7_75t_L g764 ( .A(n_605), .Y(n_764) );
A2O1A1Ixp33_ASAP7_75t_L g765 ( .A1(n_598), .A2(n_548), .B(n_555), .C(n_547), .Y(n_765) );
INVx3_ASAP7_75t_L g766 ( .A(n_631), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_662), .A2(n_666), .B1(n_677), .B2(n_687), .Y(n_767) );
OAI22xp33_ASAP7_75t_L g768 ( .A1(n_619), .A2(n_580), .B1(n_582), .B2(n_578), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_609), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_625), .A2(n_557), .B1(n_562), .B2(n_544), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_625), .A2(n_652), .B1(n_661), .B2(n_609), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_652), .A2(n_557), .B1(n_562), .B2(n_544), .Y(n_772) );
NAND2xp33_ASAP7_75t_L g773 ( .A(n_638), .B(n_580), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g774 ( .A(n_705), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_687), .A2(n_581), .B1(n_580), .B2(n_557), .Y(n_775) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_631), .A2(n_430), .B1(n_580), .B2(n_382), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_603), .A2(n_548), .B1(n_560), .B2(n_555), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_684), .B(n_404), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_618), .B(n_560), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_673), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_661), .A2(n_557), .B1(n_562), .B2(n_544), .Y(n_781) );
OR2x2_ASAP7_75t_L g782 ( .A(n_646), .B(n_544), .Y(n_782) );
BUFx6f_ASAP7_75t_L g783 ( .A(n_605), .Y(n_783) );
OAI22xp33_ASAP7_75t_L g784 ( .A1(n_714), .A2(n_580), .B1(n_562), .B2(n_558), .Y(n_784) );
A2O1A1Ixp33_ASAP7_75t_L g785 ( .A1(n_618), .A2(n_564), .B(n_558), .C(n_552), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_620), .B(n_562), .Y(n_786) );
OAI21xp5_ASAP7_75t_L g787 ( .A1(n_617), .A2(n_564), .B(n_552), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_659), .A2(n_526), .B1(n_529), .B2(n_514), .Y(n_788) );
OR2x2_ASAP7_75t_L g789 ( .A(n_660), .B(n_421), .Y(n_789) );
A2O1A1Ixp33_ASAP7_75t_L g790 ( .A1(n_711), .A2(n_526), .B(n_536), .C(n_529), .Y(n_790) );
INVx4_ASAP7_75t_SL g791 ( .A(n_638), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_660), .B(n_426), .Y(n_792) );
AND2x4_ASAP7_75t_L g793 ( .A(n_610), .B(n_536), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_637), .A2(n_539), .B1(n_516), .B2(n_565), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g795 ( .A1(n_606), .A2(n_375), .B1(n_316), .B2(n_329), .C(n_328), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_673), .Y(n_796) );
INVx6_ASAP7_75t_L g797 ( .A(n_710), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_623), .A2(n_565), .B1(n_375), .B2(n_313), .Y(n_798) );
OAI22xp33_ASAP7_75t_L g799 ( .A1(n_719), .A2(n_720), .B1(n_685), .B2(n_699), .Y(n_799) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_639), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_623), .A2(n_331), .B1(n_336), .B2(n_333), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_720), .A2(n_539), .B1(n_516), .B2(n_380), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_606), .A2(n_380), .B1(n_399), .B2(n_354), .Y(n_803) );
CKINVDCx6p67_ASAP7_75t_R g804 ( .A(n_715), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_604), .Y(n_805) );
CKINVDCx11_ASAP7_75t_R g806 ( .A(n_690), .Y(n_806) );
OR2x2_ASAP7_75t_L g807 ( .A(n_706), .B(n_694), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_690), .Y(n_808) );
AND2x4_ASAP7_75t_L g809 ( .A(n_697), .B(n_567), .Y(n_809) );
BUFx3_ASAP7_75t_L g810 ( .A(n_650), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_637), .A2(n_399), .B1(n_400), .B2(n_354), .Y(n_811) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_713), .Y(n_812) );
AOI221xp5_ASAP7_75t_L g813 ( .A1(n_711), .A2(n_408), .B1(n_381), .B2(n_337), .C(n_384), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_675), .A2(n_348), .B1(n_353), .B2(n_339), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_682), .A2(n_361), .B1(n_363), .B2(n_356), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_665), .A2(n_370), .B1(n_377), .B2(n_366), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_599), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_700), .A2(n_390), .B1(n_393), .B2(n_385), .Y(n_818) );
INVx3_ASAP7_75t_L g819 ( .A(n_671), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_665), .A2(n_402), .B1(n_405), .B2(n_398), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_608), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_718), .A2(n_411), .B1(n_425), .B2(n_400), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_680), .B(n_411), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_621), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_704), .A2(n_407), .B1(n_410), .B2(n_406), .Y(n_825) );
INVx3_ASAP7_75t_L g826 ( .A(n_695), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_613), .A2(n_416), .B1(n_418), .B2(n_414), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_617), .B(n_567), .Y(n_828) );
AOI221xp5_ASAP7_75t_L g829 ( .A1(n_709), .A2(n_424), .B1(n_427), .B2(n_433), .C(n_403), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_709), .A2(n_698), .B1(n_707), .B2(n_632), .Y(n_830) );
OAI22xp33_ASAP7_75t_L g831 ( .A1(n_654), .A2(n_425), .B1(n_335), .B2(n_349), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_636), .A2(n_352), .B1(n_373), .B2(n_347), .Y(n_832) );
NAND2x1p5_ASAP7_75t_L g833 ( .A(n_624), .B(n_345), .Y(n_833) );
O2A1O1Ixp33_ASAP7_75t_SL g834 ( .A1(n_632), .A2(n_362), .B(n_374), .C(n_338), .Y(n_834) );
OR2x2_ASAP7_75t_L g835 ( .A(n_680), .B(n_12), .Y(n_835) );
AOI221xp5_ASAP7_75t_L g836 ( .A1(n_688), .A2(n_686), .B1(n_698), .B2(n_707), .C(n_674), .Y(n_836) );
OAI21x1_ASAP7_75t_L g837 ( .A1(n_633), .A2(n_352), .B(n_347), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_657), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_672), .B(n_373), .Y(n_839) );
AOI22xp5_ASAP7_75t_L g840 ( .A1(n_708), .A2(n_419), .B1(n_415), .B2(n_308), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_629), .Y(n_841) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_713), .Y(n_842) );
OR2x6_ASAP7_75t_L g843 ( .A(n_670), .B(n_419), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_708), .A2(n_415), .B1(n_449), .B2(n_434), .Y(n_844) );
NOR2xp67_ASAP7_75t_SL g845 ( .A(n_624), .B(n_415), .Y(n_845) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_616), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_679), .Y(n_847) );
OA21x2_ASAP7_75t_L g848 ( .A1(n_688), .A2(n_471), .B(n_467), .Y(n_848) );
OAI221xp5_ASAP7_75t_L g849 ( .A1(n_686), .A2(n_454), .B1(n_434), .B2(n_449), .C(n_442), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_643), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_645), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_624), .A2(n_442), .B1(n_448), .B2(n_439), .Y(n_852) );
BUFx8_ASAP7_75t_L g853 ( .A(n_689), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_691), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_733), .B(n_693), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_728), .B(n_616), .Y(n_856) );
OR2x2_ASAP7_75t_L g857 ( .A(n_808), .B(n_738), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_741), .A2(n_638), .B1(n_708), .B2(n_627), .Y(n_858) );
BUFx6f_ASAP7_75t_L g859 ( .A(n_730), .Y(n_859) );
AOI21xp5_ASAP7_75t_L g860 ( .A1(n_828), .A2(n_653), .B(n_651), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_751), .B(n_622), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_743), .B(n_622), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_753), .B(n_627), .Y(n_863) );
NOR2x1_ASAP7_75t_R g864 ( .A(n_749), .B(n_624), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_780), .Y(n_865) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_722), .Y(n_866) );
INVx8_ASAP7_75t_L g867 ( .A(n_758), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_757), .A2(n_638), .B1(n_708), .B2(n_647), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_760), .A2(n_638), .B1(n_708), .B2(n_647), .Y(n_869) );
OAI21x1_ASAP7_75t_L g870 ( .A1(n_828), .A2(n_653), .B(n_630), .Y(n_870) );
INVx3_ASAP7_75t_L g871 ( .A(n_725), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_796), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_778), .B(n_630), .Y(n_873) );
OAI21xp5_ASAP7_75t_SL g874 ( .A1(n_734), .A2(n_701), .B(n_663), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_835), .A2(n_667), .B1(n_668), .B2(n_655), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_792), .B(n_669), .Y(n_876) );
BUFx12f_ASAP7_75t_L g877 ( .A(n_723), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_817), .Y(n_878) );
AND2x4_ASAP7_75t_L g879 ( .A(n_740), .B(n_656), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_721), .A2(n_692), .B1(n_696), .B2(n_681), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_727), .A2(n_663), .B1(n_701), .B2(n_656), .Y(n_881) );
OAI22xp33_ASAP7_75t_L g882 ( .A1(n_843), .A2(n_744), .B1(n_807), .B2(n_763), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_839), .Y(n_883) );
BUFx8_ASAP7_75t_L g884 ( .A(n_756), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_838), .Y(n_885) );
AOI21xp33_ASAP7_75t_L g886 ( .A1(n_799), .A2(n_701), .B(n_663), .Y(n_886) );
OAI211xp5_ASAP7_75t_L g887 ( .A1(n_795), .A2(n_442), .B(n_448), .C(n_439), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_729), .A2(n_701), .B1(n_663), .B2(n_611), .Y(n_888) );
A2O1A1Ixp33_ASAP7_75t_L g889 ( .A1(n_726), .A2(n_651), .B(n_611), .C(n_703), .Y(n_889) );
AOI222xp33_ASAP7_75t_L g890 ( .A1(n_806), .A2(n_454), .B1(n_434), .B2(n_449), .C1(n_415), .C2(n_448), .Y(n_890) );
BUFx6f_ASAP7_75t_L g891 ( .A(n_730), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_749), .A2(n_611), .B1(n_651), .B2(n_703), .Y(n_892) );
INVx3_ASAP7_75t_L g893 ( .A(n_725), .Y(n_893) );
OAI221xp5_ASAP7_75t_L g894 ( .A1(n_742), .A2(n_454), .B1(n_449), .B2(n_434), .C(n_611), .Y(n_894) );
OAI33xp33_ASAP7_75t_L g895 ( .A1(n_801), .A2(n_439), .A3(n_442), .B1(n_448), .B2(n_458), .B3(n_462), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_823), .B(n_12), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_749), .A2(n_651), .B1(n_717), .B2(n_703), .Y(n_897) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_843), .A2(n_648), .B1(n_717), .B2(n_703), .Y(n_898) );
BUFx3_ASAP7_75t_L g899 ( .A(n_804), .Y(n_899) );
OAI22xp33_ASAP7_75t_L g900 ( .A1(n_843), .A2(n_648), .B1(n_717), .B2(n_415), .Y(n_900) );
AO21x2_ASAP7_75t_L g901 ( .A1(n_787), .A2(n_458), .B(n_439), .Y(n_901) );
OAI211xp5_ASAP7_75t_SL g902 ( .A1(n_813), .A2(n_449), .B(n_454), .C(n_434), .Y(n_902) );
AO31x2_ASAP7_75t_L g903 ( .A1(n_830), .A2(n_462), .A3(n_466), .B(n_458), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_763), .A2(n_648), .B1(n_717), .B2(n_462), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_795), .A2(n_454), .B1(n_462), .B2(n_458), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_839), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_813), .B(n_14), .Y(n_907) );
INVxp67_ASAP7_75t_L g908 ( .A(n_754), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_847), .Y(n_909) );
AOI221xp5_ASAP7_75t_L g910 ( .A1(n_801), .A2(n_466), .B1(n_451), .B2(n_457), .C(n_492), .Y(n_910) );
AOI21xp33_ASAP7_75t_L g911 ( .A1(n_830), .A2(n_466), .B(n_14), .Y(n_911) );
AOI22xp33_ASAP7_75t_SL g912 ( .A1(n_797), .A2(n_767), .B1(n_762), .B2(n_816), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_767), .A2(n_466), .B1(n_457), .B2(n_451), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_737), .Y(n_914) );
OR2x2_ASAP7_75t_L g915 ( .A(n_800), .B(n_15), .Y(n_915) );
OAI21xp33_ASAP7_75t_L g916 ( .A1(n_811), .A2(n_457), .B(n_451), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_854), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_822), .B(n_15), .Y(n_918) );
HB1xp67_ASAP7_75t_L g919 ( .A(n_724), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_836), .A2(n_451), .B1(n_457), .B2(n_495), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_789), .Y(n_921) );
OAI211xp5_ASAP7_75t_SL g922 ( .A1(n_829), .A2(n_503), .B(n_495), .C(n_492), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_829), .A2(n_457), .B1(n_503), .B2(n_495), .C(n_492), .Y(n_923) );
AOI21xp5_ASAP7_75t_L g924 ( .A1(n_787), .A2(n_506), .B(n_471), .Y(n_924) );
NAND3xp33_ASAP7_75t_L g925 ( .A(n_776), .B(n_457), .C(n_468), .Y(n_925) );
OAI22xp5_ASAP7_75t_SL g926 ( .A1(n_797), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_732), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_836), .A2(n_457), .B1(n_503), .B2(n_479), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_761), .A2(n_457), .B1(n_18), .B2(n_19), .Y(n_929) );
CKINVDCx20_ASAP7_75t_R g930 ( .A(n_750), .Y(n_930) );
OAI22xp33_ASAP7_75t_L g931 ( .A1(n_803), .A2(n_17), .B1(n_19), .B2(n_20), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_735), .Y(n_932) );
INVx2_ASAP7_75t_SL g933 ( .A(n_797), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_779), .A2(n_506), .B1(n_479), .B2(n_467), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_779), .A2(n_506), .B1(n_479), .B2(n_475), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_768), .A2(n_468), .B1(n_475), .B2(n_22), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_848), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_782), .A2(n_475), .B1(n_468), .B2(n_473), .Y(n_938) );
AOI221xp5_ASAP7_75t_L g939 ( .A1(n_816), .A2(n_475), .B1(n_468), .B2(n_489), .C(n_473), .Y(n_939) );
OAI22xp33_ASAP7_75t_L g940 ( .A1(n_820), .A2(n_20), .B1(n_21), .B2(n_22), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_820), .A2(n_468), .B1(n_475), .B2(n_25), .Y(n_941) );
INVx2_ASAP7_75t_L g942 ( .A(n_848), .Y(n_942) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_739), .B(n_23), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_771), .A2(n_475), .B1(n_468), .B2(n_489), .Y(n_944) );
OAI221xp5_ASAP7_75t_L g945 ( .A1(n_814), .A2(n_475), .B1(n_468), .B2(n_489), .C(n_473), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_805), .Y(n_946) );
INVx2_ASAP7_75t_L g947 ( .A(n_821), .Y(n_947) );
OAI221xp5_ASAP7_75t_L g948 ( .A1(n_815), .A2(n_818), .B1(n_825), .B2(n_827), .C(n_777), .Y(n_948) );
OR2x2_ASAP7_75t_L g949 ( .A(n_747), .B(n_24), .Y(n_949) );
INVx2_ASAP7_75t_L g950 ( .A(n_824), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_841), .Y(n_951) );
BUFx6f_ASAP7_75t_L g952 ( .A(n_730), .Y(n_952) );
OAI22xp33_ASAP7_75t_L g953 ( .A1(n_833), .A2(n_24), .B1(n_26), .B2(n_27), .Y(n_953) );
OAI21x1_ASAP7_75t_L g954 ( .A1(n_745), .A2(n_91), .B(n_90), .Y(n_954) );
OAI211xp5_ASAP7_75t_L g955 ( .A1(n_832), .A2(n_489), .B(n_488), .C(n_473), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_798), .A2(n_26), .B1(n_29), .B2(n_30), .Y(n_956) );
INVxp67_ASAP7_75t_L g957 ( .A(n_853), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_850), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_769), .B(n_31), .Y(n_959) );
INVx4_ASAP7_75t_L g960 ( .A(n_740), .Y(n_960) );
AOI332xp33_ASAP7_75t_L g961 ( .A1(n_794), .A2(n_32), .A3(n_33), .B1(n_34), .B2(n_35), .B3(n_36), .C1(n_37), .C2(n_39), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_849), .A2(n_34), .B1(n_35), .B2(n_36), .Y(n_962) );
HB1xp67_ASAP7_75t_L g963 ( .A(n_786), .Y(n_963) );
OAI221xp5_ASAP7_75t_L g964 ( .A1(n_736), .A2(n_489), .B1(n_488), .B2(n_473), .C(n_41), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_849), .A2(n_37), .B1(n_39), .B2(n_40), .Y(n_965) );
NAND2xp33_ASAP7_75t_R g966 ( .A(n_774), .B(n_40), .Y(n_966) );
OAI22xp33_ASAP7_75t_L g967 ( .A1(n_833), .A2(n_42), .B1(n_45), .B2(n_46), .Y(n_967) );
AOI22xp33_ASAP7_75t_SL g968 ( .A1(n_758), .A2(n_46), .B1(n_47), .B2(n_48), .Y(n_968) );
AO21x2_ASAP7_75t_L g969 ( .A1(n_837), .A2(n_95), .B(n_92), .Y(n_969) );
AOI21x1_ASAP7_75t_L g970 ( .A1(n_775), .A2(n_97), .B(n_96), .Y(n_970) );
CKINVDCx5p33_ASAP7_75t_R g971 ( .A(n_853), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_755), .A2(n_488), .B1(n_473), .B2(n_489), .Y(n_972) );
AOI211xp5_ASAP7_75t_L g973 ( .A1(n_831), .A2(n_47), .B(n_50), .C(n_51), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_798), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_759), .B(n_52), .Y(n_975) );
AOI22xp5_ASAP7_75t_L g976 ( .A1(n_766), .A2(n_489), .B1(n_488), .B2(n_473), .Y(n_976) );
OAI21xp5_ASAP7_75t_L g977 ( .A1(n_785), .A2(n_488), .B(n_53), .Y(n_977) );
OAI22xp33_ASAP7_75t_L g978 ( .A1(n_758), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_909), .Y(n_979) );
OR2x2_ASAP7_75t_L g980 ( .A(n_857), .B(n_810), .Y(n_980) );
INVxp67_ASAP7_75t_SL g981 ( .A(n_900), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g982 ( .A1(n_912), .A2(n_812), .B1(n_842), .B2(n_758), .Y(n_982) );
AOI22xp5_ASAP7_75t_L g983 ( .A1(n_948), .A2(n_766), .B1(n_793), .B2(n_740), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_882), .A2(n_775), .B1(n_840), .B2(n_802), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_937), .Y(n_985) );
INVx2_ASAP7_75t_L g986 ( .A(n_942), .Y(n_986) );
AO21x2_ASAP7_75t_L g987 ( .A1(n_911), .A2(n_834), .B(n_765), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_903), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_885), .Y(n_989) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_866), .Y(n_990) );
OAI31xp33_ASAP7_75t_L g991 ( .A1(n_940), .A2(n_790), .A3(n_731), .B(n_784), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_917), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g993 ( .A1(n_882), .A2(n_793), .B1(n_752), .B2(n_809), .Y(n_993) );
AOI221xp5_ASAP7_75t_L g994 ( .A1(n_921), .A2(n_852), .B1(n_788), .B2(n_844), .C(n_809), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_855), .A2(n_819), .B1(n_826), .B2(n_851), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_931), .A2(n_819), .B1(n_826), .B2(n_846), .Y(n_996) );
NAND5xp2_ASAP7_75t_SL g997 ( .A(n_971), .B(n_55), .C(n_56), .D(n_57), .E(n_58), .Y(n_997) );
INVx2_ASAP7_75t_L g998 ( .A(n_903), .Y(n_998) );
OA21x2_ASAP7_75t_L g999 ( .A1(n_870), .A2(n_781), .B(n_772), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_866), .B(n_746), .Y(n_1000) );
OR2x2_ASAP7_75t_SL g1001 ( .A(n_915), .B(n_57), .Y(n_1001) );
OAI33xp33_ASAP7_75t_L g1002 ( .A1(n_940), .A2(n_852), .A3(n_59), .B1(n_61), .B2(n_63), .B3(n_64), .Y(n_1002) );
AOI221xp5_ASAP7_75t_L g1003 ( .A1(n_931), .A2(n_752), .B1(n_770), .B2(n_731), .C(n_845), .Y(n_1003) );
INVxp67_ASAP7_75t_L g1004 ( .A(n_884), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_878), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_907), .B(n_896), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_919), .B(n_746), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1008 ( .A1(n_941), .A2(n_900), .B1(n_973), .B2(n_936), .Y(n_1008) );
OAI33xp33_ASAP7_75t_L g1009 ( .A1(n_978), .A2(n_58), .A3(n_64), .B1(n_65), .B2(n_66), .B3(n_67), .Y(n_1009) );
AOI33xp33_ASAP7_75t_L g1010 ( .A1(n_962), .A2(n_67), .A3(n_68), .B1(n_69), .B2(n_70), .B3(n_71), .Y(n_1010) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_949), .B(n_71), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_873), .B(n_72), .Y(n_1012) );
AOI221xp5_ASAP7_75t_L g1013 ( .A1(n_953), .A2(n_746), .B1(n_773), .B2(n_764), .C(n_748), .Y(n_1013) );
OAI211xp5_ASAP7_75t_L g1014 ( .A1(n_961), .A2(n_488), .B(n_783), .C(n_764), .Y(n_1014) );
AOI211xp5_ASAP7_75t_L g1015 ( .A1(n_926), .A2(n_748), .B(n_764), .C(n_783), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g1016 ( .A(n_919), .Y(n_1016) );
INVx3_ASAP7_75t_L g1017 ( .A(n_867), .Y(n_1017) );
NOR3xp33_ASAP7_75t_SL g1018 ( .A(n_966), .B(n_791), .C(n_73), .Y(n_1018) );
INVx2_ASAP7_75t_L g1019 ( .A(n_903), .Y(n_1019) );
OAI31xp33_ASAP7_75t_SL g1020 ( .A1(n_953), .A2(n_791), .A3(n_74), .B(n_75), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_865), .Y(n_1021) );
NAND3xp33_ASAP7_75t_L g1022 ( .A(n_890), .B(n_748), .C(n_783), .Y(n_1022) );
OAI221xp5_ASAP7_75t_L g1023 ( .A1(n_962), .A2(n_791), .B1(n_488), .B2(n_76), .C(n_77), .Y(n_1023) );
INVx2_ASAP7_75t_L g1024 ( .A(n_903), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_918), .A2(n_72), .B1(n_74), .B2(n_77), .Y(n_1025) );
NOR2xp33_ASAP7_75t_L g1026 ( .A(n_856), .B(n_78), .Y(n_1026) );
NAND4xp25_ASAP7_75t_L g1027 ( .A(n_965), .B(n_78), .C(n_79), .D(n_80), .Y(n_1027) );
AOI221xp5_ASAP7_75t_L g1028 ( .A1(n_967), .A2(n_79), .B1(n_80), .B2(n_81), .C(n_82), .Y(n_1028) );
INVxp67_ASAP7_75t_SL g1029 ( .A(n_963), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_947), .B(n_81), .Y(n_1030) );
BUFx12f_ASAP7_75t_L g1031 ( .A(n_884), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_872), .Y(n_1032) );
OAI22xp5_ASAP7_75t_SL g1033 ( .A1(n_957), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_950), .B(n_951), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_927), .B(n_84), .Y(n_1035) );
OAI21xp5_ASAP7_75t_L g1036 ( .A1(n_977), .A2(n_85), .B(n_86), .Y(n_1036) );
OAI221xp5_ASAP7_75t_L g1037 ( .A1(n_965), .A2(n_86), .B1(n_87), .B2(n_98), .C(n_100), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_932), .Y(n_1038) );
OAI221xp5_ASAP7_75t_SL g1039 ( .A1(n_974), .A2(n_978), .B1(n_967), .B2(n_941), .C(n_936), .Y(n_1039) );
OA21x2_ASAP7_75t_L g1040 ( .A1(n_889), .A2(n_189), .B(n_102), .Y(n_1040) );
NAND3xp33_ASAP7_75t_L g1041 ( .A(n_968), .B(n_87), .C(n_105), .Y(n_1041) );
AOI33xp33_ASAP7_75t_L g1042 ( .A1(n_974), .A2(n_106), .A3(n_108), .B1(n_111), .B2(n_112), .B3(n_114), .Y(n_1042) );
OAI21xp5_ASAP7_75t_L g1043 ( .A1(n_964), .A2(n_116), .B(n_118), .Y(n_1043) );
AOI222xp33_ASAP7_75t_L g1044 ( .A1(n_956), .A2(n_119), .B1(n_122), .B2(n_124), .C1(n_126), .C2(n_127), .Y(n_1044) );
OAI221xp5_ASAP7_75t_L g1045 ( .A1(n_880), .A2(n_128), .B1(n_130), .B2(n_134), .C(n_135), .Y(n_1045) );
HB1xp67_ASAP7_75t_L g1046 ( .A(n_963), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1047 ( .A1(n_875), .A2(n_136), .B1(n_137), .B2(n_138), .Y(n_1047) );
NAND3xp33_ASAP7_75t_L g1048 ( .A(n_943), .B(n_139), .C(n_140), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_875), .A2(n_141), .B1(n_144), .B2(n_145), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_883), .A2(n_148), .B1(n_149), .B2(n_150), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_946), .B(n_151), .Y(n_1051) );
AND2x2_ASAP7_75t_SL g1052 ( .A(n_960), .B(n_152), .Y(n_1052) );
AO21x2_ASAP7_75t_L g1053 ( .A1(n_901), .A2(n_155), .B(n_157), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_958), .Y(n_1054) );
OAI31xp33_ASAP7_75t_SL g1055 ( .A1(n_898), .A2(n_913), .A3(n_929), .B(n_902), .Y(n_1055) );
INVx2_ASAP7_75t_SL g1056 ( .A(n_867), .Y(n_1056) );
OAI211xp5_ASAP7_75t_L g1057 ( .A1(n_975), .A2(n_158), .B(n_159), .C(n_160), .Y(n_1057) );
OAI211xp5_ASAP7_75t_SL g1058 ( .A1(n_908), .A2(n_161), .B(n_162), .C(n_164), .Y(n_1058) );
INVx2_ASAP7_75t_L g1059 ( .A(n_901), .Y(n_1059) );
BUFx2_ASAP7_75t_L g1060 ( .A(n_867), .Y(n_1060) );
AOI221xp5_ASAP7_75t_L g1061 ( .A1(n_876), .A2(n_165), .B1(n_168), .B2(n_171), .C(n_174), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_906), .A2(n_175), .B1(n_177), .B2(n_179), .Y(n_1062) );
AOI22xp33_ASAP7_75t_SL g1063 ( .A1(n_960), .A2(n_181), .B1(n_182), .B2(n_183), .Y(n_1063) );
OAI31xp33_ASAP7_75t_SL g1064 ( .A1(n_879), .A2(n_184), .A3(n_188), .B(n_190), .Y(n_1064) );
OAI21xp5_ASAP7_75t_L g1065 ( .A1(n_916), .A2(n_194), .B(n_195), .Y(n_1065) );
AOI22xp5_ASAP7_75t_L g1066 ( .A1(n_861), .A2(n_196), .B1(n_199), .B2(n_201), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_959), .B(n_871), .Y(n_1067) );
OR2x2_ASAP7_75t_L g1068 ( .A(n_871), .B(n_287), .Y(n_1068) );
INVx3_ASAP7_75t_L g1069 ( .A(n_879), .Y(n_1069) );
OAI21xp5_ASAP7_75t_L g1070 ( .A1(n_905), .A2(n_205), .B(n_206), .Y(n_1070) );
INVx2_ASAP7_75t_SL g1071 ( .A(n_893), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_895), .A2(n_209), .B1(n_211), .B2(n_212), .Y(n_1072) );
NAND3xp33_ASAP7_75t_L g1073 ( .A(n_920), .B(n_220), .C(n_223), .Y(n_1073) );
OAI21xp5_ASAP7_75t_L g1074 ( .A1(n_905), .A2(n_228), .B(n_229), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_863), .A2(n_233), .B1(n_234), .B2(n_235), .Y(n_1075) );
HB1xp67_ASAP7_75t_L g1076 ( .A(n_893), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_933), .B(n_239), .Y(n_1077) );
NOR2x1_ASAP7_75t_SL g1078 ( .A(n_864), .B(n_241), .Y(n_1078) );
AOI221xp5_ASAP7_75t_L g1079 ( .A1(n_920), .A2(n_242), .B1(n_244), .B2(n_246), .C(n_248), .Y(n_1079) );
AOI33xp33_ASAP7_75t_L g1080 ( .A1(n_928), .A2(n_249), .A3(n_252), .B1(n_254), .B2(n_255), .B3(n_256), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_862), .B(n_260), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_979), .Y(n_1082) );
INVx2_ASAP7_75t_L g1083 ( .A(n_985), .Y(n_1083) );
INVx2_ASAP7_75t_L g1084 ( .A(n_985), .Y(n_1084) );
OAI33xp33_ASAP7_75t_L g1085 ( .A1(n_1033), .A2(n_922), .A3(n_904), .B1(n_925), .B2(n_887), .B3(n_899), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_992), .Y(n_1086) );
INVxp67_ASAP7_75t_L g1087 ( .A(n_1060), .Y(n_1087) );
NAND2xp5_ASAP7_75t_SL g1088 ( .A(n_1052), .B(n_891), .Y(n_1088) );
INVx1_ASAP7_75t_SL g1089 ( .A(n_980), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_989), .Y(n_1090) );
INVx2_ASAP7_75t_L g1091 ( .A(n_986), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1005), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1000), .B(n_928), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1054), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1021), .Y(n_1095) );
AND3x2_ASAP7_75t_L g1096 ( .A(n_1020), .B(n_877), .C(n_930), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1000), .B(n_859), .Y(n_1097) );
NAND3xp33_ASAP7_75t_L g1098 ( .A(n_1018), .B(n_888), .C(n_944), .Y(n_1098) );
INVx1_ASAP7_75t_SL g1099 ( .A(n_1056), .Y(n_1099) );
AOI211xp5_ASAP7_75t_L g1100 ( .A1(n_1039), .A2(n_874), .B(n_886), .C(n_894), .Y(n_1100) );
AOI221xp5_ASAP7_75t_L g1101 ( .A1(n_1009), .A2(n_910), .B1(n_923), .B2(n_939), .C(n_858), .Y(n_1101) );
NAND2xp67_ASAP7_75t_L g1102 ( .A(n_1012), .B(n_860), .Y(n_1102) );
INVx2_ASAP7_75t_L g1103 ( .A(n_986), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1032), .Y(n_1104) );
INVx2_ASAP7_75t_L g1105 ( .A(n_988), .Y(n_1105) );
HB1xp67_ASAP7_75t_L g1106 ( .A(n_990), .Y(n_1106) );
NAND3xp33_ASAP7_75t_SL g1107 ( .A(n_1010), .B(n_914), .C(n_868), .Y(n_1107) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_1029), .B(n_859), .Y(n_1108) );
BUFx2_ASAP7_75t_L g1109 ( .A(n_1046), .Y(n_1109) );
OAI221xp5_ASAP7_75t_L g1110 ( .A1(n_1027), .A2(n_858), .B1(n_869), .B2(n_868), .C(n_881), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1038), .Y(n_1111) );
BUFx2_ASAP7_75t_L g1112 ( .A(n_1016), .Y(n_1112) );
AO21x2_ASAP7_75t_L g1113 ( .A1(n_1036), .A2(n_970), .B(n_969), .Y(n_1113) );
AOI22xp33_ASAP7_75t_SL g1114 ( .A1(n_1052), .A2(n_969), .B1(n_954), .B2(n_859), .Y(n_1114) );
OAI21xp5_ASAP7_75t_SL g1115 ( .A1(n_1064), .A2(n_869), .B(n_897), .Y(n_1115) );
OAI221xp5_ASAP7_75t_L g1116 ( .A1(n_983), .A2(n_1006), .B1(n_996), .B2(n_1025), .C(n_1014), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1034), .B(n_938), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1007), .B(n_952), .Y(n_1118) );
OAI31xp33_ASAP7_75t_L g1119 ( .A1(n_1008), .A2(n_955), .A3(n_945), .B(n_892), .Y(n_1119) );
AOI22xp5_ASAP7_75t_L g1120 ( .A1(n_1026), .A2(n_935), .B1(n_934), .B2(n_976), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1007), .B(n_952), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1034), .B(n_952), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_988), .B(n_952), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1026), .B(n_891), .Y(n_1124) );
OR2x2_ASAP7_75t_L g1125 ( .A(n_998), .B(n_891), .Y(n_1125) );
OR2x2_ASAP7_75t_L g1126 ( .A(n_998), .B(n_891), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1030), .Y(n_1127) );
NOR3xp33_ASAP7_75t_SL g1128 ( .A(n_1002), .B(n_924), .C(n_262), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1067), .B(n_859), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1019), .B(n_934), .Y(n_1130) );
OA21x2_ASAP7_75t_L g1131 ( .A1(n_1013), .A2(n_935), .B(n_972), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1030), .B(n_286), .Y(n_1132) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_1019), .B(n_261), .Y(n_1133) );
NOR2xp33_ASAP7_75t_SL g1134 ( .A(n_1031), .B(n_264), .Y(n_1134) );
AOI21xp5_ASAP7_75t_L g1135 ( .A1(n_1065), .A2(n_265), .B(n_266), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1035), .Y(n_1136) );
OR2x2_ASAP7_75t_L g1137 ( .A(n_1024), .B(n_267), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1010), .Y(n_1138) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1024), .Y(n_1139) );
AND2x4_ASAP7_75t_L g1140 ( .A(n_1069), .B(n_268), .Y(n_1140) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_1076), .Y(n_1141) );
NAND2x1p5_ASAP7_75t_L g1142 ( .A(n_1017), .B(n_269), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1011), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1051), .Y(n_1144) );
HB1xp67_ASAP7_75t_L g1145 ( .A(n_1069), .Y(n_1145) );
OAI31xp33_ASAP7_75t_SL g1146 ( .A1(n_982), .A2(n_270), .A3(n_271), .B(n_272), .Y(n_1146) );
OAI221xp5_ASAP7_75t_L g1147 ( .A1(n_996), .A2(n_273), .B1(n_274), .B2(n_276), .C(n_278), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1069), .B(n_995), .Y(n_1148) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1059), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1051), .Y(n_1150) );
INVx1_ASAP7_75t_SL g1151 ( .A(n_1056), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1152 ( .A(n_995), .B(n_280), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1068), .Y(n_1153) );
OAI33xp33_ASAP7_75t_L g1154 ( .A1(n_1004), .A2(n_282), .A3(n_283), .B1(n_284), .B2(n_984), .B3(n_997), .Y(n_1154) );
OA21x2_ASAP7_75t_L g1155 ( .A1(n_1059), .A2(n_1072), .B(n_981), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1081), .B(n_1071), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1001), .B(n_1071), .Y(n_1157) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1040), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_993), .B(n_1017), .Y(n_1159) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1040), .Y(n_1160) );
AOI221xp5_ASAP7_75t_L g1161 ( .A1(n_1025), .A2(n_1028), .B1(n_1023), .B2(n_1037), .C(n_994), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1017), .Y(n_1162) );
INVx2_ASAP7_75t_L g1163 ( .A(n_1040), .Y(n_1163) );
OAI221xp5_ASAP7_75t_L g1164 ( .A1(n_1015), .A2(n_991), .B1(n_1055), .B2(n_1041), .C(n_1043), .Y(n_1164) );
NAND3xp33_ASAP7_75t_L g1165 ( .A(n_1044), .B(n_1042), .C(n_1080), .Y(n_1165) );
HB1xp67_ASAP7_75t_L g1166 ( .A(n_1081), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1042), .B(n_1077), .Y(n_1167) );
INVx2_ASAP7_75t_L g1168 ( .A(n_1149), .Y(n_1168) );
INVxp67_ASAP7_75t_L g1169 ( .A(n_1109), .Y(n_1169) );
OR2x2_ASAP7_75t_L g1170 ( .A(n_1112), .B(n_987), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1097), .B(n_987), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1097), .B(n_999), .Y(n_1172) );
NOR2xp33_ASAP7_75t_L g1173 ( .A(n_1089), .B(n_1031), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1118), .B(n_999), .Y(n_1174) );
NAND4xp25_ASAP7_75t_L g1175 ( .A(n_1157), .B(n_1003), .C(n_1080), .D(n_1075), .Y(n_1175) );
INVxp67_ASAP7_75t_L g1176 ( .A(n_1109), .Y(n_1176) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1149), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1082), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1118), .B(n_999), .Y(n_1179) );
HB1xp67_ASAP7_75t_L g1180 ( .A(n_1112), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1083), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1121), .B(n_1053), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1086), .Y(n_1183) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1106), .B(n_1053), .Y(n_1184) );
NAND4xp25_ASAP7_75t_L g1185 ( .A(n_1157), .B(n_1075), .C(n_1061), .D(n_1079), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1121), .B(n_1072), .Y(n_1186) );
INVx1_ASAP7_75t_SL g1187 ( .A(n_1099), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1095), .Y(n_1188) );
AOI21xp5_ASAP7_75t_L g1189 ( .A1(n_1088), .A2(n_1022), .B(n_1074), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1083), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1084), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1093), .B(n_1070), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_1127), .B(n_1078), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1084), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1091), .B(n_1048), .Y(n_1195) );
NAND4xp25_ASAP7_75t_L g1196 ( .A(n_1107), .B(n_1066), .C(n_1063), .D(n_1058), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1093), .B(n_1047), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1123), .B(n_1049), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1104), .Y(n_1199) );
INVxp67_ASAP7_75t_SL g1200 ( .A(n_1108), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1123), .B(n_1050), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1090), .B(n_1062), .Y(n_1202) );
INVx1_ASAP7_75t_SL g1203 ( .A(n_1151), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_1154), .A2(n_1045), .B1(n_1073), .B2(n_1057), .Y(n_1204) );
INVx5_ASAP7_75t_L g1205 ( .A(n_1140), .Y(n_1205) );
OAI21xp5_ASAP7_75t_L g1206 ( .A1(n_1165), .A2(n_1164), .B(n_1128), .Y(n_1206) );
INVxp67_ASAP7_75t_L g1207 ( .A(n_1141), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1111), .Y(n_1208) );
NAND2xp33_ASAP7_75t_SL g1209 ( .A(n_1088), .B(n_1166), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1092), .B(n_1143), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_1091), .B(n_1103), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1103), .B(n_1139), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1105), .B(n_1139), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1105), .B(n_1130), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1094), .Y(n_1215) );
NOR2xp33_ASAP7_75t_L g1216 ( .A(n_1087), .B(n_1096), .Y(n_1216) );
INVx1_ASAP7_75t_SL g1217 ( .A(n_1108), .Y(n_1217) );
OR2x2_ASAP7_75t_L g1218 ( .A(n_1148), .B(n_1125), .Y(n_1218) );
INVx3_ASAP7_75t_SL g1219 ( .A(n_1140), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1136), .B(n_1138), .Y(n_1220) );
NOR3xp33_ASAP7_75t_SL g1221 ( .A(n_1116), .B(n_1115), .C(n_1110), .Y(n_1221) );
AOI21xp5_ASAP7_75t_L g1222 ( .A1(n_1167), .A2(n_1114), .B(n_1146), .Y(n_1222) );
HB1xp67_ASAP7_75t_L g1223 ( .A(n_1145), .Y(n_1223) );
INVx3_ASAP7_75t_SL g1224 ( .A(n_1140), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1159), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1159), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1130), .B(n_1148), .Y(n_1227) );
HB1xp67_ASAP7_75t_L g1228 ( .A(n_1122), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1125), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1144), .B(n_1150), .Y(n_1230) );
NAND4xp25_ASAP7_75t_L g1231 ( .A(n_1161), .B(n_1100), .C(n_1134), .D(n_1098), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1126), .B(n_1156), .Y(n_1232) );
NOR2xp33_ASAP7_75t_L g1233 ( .A(n_1162), .B(n_1124), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1227), .B(n_1126), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1181), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1227), .B(n_1163), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1181), .Y(n_1237) );
OR2x2_ASAP7_75t_L g1238 ( .A(n_1218), .B(n_1129), .Y(n_1238) );
AOI22xp5_ASAP7_75t_L g1239 ( .A1(n_1231), .A2(n_1085), .B1(n_1156), .B2(n_1153), .Y(n_1239) );
NOR2x1_ASAP7_75t_L g1240 ( .A(n_1187), .B(n_1137), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1225), .B(n_1102), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1218), .B(n_1226), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1190), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1171), .B(n_1163), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1171), .B(n_1160), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1230), .B(n_1102), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1190), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1232), .B(n_1160), .Y(n_1248) );
NAND4xp25_ASAP7_75t_L g1249 ( .A(n_1206), .B(n_1119), .C(n_1152), .D(n_1120), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1180), .B(n_1117), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1220), .B(n_1137), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1232), .B(n_1174), .Y(n_1252) );
INVxp67_ASAP7_75t_L g1253 ( .A(n_1203), .Y(n_1253) );
INVx1_ASAP7_75t_SL g1254 ( .A(n_1219), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1207), .B(n_1133), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1191), .Y(n_1256) );
HB1xp67_ASAP7_75t_L g1257 ( .A(n_1217), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1210), .B(n_1133), .Y(n_1258) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_1200), .B(n_1158), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1191), .Y(n_1260) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1168), .Y(n_1261) );
NOR2x1_ASAP7_75t_L g1262 ( .A(n_1175), .B(n_1152), .Y(n_1262) );
OAI22xp5_ASAP7_75t_L g1263 ( .A1(n_1219), .A2(n_1142), .B1(n_1147), .B2(n_1132), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1172), .B(n_1155), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1172), .B(n_1155), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1194), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1174), .B(n_1179), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1169), .B(n_1131), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1176), .B(n_1228), .Y(n_1269) );
INVx1_ASAP7_75t_SL g1270 ( .A(n_1173), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1229), .B(n_1131), .Y(n_1271) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1168), .Y(n_1272) );
AOI21xp5_ASAP7_75t_L g1273 ( .A1(n_1209), .A2(n_1135), .B(n_1113), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1179), .B(n_1155), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1178), .B(n_1131), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1183), .B(n_1113), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1188), .B(n_1113), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1242), .B(n_1208), .Y(n_1278) );
NOR2xp33_ASAP7_75t_L g1279 ( .A(n_1270), .B(n_1216), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_1249), .A2(n_1222), .B1(n_1197), .B2(n_1192), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1281 ( .A(n_1242), .B(n_1199), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1267), .B(n_1214), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1235), .Y(n_1283) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1261), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1267), .B(n_1214), .Y(n_1285) );
NOR2xp33_ASAP7_75t_L g1286 ( .A(n_1253), .B(n_1193), .Y(n_1286) );
OAI321xp33_ASAP7_75t_L g1287 ( .A1(n_1249), .A2(n_1196), .A3(n_1185), .B1(n_1170), .B2(n_1233), .C(n_1184), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1250), .B(n_1215), .Y(n_1288) );
AND4x1_ASAP7_75t_L g1289 ( .A(n_1262), .B(n_1221), .C(n_1189), .D(n_1204), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_1252), .B(n_1170), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1234), .B(n_1223), .Y(n_1291) );
OR2x2_ASAP7_75t_L g1292 ( .A(n_1252), .B(n_1211), .Y(n_1292) );
INVxp33_ASAP7_75t_L g1293 ( .A(n_1257), .Y(n_1293) );
INVxp67_ASAP7_75t_SL g1294 ( .A(n_1240), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1295 ( .A(n_1269), .B(n_1211), .Y(n_1295) );
OAI22xp5_ASAP7_75t_L g1296 ( .A1(n_1262), .A2(n_1224), .B1(n_1205), .B2(n_1184), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1235), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1236), .B(n_1212), .Y(n_1298) );
OAI21xp5_ASAP7_75t_SL g1299 ( .A1(n_1254), .A2(n_1142), .B(n_1224), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1248), .B(n_1182), .Y(n_1300) );
AOI21xp5_ASAP7_75t_L g1301 ( .A1(n_1263), .A2(n_1209), .B(n_1205), .Y(n_1301) );
INVx2_ASAP7_75t_L g1302 ( .A(n_1261), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1237), .Y(n_1303) );
INVx2_ASAP7_75t_SL g1304 ( .A(n_1254), .Y(n_1304) );
XOR2x2_ASAP7_75t_L g1305 ( .A(n_1239), .B(n_1202), .Y(n_1305) );
OAI211xp5_ASAP7_75t_L g1306 ( .A1(n_1239), .A2(n_1205), .B(n_1182), .C(n_1201), .Y(n_1306) );
OA22x2_ASAP7_75t_L g1307 ( .A1(n_1246), .A2(n_1201), .B1(n_1198), .B2(n_1194), .Y(n_1307) );
INVx2_ASAP7_75t_SL g1308 ( .A(n_1259), .Y(n_1308) );
XNOR2x1_ASAP7_75t_L g1309 ( .A(n_1238), .B(n_1198), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1271), .B(n_1212), .Y(n_1310) );
HB1xp67_ASAP7_75t_L g1311 ( .A(n_1259), .Y(n_1311) );
AOI21xp5_ASAP7_75t_L g1312 ( .A1(n_1240), .A2(n_1205), .B(n_1195), .Y(n_1312) );
OAI22xp5_ASAP7_75t_L g1313 ( .A1(n_1258), .A2(n_1205), .B1(n_1195), .B2(n_1177), .Y(n_1313) );
AOI211xp5_ASAP7_75t_L g1314 ( .A1(n_1241), .A2(n_1186), .B(n_1101), .C(n_1213), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1237), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1238), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1317 ( .A(n_1275), .B(n_1186), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1243), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1268), .B(n_1244), .Y(n_1319) );
NAND2xp5_ASAP7_75t_L g1320 ( .A(n_1245), .B(n_1251), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1243), .Y(n_1321) );
AOI32xp33_ASAP7_75t_L g1322 ( .A1(n_1264), .A2(n_1274), .A3(n_1265), .B1(n_1255), .B2(n_1266), .Y(n_1322) );
O2A1O1Ixp33_ASAP7_75t_L g1323 ( .A1(n_1287), .A2(n_1280), .B(n_1279), .C(n_1304), .Y(n_1323) );
AOI211xp5_ASAP7_75t_L g1324 ( .A1(n_1287), .A2(n_1299), .B(n_1296), .C(n_1306), .Y(n_1324) );
NAND4xp25_ASAP7_75t_SL g1325 ( .A(n_1322), .B(n_1301), .C(n_1312), .D(n_1314), .Y(n_1325) );
AOI21xp5_ASAP7_75t_L g1326 ( .A1(n_1299), .A2(n_1307), .B(n_1294), .Y(n_1326) );
NOR2x1_ASAP7_75t_L g1327 ( .A(n_1309), .B(n_1286), .Y(n_1327) );
OAI321xp33_ASAP7_75t_L g1328 ( .A1(n_1313), .A2(n_1308), .A3(n_1289), .B1(n_1317), .B2(n_1290), .C(n_1265), .Y(n_1328) );
AOI22x1_ASAP7_75t_L g1329 ( .A1(n_1311), .A2(n_1308), .B1(n_1289), .B2(n_1290), .Y(n_1329) );
NAND2xp5_ASAP7_75t_SL g1330 ( .A(n_1293), .B(n_1305), .Y(n_1330) );
AOI221xp5_ASAP7_75t_L g1331 ( .A1(n_1288), .A2(n_1316), .B1(n_1278), .B2(n_1281), .C(n_1319), .Y(n_1331) );
NOR2xp33_ASAP7_75t_R g1332 ( .A(n_1291), .B(n_1295), .Y(n_1332) );
INVxp67_ASAP7_75t_L g1333 ( .A(n_1295), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1333), .Y(n_1334) );
AO22x2_ASAP7_75t_L g1335 ( .A1(n_1330), .A2(n_1273), .B1(n_1292), .B2(n_1285), .Y(n_1335) );
NOR3xp33_ASAP7_75t_SL g1336 ( .A(n_1325), .B(n_1276), .C(n_1277), .Y(n_1336) );
HB1xp67_ASAP7_75t_L g1337 ( .A(n_1332), .Y(n_1337) );
AOI221xp5_ASAP7_75t_L g1338 ( .A1(n_1328), .A2(n_1320), .B1(n_1310), .B2(n_1318), .C(n_1321), .Y(n_1338) );
AOI21xp5_ASAP7_75t_L g1339 ( .A1(n_1326), .A2(n_1298), .B(n_1282), .Y(n_1339) );
NAND2xp5_ASAP7_75t_SL g1340 ( .A(n_1329), .B(n_1284), .Y(n_1340) );
AOI21x1_ASAP7_75t_L g1341 ( .A1(n_1337), .A2(n_1327), .B(n_1323), .Y(n_1341) );
OAI22x1_ASAP7_75t_L g1342 ( .A1(n_1340), .A2(n_1324), .B1(n_1332), .B2(n_1331), .Y(n_1342) );
OAI221xp5_ASAP7_75t_L g1343 ( .A1(n_1336), .A2(n_1315), .B1(n_1303), .B2(n_1297), .C(n_1283), .Y(n_1343) );
OAI211xp5_ASAP7_75t_L g1344 ( .A1(n_1338), .A2(n_1283), .B(n_1297), .C(n_1300), .Y(n_1344) );
INVx5_ASAP7_75t_L g1345 ( .A(n_1341), .Y(n_1345) );
NOR3xp33_ASAP7_75t_SL g1346 ( .A(n_1344), .B(n_1339), .C(n_1334), .Y(n_1346) );
INVx2_ASAP7_75t_SL g1347 ( .A(n_1342), .Y(n_1347) );
NOR2x1_ASAP7_75t_L g1348 ( .A(n_1343), .B(n_1335), .Y(n_1348) );
INVx1_ASAP7_75t_SL g1349 ( .A(n_1347), .Y(n_1349) );
NAND3xp33_ASAP7_75t_L g1350 ( .A(n_1345), .B(n_1346), .C(n_1348), .Y(n_1350) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1349), .Y(n_1351) );
XNOR2xp5_ASAP7_75t_L g1352 ( .A(n_1350), .B(n_1335), .Y(n_1352) );
OAI21xp5_ASAP7_75t_L g1353 ( .A1(n_1352), .A2(n_1302), .B(n_1284), .Y(n_1353) );
AOI222xp33_ASAP7_75t_L g1354 ( .A1(n_1351), .A2(n_1247), .B1(n_1256), .B2(n_1260), .C1(n_1266), .C2(n_1302), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1353), .Y(n_1355) );
AOI21xp5_ASAP7_75t_L g1356 ( .A1(n_1355), .A2(n_1354), .B(n_1272), .Y(n_1356) );
endmodule