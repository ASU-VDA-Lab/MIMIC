module real_jpeg_23849_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_288;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

INVx6_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_2),
.A2(n_39),
.B1(n_66),
.B2(n_67),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_2),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_3),
.A2(n_52),
.B1(n_66),
.B2(n_67),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_7),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_55),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_7),
.A2(n_55),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_8),
.A2(n_66),
.B1(n_67),
.B2(n_80),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_80),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_9),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_110),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_110),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_9),
.A2(n_66),
.B1(n_67),
.B2(n_110),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_11),
.B(n_43),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_11),
.B(n_66),
.C(n_74),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_159),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_11),
.B(n_107),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_11),
.A2(n_69),
.B1(n_177),
.B2(n_230),
.Y(n_229)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_13),
.A2(n_156),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_13),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_164),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_164),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_13),
.A2(n_66),
.B1(n_67),
.B2(n_164),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_15),
.A2(n_42),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_42),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_15),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_139),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_137),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_19),
.B(n_111),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_82),
.C(n_91),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_20),
.B(n_82),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_58),
.B2(n_81),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_44),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_23),
.B(n_44),
.C(n_81),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_37),
.B(n_40),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_24),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_24),
.A2(n_26),
.B1(n_162),
.B2(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_25),
.A2(n_38),
.B1(n_43),
.B2(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_25),
.A2(n_43),
.B1(n_155),
.B2(n_161),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_36),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_27),
.A2(n_30),
.B(n_160),
.C(n_179),
.Y(n_178)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_28),
.B(n_29),
.C(n_36),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_29),
.A2(n_30),
.B1(n_46),
.B2(n_50),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g245 ( 
.A(n_30),
.B(n_159),
.CON(n_245),
.SN(n_245)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_30),
.B(n_47),
.C(n_50),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_35),
.Y(n_123)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_35),
.Y(n_158)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_36),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_41),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_43),
.B(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_51),
.B(n_53),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_45),
.A2(n_105),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_45)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_46),
.A2(n_48),
.B(n_245),
.C(n_246),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_48),
.B1(n_74),
.B2(n_76),
.Y(n_73)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_48),
.B(n_204),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_51),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_54),
.B(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_56),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_56),
.A2(n_107),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_56),
.A2(n_107),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_56),
.A2(n_107),
.B1(n_189),
.B2(n_245),
.Y(n_254)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_71),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_59),
.A2(n_60),
.B1(n_71),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_62),
.A2(n_69),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_63),
.Y(n_177)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_66),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_69),
.B(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g195 ( 
.A(n_64),
.Y(n_195)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_64),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_65),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_65),
.A2(n_96),
.B(n_221),
.Y(n_247)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_67),
.B1(n_74),
.B2(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_67),
.B(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_68),
.A2(n_176),
.B(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_69),
.A2(n_94),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_69),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_69),
.A2(n_97),
.B1(n_223),
.B2(n_230),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_97),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_71),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_79),
.B(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_72),
.A2(n_87),
.B(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_72),
.A2(n_77),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_72),
.A2(n_77),
.B1(n_208),
.B2(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_72),
.A2(n_129),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_78),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_77),
.B(n_159),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_86),
.B2(n_90),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_84),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_86),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_89),
.B(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_89),
.A2(n_100),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_91),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_101),
.C(n_108),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_92),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_93),
.B(n_98),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_101),
.A2(n_102),
.B1(n_108),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B(n_106),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_104),
.B(n_107),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_105),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_108),
.Y(n_283)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_136),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_126),
.B2(n_127),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_125),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_123),
.B(n_159),
.Y(n_160)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_131),
.B(n_135),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_290),
.B(n_294),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_196),
.B(n_277),
.C(n_289),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_181),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_142),
.B(n_181),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_165),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_144),
.B(n_147),
.C(n_165),
.Y(n_278)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.C(n_154),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_152),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_154),
.B(n_183),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_159),
.B(n_160),
.Y(n_155)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_159),
.B(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_173),
.B2(n_180),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_168),
.B(n_170),
.C(n_180),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_173),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_178),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.C(n_186),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_182),
.B(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_185),
.B(n_186),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.C(n_193),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_187),
.B(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_221),
.B1(n_222),
.B2(n_224),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_276),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_271),
.B(n_275),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_257),
.B(n_270),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_241),
.B(n_256),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_218),
.B(n_240),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_209),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_205),
.B1(n_206),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_216),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_214),
.C(n_216),
.Y(n_255)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_217),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_227),
.B(n_239),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_225),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_235),
.B(n_238),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_255),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_255),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_250),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_251),
.C(n_254),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_253),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_258),
.B(n_259),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_266),
.C(n_268),
.Y(n_274)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_274),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_279),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_288),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_284),
.B1(n_286),
.B2(n_287),
.Y(n_280)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_281),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_286),
.C(n_288),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);


endmodule