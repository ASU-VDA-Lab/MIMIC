module real_jpeg_26316_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_1),
.A2(n_19),
.B1(n_21),
.B2(n_56),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_1),
.B(n_24),
.C(n_29),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_39),
.B1(n_88),
.B2(n_95),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_4),
.A2(n_19),
.B1(n_21),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_5),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_20),
.B1(n_52),
.B2(n_53),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_5),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_9),
.A2(n_19),
.B1(n_21),
.B2(n_44),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_11),
.Y(n_89)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_11),
.Y(n_98)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_72),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_70),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_49),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_15),
.B(n_49),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_33),
.C(n_38),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_16),
.A2(n_17),
.B1(n_33),
.B2(n_34),
.Y(n_80)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_18),
.A2(n_22),
.B1(n_30),
.B2(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_19),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_23)
);

AO22x1_ASAP7_75t_L g35 ( 
.A1(n_19),
.A2(n_21),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g51 ( 
.A1(n_19),
.A2(n_36),
.A3(n_52),
.B1(n_55),
.B2(n_57),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_19),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_21),
.B(n_37),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_22),
.A2(n_30),
.B1(n_31),
.B2(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.Y(n_22)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_27),
.B(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_28),
.B(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_55),
.B1(n_67),
.B2(n_69),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_36),
.A2(n_37),
.B1(n_52),
.B2(n_53),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B(n_45),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_59),
.B(n_60),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_39),
.A2(n_85),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_40),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_63),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

HAxp5_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_56),
.CON(n_55),
.SN(n_55)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_81),
.B(n_106),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_74),
.B(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_77),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_91),
.B(n_105),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_90),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_90),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_99),
.B(n_104),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);


endmodule