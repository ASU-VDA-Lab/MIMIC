module fake_jpeg_439_n_186 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_1),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_28),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_42),
.C(n_23),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_75),
.Y(n_86)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_46),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_60),
.Y(n_83)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_62),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_86),
.Y(n_91)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_18),
.A3(n_43),
.B1(n_41),
.B2(n_40),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_75),
.C(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_93),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_49),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_108),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_50),
.B1(n_60),
.B2(n_59),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_54),
.B1(n_52),
.B2(n_58),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_68),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_61),
.Y(n_116)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_67),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_33),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_71),
.B1(n_84),
.B2(n_72),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_44),
.B1(n_39),
.B2(n_38),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_72),
.B(n_69),
.C(n_64),
.Y(n_111)
);

INVxp33_ASAP7_75t_SL g146 ( 
.A(n_111),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_62),
.B(n_63),
.C(n_56),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_114),
.B(n_126),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_66),
.B(n_64),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_124),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_55),
.B(n_57),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_4),
.B(n_5),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_65),
.B1(n_69),
.B2(n_54),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_120),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_55),
.Y(n_120)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_97),
.B1(n_98),
.B2(n_2),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_25),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_97),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_129),
.C(n_144),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_32),
.C(n_30),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_0),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_0),
.Y(n_137)
);

OAI21x1_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_1),
.B(n_2),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_138),
.A2(n_143),
.B(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_4),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_140),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_24),
.C(n_21),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_20),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_19),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_8),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_5),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_9),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_157),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_150),
.B(n_153),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_119),
.B(n_7),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_158),
.B(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_148),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_141),
.B1(n_151),
.B2(n_152),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_156),
.B(n_161),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_131),
.A2(n_16),
.B(n_10),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_162),
.A2(n_133),
.B1(n_146),
.B2(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_164),
.B(n_170),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_165),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_142),
.B1(n_13),
.B2(n_14),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_129),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_159),
.C(n_156),
.Y(n_171)
);

BUFx12_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_175),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_159),
.C(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_176),
.B(n_168),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_178),
.A2(n_15),
.B1(n_170),
.B2(n_177),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_163),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_174),
.B(n_172),
.C(n_180),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g184 ( 
.A(n_183),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_182),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_170),
.Y(n_186)
);


endmodule