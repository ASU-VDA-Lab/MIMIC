module fake_jpeg_134_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_0),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx2_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_35),
.B1(n_43),
.B2(n_41),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_62),
.B1(n_56),
.B2(n_55),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_40),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_36),
.C(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_37),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_63),
.B(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_75),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_61),
.B1(n_38),
.B2(n_41),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_89),
.B1(n_1),
.B2(n_2),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_81),
.B(n_83),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_1),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_62),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_77),
.C(n_85),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_44),
.B1(n_42),
.B2(n_39),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_67),
.B1(n_65),
.B2(n_46),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_76),
.B1(n_57),
.B2(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_34),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_95),
.C(n_97),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_86),
.B(n_87),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_2),
.B(n_3),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_33),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_98),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_102),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_101),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_25),
.B1(n_24),
.B2(n_23),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_97),
.B(n_18),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_110),
.C(n_5),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_100),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_16),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_6),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_4),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_113),
.B(n_102),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_117),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_118),
.B(n_120),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_5),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_15),
.C(n_7),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_121),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_108),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_119),
.A2(n_105),
.B1(n_104),
.B2(n_103),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_126),
.A2(n_106),
.B(n_110),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_114),
.B(n_109),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_123),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_129),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_125),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_6),
.C2(n_12),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_131),
.C(n_12),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_13),
.C(n_14),
.Y(n_135)
);


endmodule