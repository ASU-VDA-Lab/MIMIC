module fake_jpeg_29685_n_538 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_538);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_538;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_20),
.B(n_7),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_47),
.C(n_48),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_7),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_59),
.B(n_69),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_64),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_22),
.B(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_68),
.B(n_85),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_37),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_83),
.Y(n_155)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_7),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_23),
.B(n_8),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_24),
.A2(n_6),
.B1(n_13),
.B2(n_2),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_53),
.B1(n_40),
.B2(n_45),
.Y(n_129)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

BUFx4f_ASAP7_75t_SL g156 ( 
.A(n_100),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_24),
.B(n_6),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_30),
.B(n_6),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_105),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_40),
.B(n_9),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_84),
.A2(n_26),
.B1(n_46),
.B2(n_44),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_120),
.A2(n_144),
.B1(n_92),
.B2(n_90),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_69),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_123),
.B(n_126),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_53),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_127),
.B(n_150),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_129),
.A2(n_138),
.B1(n_49),
.B2(n_51),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_45),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_132),
.B(n_137),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_47),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_86),
.A2(n_44),
.B1(n_33),
.B2(n_37),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_54),
.A2(n_44),
.B1(n_33),
.B2(n_48),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_140),
.A2(n_87),
.B1(n_93),
.B2(n_78),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_145),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_91),
.A2(n_44),
.B1(n_33),
.B2(n_48),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_65),
.B(n_28),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_103),
.Y(n_150)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_155),
.A2(n_67),
.B1(n_66),
.B2(n_100),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_168),
.A2(n_217),
.B1(n_218),
.B2(n_151),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_116),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_169),
.B(n_181),
.Y(n_223)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_170),
.Y(n_241)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

BUFx4f_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_172),
.Y(n_255)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_175),
.B(n_176),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_122),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_166),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_177),
.B(n_178),
.Y(n_233)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_39),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_180),
.B(n_187),
.Y(n_248)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_155),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_189),
.B(n_190),
.Y(n_256)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_134),
.A2(n_39),
.B1(n_52),
.B2(n_51),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_197),
.Y(n_235)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_194),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_148),
.B(n_38),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_198),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_106),
.B(n_35),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_200),
.Y(n_257)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_143),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_134),
.B(n_112),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_136),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_211),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_111),
.B(n_83),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_213),
.Y(n_254)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_135),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_62),
.B1(n_56),
.B2(n_72),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_35),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_216),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_125),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_113),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_141),
.B(n_43),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_219),
.B(n_220),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_157),
.B(n_28),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_138),
.B(n_52),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_43),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_236),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_38),
.B(n_18),
.C(n_29),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_234),
.B(n_29),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_109),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_181),
.A2(n_152),
.B1(n_154),
.B2(n_131),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_238),
.A2(n_244),
.B1(n_262),
.B2(n_263),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_204),
.A2(n_120),
.B(n_144),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_243),
.A2(n_168),
.B(n_166),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_109),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_260),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_173),
.B(n_124),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_214),
.A2(n_114),
.B1(n_124),
.B2(n_119),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_191),
.A2(n_140),
.B1(n_64),
.B2(n_74),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_130),
.B1(n_114),
.B2(n_164),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_265),
.A2(n_280),
.B1(n_287),
.B2(n_255),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_242),
.A2(n_217),
.B1(n_203),
.B2(n_174),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_266),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_237),
.A2(n_209),
.B1(n_205),
.B2(n_171),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_268),
.A2(n_283),
.B(n_292),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_215),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_271),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_204),
.C(n_212),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_294),
.C(n_222),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_199),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_272),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_275),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_223),
.A2(n_131),
.B1(n_154),
.B2(n_213),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_277),
.A2(n_289),
.B1(n_293),
.B2(n_296),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_228),
.B(n_200),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_290),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_279),
.B(n_284),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_235),
.A2(n_211),
.B1(n_149),
.B2(n_60),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_286),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_235),
.A2(n_193),
.B1(n_185),
.B2(n_192),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_241),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_288),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_235),
.A2(n_218),
.B1(n_195),
.B2(n_184),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_239),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_227),
.B(n_186),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_260),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_243),
.A2(n_223),
.B(n_254),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_223),
.A2(n_216),
.B1(n_179),
.B2(n_182),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_201),
.C(n_194),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_258),
.A2(n_156),
.B(n_49),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_295),
.A2(n_229),
.B(n_172),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_236),
.A2(n_133),
.B1(n_157),
.B2(n_33),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_230),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_237),
.A2(n_183),
.B1(n_188),
.B2(n_169),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_255),
.B1(n_172),
.B2(n_242),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_263),
.A2(n_125),
.B1(n_70),
.B2(n_33),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_299),
.A2(n_255),
.B1(n_222),
.B2(n_259),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_306),
.B(n_44),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_244),
.B1(n_233),
.B2(n_242),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_307),
.A2(n_320),
.B1(n_282),
.B2(n_232),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_233),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_308),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_309),
.B(n_310),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_279),
.B(n_230),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_331),
.Y(n_363)
);

NAND3xp33_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_225),
.C(n_248),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_L g343 ( 
.A1(n_312),
.A2(n_264),
.B(n_267),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_313),
.A2(n_319),
.B(n_298),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_248),
.C(n_231),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_294),
.C(n_269),
.Y(n_339)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_322),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_292),
.A2(n_229),
.B(n_234),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_323),
.A2(n_334),
.B(n_295),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_325),
.A2(n_333),
.B1(n_265),
.B2(n_290),
.Y(n_345)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_326),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_249),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_327),
.Y(n_347)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_275),
.Y(n_328)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_328),
.Y(n_342)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_285),
.Y(n_329)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_329),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_276),
.A2(n_237),
.B1(n_259),
.B2(n_239),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_276),
.A2(n_249),
.B1(n_240),
.B2(n_232),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_283),
.A2(n_252),
.B(n_246),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_336),
.A2(n_341),
.B(n_350),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_337),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_301),
.B(n_291),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_338),
.B(n_351),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_356),
.C(n_367),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_303),
.A2(n_281),
.B(n_287),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_343),
.B(n_361),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_304),
.A2(n_267),
.B1(n_280),
.B2(n_264),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_344),
.A2(n_345),
.B1(n_349),
.B2(n_351),
.Y(n_385)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_318),
.Y(n_349)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_349),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_324),
.A2(n_293),
.B1(n_296),
.B2(n_299),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_318),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_352),
.A2(n_304),
.B1(n_325),
.B2(n_320),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_303),
.A2(n_288),
.B(n_290),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_353),
.A2(n_354),
.B(n_355),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_319),
.A2(n_288),
.B(n_268),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_334),
.A2(n_247),
.B(n_246),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_306),
.B(n_247),
.C(n_252),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_308),
.A2(n_156),
.B(n_241),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_357),
.A2(n_366),
.B(n_314),
.Y(n_397)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_302),
.Y(n_360)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_308),
.A2(n_286),
.B(n_226),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_302),
.Y(n_362)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_315),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_365),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_300),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_324),
.A2(n_183),
.B(n_226),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_315),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_368),
.B(n_332),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_399),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_311),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_373),
.B(n_377),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_346),
.A2(n_323),
.B1(n_305),
.B2(n_322),
.Y(n_374)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_316),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_359),
.A2(n_305),
.B1(n_331),
.B2(n_333),
.Y(n_378)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_378),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_326),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_379),
.B(n_391),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_346),
.B(n_330),
.Y(n_380)
);

NAND3xp33_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_340),
.C(n_360),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_329),
.Y(n_381)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

NAND2x1p5_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_328),
.Y(n_382)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_382),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_321),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_348),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_385),
.A2(n_392),
.B1(n_376),
.B2(n_378),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_347),
.B(n_330),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_386),
.B(n_398),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_363),
.A2(n_321),
.B1(n_317),
.B2(n_314),
.Y(n_389)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_389),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_336),
.B(n_317),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_257),
.C(n_332),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_392),
.B(n_368),
.C(n_340),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_357),
.B(n_341),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_19),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_355),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_335),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_335),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_400),
.B(n_342),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_352),
.A2(n_300),
.B1(n_273),
.B2(n_282),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_401),
.B(n_345),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_382),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_403),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_381),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_404),
.B(n_406),
.Y(n_445)
);

INVx13_ASAP7_75t_L g406 ( 
.A(n_395),
.Y(n_406)
);

AOI322xp5_ASAP7_75t_L g407 ( 
.A1(n_371),
.A2(n_337),
.A3(n_353),
.B1(n_338),
.B2(n_354),
.C1(n_350),
.C2(n_364),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_407),
.A2(n_369),
.B1(n_397),
.B2(n_396),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_408),
.Y(n_432)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_410),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_411),
.A2(n_422),
.B(n_396),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_373),
.C(n_375),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_348),
.Y(n_415)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_379),
.B(n_362),
.Y(n_416)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_416),
.Y(n_447)
);

XOR2x2_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_366),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_389),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_421),
.B(n_429),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_376),
.A2(n_342),
.B(n_365),
.Y(n_422)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_423),
.Y(n_448)
);

INVx13_ASAP7_75t_L g425 ( 
.A(n_395),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_427),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_372),
.B(n_358),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_393),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_428),
.B(n_415),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_430),
.A2(n_370),
.B1(n_394),
.B2(n_391),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_431),
.B(n_453),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_433),
.A2(n_411),
.B(n_417),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_421),
.Y(n_455)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_414),
.B(n_375),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_442),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_385),
.Y(n_441)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_441),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_377),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_443),
.A2(n_450),
.B1(n_454),
.B2(n_413),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_444),
.B(n_452),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_390),
.Y(n_449)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_449),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_409),
.A2(n_401),
.B1(n_382),
.B2(n_387),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_413),
.B(n_273),
.Y(n_451)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_170),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_224),
.C(n_19),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_402),
.A2(n_224),
.B1(n_1),
.B2(n_0),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_470),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_432),
.B(n_429),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_457),
.Y(n_489)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_448),
.Y(n_457)
);

FAx1_ASAP7_75t_SL g458 ( 
.A(n_439),
.B(n_422),
.CI(n_411),
.CON(n_458),
.SN(n_458)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_458),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_460),
.B(n_436),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_466),
.A2(n_444),
.B1(n_417),
.B2(n_443),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_446),
.A2(n_402),
.B1(n_426),
.B2(n_418),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_473),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_412),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_437),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_447),
.Y(n_469)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_469),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_419),
.Y(n_470)
);

BUFx24_ASAP7_75t_SL g471 ( 
.A(n_440),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_471),
.A2(n_464),
.B(n_465),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_442),
.B(n_426),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_476),
.B(n_480),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_461),
.A2(n_438),
.B1(n_446),
.B2(n_419),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_477),
.A2(n_478),
.B1(n_488),
.B2(n_490),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_452),
.C(n_433),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_482),
.C(n_487),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_450),
.C(n_451),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_463),
.A2(n_441),
.B1(n_405),
.B2(n_410),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_483),
.A2(n_479),
.B1(n_485),
.B2(n_487),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_486),
.Y(n_505)
);

OAI21xp33_ASAP7_75t_L g486 ( 
.A1(n_458),
.A2(n_403),
.B(n_449),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_462),
.B(n_439),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_472),
.A2(n_473),
.B1(n_462),
.B2(n_405),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_467),
.A2(n_454),
.B1(n_435),
.B2(n_427),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_459),
.B(n_453),
.C(n_435),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_32),
.C(n_9),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_475),
.A2(n_460),
.B1(n_459),
.B2(n_425),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_493),
.A2(n_499),
.B1(n_495),
.B2(n_497),
.Y(n_513)
);

BUFx24_ASAP7_75t_SL g494 ( 
.A(n_489),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g511 ( 
.A(n_494),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_486),
.A2(n_406),
.B1(n_224),
.B2(n_49),
.Y(n_495)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_495),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_484),
.A2(n_224),
.B(n_11),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_497),
.A2(n_506),
.B(n_12),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_498),
.B(n_504),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_477),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_474),
.A2(n_11),
.B(n_15),
.Y(n_500)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_500),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_481),
.A2(n_11),
.B(n_15),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_501),
.A2(n_503),
.B(n_491),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_480),
.B(n_32),
.C(n_1),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_482),
.A2(n_5),
.B(n_13),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_513),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_509),
.B(n_515),
.Y(n_525)
);

MAJx2_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_485),
.C(n_12),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_506),
.C(n_498),
.Y(n_523)
);

BUFx24_ASAP7_75t_SL g512 ( 
.A(n_496),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_512),
.B(n_517),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_492),
.A2(n_2),
.B(n_3),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_3),
.Y(n_521)
);

BUFx24_ASAP7_75t_SL g517 ( 
.A(n_505),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_505),
.A2(n_3),
.B(n_12),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_493),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_521),
.B(n_523),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_502),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_522),
.A2(n_520),
.B(n_507),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_524),
.B(n_503),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_525),
.A2(n_511),
.B(n_32),
.Y(n_529)
);

AO21x1_ASAP7_75t_L g531 ( 
.A1(n_526),
.A2(n_528),
.B(n_529),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_527),
.A2(n_522),
.B(n_519),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_530),
.A2(n_532),
.B(n_32),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_528),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_531),
.C(n_1),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_534),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_12),
.B(n_13),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_0),
.C(n_32),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_0),
.Y(n_538)
);


endmodule