module fake_jpeg_18075_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g15 ( 
.A(n_12),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_40),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_51),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx2_ASAP7_75t_SL g58 ( 
.A(n_47),
.Y(n_58)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_23),
.B1(n_17),
.B2(n_26),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_39),
.B1(n_32),
.B2(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_63),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_68),
.B1(n_39),
.B2(n_50),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_67),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_70),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_30),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_42),
.B(n_27),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_70),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_41),
.A2(n_35),
.B1(n_37),
.B2(n_33),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_41),
.B1(n_44),
.B2(n_49),
.Y(n_104)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_26),
.B1(n_17),
.B2(n_23),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_89),
.B(n_96),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_95),
.B1(n_113),
.B2(n_56),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_41),
.B1(n_44),
.B2(n_49),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_35),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_110),
.Y(n_121)
);

AOI32xp33_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_33),
.A3(n_39),
.B1(n_32),
.B2(n_19),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_15),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_50),
.B1(n_77),
.B2(n_85),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_41),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_46),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_79),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_44),
.B1(n_23),
.B2(n_17),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_18),
.B(n_27),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_116),
.A2(n_126),
.B(n_131),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_117),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_50),
.B1(n_69),
.B2(n_76),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_129),
.B1(n_130),
.B2(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_128),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_136),
.B1(n_139),
.B2(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

AND2x4_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_32),
.Y(n_126)
);

OAI31xp33_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_24),
.A3(n_32),
.B(n_38),
.Y(n_127)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_140),
.B(n_82),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_62),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_91),
.A2(n_26),
.B1(n_56),
.B2(n_57),
.Y(n_130)
);

NOR2xp67_ASAP7_75t_R g131 ( 
.A(n_89),
.B(n_38),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_24),
.B(n_31),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g133 ( 
.A(n_108),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_106),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_34),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_72),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_80),
.B1(n_23),
.B2(n_34),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_36),
.B1(n_16),
.B2(n_27),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_137),
.A2(n_103),
.B1(n_100),
.B2(n_90),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_88),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_142),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_112),
.A2(n_36),
.B1(n_15),
.B2(n_38),
.Y(n_139)
);

AOI22x1_ASAP7_75t_L g140 ( 
.A1(n_87),
.A2(n_38),
.B1(n_36),
.B2(n_31),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_36),
.B1(n_15),
.B2(n_71),
.Y(n_141)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_114),
.B(n_86),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_152),
.B(n_161),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_86),
.C(n_114),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_28),
.C(n_82),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_146),
.B1(n_155),
.B2(n_122),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_111),
.B(n_103),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_172),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_22),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_168),
.C(n_20),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_100),
.B1(n_111),
.B2(n_105),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_105),
.B1(n_99),
.B2(n_94),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_SL g185 ( 
.A1(n_156),
.A2(n_160),
.B(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_119),
.A2(n_117),
.B(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_167),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_121),
.A2(n_24),
.B(n_31),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_164),
.A2(n_137),
.B(n_140),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_99),
.Y(n_166)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_127),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_22),
.C(n_31),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_140),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_31),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_20),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_16),
.B1(n_22),
.B2(n_82),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_16),
.B1(n_82),
.B2(n_21),
.Y(n_186)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_180),
.A2(n_197),
.B(n_202),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_139),
.Y(n_181)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_187),
.C(n_4),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_184),
.A2(n_206),
.B1(n_170),
.B2(n_174),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_205),
.B1(n_146),
.B2(n_165),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_28),
.C(n_21),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_29),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_190),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_20),
.B1(n_29),
.B2(n_2),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_192),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_193),
.B(n_195),
.Y(n_213)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_169),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_148),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_204),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_165),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_198)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_150),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_201),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_143),
.A2(n_0),
.B(n_1),
.Y(n_202)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_154),
.B(n_8),
.CI(n_13),
.CON(n_203),
.SN(n_203)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_173),
.A2(n_9),
.A3(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_204)
);

AOI22x1_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_3),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_208),
.A2(n_214),
.B1(n_210),
.B2(n_222),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_179),
.B1(n_182),
.B2(n_176),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_212),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_196),
.B(n_161),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_175),
.A2(n_157),
.B(n_160),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_205),
.B(n_204),
.Y(n_244)
);

FAx1_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_157),
.CI(n_156),
.CON(n_216),
.SN(n_216)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_221),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_152),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_187),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_170),
.B1(n_163),
.B2(n_148),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_177),
.A2(n_168),
.B(n_151),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_202),
.B(n_206),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_203),
.C(n_180),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_230),
.A2(n_239),
.B1(n_245),
.B2(n_208),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_244),
.Y(n_249)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_228),
.Y(n_260)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_207),
.B(n_190),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_238),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_178),
.B1(n_181),
.B2(n_188),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_242),
.C(n_219),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_192),
.C(n_189),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_184),
.B1(n_199),
.B2(n_205),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_246),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_194),
.B(n_203),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_219),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_254),
.B1(n_258),
.B2(n_261),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_248),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_230),
.A2(n_225),
.B1(n_216),
.B2(n_228),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_255),
.B(n_260),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_225),
.B1(n_226),
.B2(n_224),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_218),
.B1(n_227),
.B2(n_216),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_212),
.CI(n_10),
.CON(n_263),
.SN(n_263)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_242),
.C(n_231),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_270),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_241),
.B1(n_240),
.B2(n_247),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_250),
.B1(n_254),
.B2(n_256),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_277),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_257),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_241),
.B1(n_234),
.B2(n_237),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_271),
.A2(n_250),
.B1(n_264),
.B2(n_259),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_244),
.C(n_236),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_273),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_10),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_14),
.Y(n_274)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_7),
.B(n_9),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_14),
.B(n_6),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_11),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

NOR2x1_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_260),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_272),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_5),
.C(n_6),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_287),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_277),
.B(n_263),
.CI(n_13),
.CON(n_287),
.SN(n_287)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_278),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_263),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_5),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_292),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_283),
.A2(n_268),
.B(n_278),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_282),
.B1(n_289),
.B2(n_279),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_270),
.B(n_5),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_287),
.B(n_6),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_296),
.B(n_282),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_285),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_301),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_295),
.C(n_293),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

OAI321xp33_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_307),
.A3(n_298),
.B1(n_304),
.B2(n_299),
.C(n_290),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_305),
.B(n_296),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_5),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_6),
.Y(n_313)
);


endmodule