module fake_ibex_58_n_1050 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1050);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1050;

wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_1031;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_375;
wire n_340;
wire n_317;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_798;
wire n_732;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_538;
wire n_464;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_1030;
wire n_791;
wire n_715;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_980;
wire n_849;
wire n_454;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_1038;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_801;
wire n_718;
wire n_918;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_554;
wire n_553;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_566;
wire n_484;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_1049;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_506;
wire n_444;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_397;
wire n_366;
wire n_283;
wire n_894;
wire n_803;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_951;
wire n_272;
wire n_881;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_195;
wire n_885;
wire n_588;
wire n_212;
wire n_513;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_874;
wire n_816;
wire n_890;
wire n_921;
wire n_912;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_56),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_49),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_71),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_14),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_156),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_57),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_66),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_68),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_8),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_145),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_126),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_38),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_25),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_120),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_11),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_45),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_50),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_155),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_87),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_26),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_147),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_86),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_137),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_63),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_64),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_48),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_153),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_76),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_115),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_144),
.B(n_178),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_34),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_70),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_93),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_43),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_84),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_91),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_160),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_16),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_3),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_138),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_96),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_13),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_5),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_170),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_21),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_44),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_80),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_81),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_161),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_47),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_158),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_19),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_100),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_118),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_40),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_117),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_143),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_72),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_83),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_101),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_109),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_141),
.B(n_51),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_116),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_25),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_104),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_172),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_121),
.B(n_79),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_176),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_103),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_181),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_75),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_44),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_67),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_135),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_132),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_127),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_125),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_162),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_55),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_136),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_124),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_89),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_26),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_11),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_183),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_110),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_129),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_151),
.Y(n_285)
);

INVx4_ASAP7_75t_R g286 ( 
.A(n_90),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_185),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_32),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_5),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_105),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_31),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_3),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_165),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_65),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_54),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_46),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_97),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_16),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_21),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_82),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_95),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_22),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_2),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_150),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_99),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_2),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_34),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_139),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_19),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_106),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_149),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_69),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_154),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_60),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_20),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_38),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_111),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_92),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_36),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_166),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_27),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_123),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_74),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_112),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_78),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_30),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_152),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_58),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_8),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_20),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_1),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_39),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_113),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_289),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_232),
.Y(n_335)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_192),
.A2(n_200),
.B1(n_332),
.B2(n_236),
.Y(n_339)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_203),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_189),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_197),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_203),
.Y(n_344)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_215),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_215),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_215),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_197),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_192),
.A2(n_200),
.B1(n_236),
.B2(n_198),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_198),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_350)
);

AND2x2_ASAP7_75t_SL g351 ( 
.A(n_194),
.B(n_4),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_215),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_321),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_201),
.B(n_6),
.Y(n_354)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_218),
.B(n_52),
.Y(n_355)
);

AND2x6_ASAP7_75t_L g356 ( 
.A(n_218),
.B(n_182),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_225),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_201),
.B(n_7),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_280),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_313),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_280),
.B(n_7),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_229),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_239),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_256),
.B(n_9),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_239),
.B(n_9),
.Y(n_365)
);

BUFx12f_ASAP7_75t_L g366 ( 
.A(n_321),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_243),
.A2(n_10),
.B1(n_12),
.B2(n_15),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_243),
.A2(n_10),
.B1(n_12),
.B2(n_15),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_261),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_261),
.B(n_17),
.Y(n_370)
);

BUFx8_ASAP7_75t_SL g371 ( 
.A(n_255),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_213),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_242),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_229),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_229),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_228),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_202),
.B(n_17),
.Y(n_377)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_229),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_212),
.B(n_18),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_187),
.B(n_18),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g381 ( 
.A1(n_207),
.A2(n_102),
.B(n_179),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_231),
.B(n_180),
.Y(n_383)
);

BUFx12f_ASAP7_75t_L g384 ( 
.A(n_233),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_237),
.Y(n_385)
);

AND2x6_ASAP7_75t_L g386 ( 
.A(n_231),
.B(n_177),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_242),
.Y(n_387)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_237),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_255),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_242),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_307),
.Y(n_392)
);

OAI21x1_ASAP7_75t_L g393 ( 
.A1(n_230),
.A2(n_98),
.B(n_174),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g394 ( 
.A1(n_230),
.A2(n_94),
.B(n_171),
.Y(n_394)
);

AOI22x1_ASAP7_75t_SL g395 ( 
.A1(n_266),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_266),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_237),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_188),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_204),
.B(n_28),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_305),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_305),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_272),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_249),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_191),
.Y(n_404)
);

BUFx12f_ASAP7_75t_L g405 ( 
.A(n_234),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_305),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_272),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_407)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_305),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_195),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_196),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_300),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_300),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_206),
.B(n_33),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_238),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_281),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_245),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_205),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_288),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_235),
.B(n_35),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_209),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_291),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_241),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_210),
.Y(n_423)
);

OAI22x1_ASAP7_75t_R g424 ( 
.A1(n_292),
.A2(n_319),
.B1(n_302),
.B2(n_331),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_211),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_252),
.B(n_269),
.Y(n_426)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_254),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_254),
.B(n_37),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_216),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_220),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_299),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_221),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_223),
.Y(n_433)
);

BUFx12f_ASAP7_75t_L g434 ( 
.A(n_303),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_282),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_306),
.Y(n_436)
);

OA21x2_ASAP7_75t_L g437 ( 
.A1(n_262),
.A2(n_278),
.B(n_271),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_271),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_309),
.B(n_42),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_437),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_360),
.B(n_193),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_437),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_398),
.B(n_278),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_365),
.Y(n_444)
);

NAND3xp33_ASAP7_75t_L g445 ( 
.A(n_377),
.B(n_329),
.C(n_315),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_360),
.B(n_335),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_398),
.B(n_308),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_382),
.B(n_227),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_404),
.B(n_308),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_355),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_438),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_404),
.B(n_328),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_L g453 ( 
.A(n_355),
.B(n_186),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_438),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_370),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_354),
.Y(n_456)
);

AO22x2_ASAP7_75t_L g457 ( 
.A1(n_395),
.A2(n_316),
.B1(n_326),
.B2(n_330),
.Y(n_457)
);

AO21x2_ASAP7_75t_L g458 ( 
.A1(n_393),
.A2(n_259),
.B(n_226),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_354),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_358),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_376),
.B(n_415),
.Y(n_461)
);

NOR2x1p5_ASAP7_75t_L g462 ( 
.A(n_366),
.B(n_199),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_438),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_341),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_361),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_361),
.Y(n_466)
);

NOR2x1p5_ASAP7_75t_L g467 ( 
.A(n_384),
.B(n_199),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_341),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_428),
.B(n_248),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_409),
.B(n_250),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_344),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_334),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_344),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_346),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_334),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_338),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_347),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_418),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_439),
.B(n_253),
.Y(n_479)
);

AND3x2_ASAP7_75t_L g480 ( 
.A(n_353),
.B(n_219),
.C(n_222),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_410),
.B(n_257),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_338),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_419),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_435),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_439),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_410),
.B(n_258),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_435),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_337),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_379),
.B(n_320),
.C(n_327),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_359),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_372),
.B(n_320),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_422),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_422),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_336),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_352),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_417),
.B(n_420),
.Y(n_496)
);

NOR2x1p5_ASAP7_75t_L g497 ( 
.A(n_405),
.B(n_322),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_371),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_340),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_362),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_411),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_362),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_420),
.B(n_265),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_362),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_374),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_356),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_423),
.B(n_324),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_423),
.B(n_325),
.Y(n_508)
);

OR2x6_ASAP7_75t_L g509 ( 
.A(n_350),
.B(n_224),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_343),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_425),
.B(n_267),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_414),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_374),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_375),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_425),
.B(n_273),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_421),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_429),
.B(n_274),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_343),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_383),
.Y(n_519)
);

INVx8_ASAP7_75t_L g520 ( 
.A(n_383),
.Y(n_520)
);

AND3x2_ASAP7_75t_L g521 ( 
.A(n_436),
.B(n_297),
.C(n_311),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_429),
.B(n_277),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_348),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_383),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_430),
.B(n_325),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_357),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_430),
.B(n_284),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_357),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_342),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_432),
.B(n_287),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_416),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_364),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_375),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_433),
.B(n_208),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_433),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_426),
.B(n_290),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_380),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_385),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_363),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_363),
.B(n_294),
.Y(n_540)
);

AOI21x1_ASAP7_75t_L g541 ( 
.A1(n_381),
.A2(n_301),
.B(n_310),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_369),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_391),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_385),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_396),
.B(n_264),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_391),
.B(n_214),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_434),
.B(n_286),
.Y(n_547)
);

NOR2x1_ASAP7_75t_L g548 ( 
.A(n_399),
.B(n_190),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_385),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_349),
.A2(n_298),
.B1(n_247),
.B2(n_295),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_392),
.B(n_217),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_413),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_397),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_552),
.B(n_383),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_441),
.B(n_446),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_535),
.B(n_386),
.Y(n_556)
);

NOR3xp33_ASAP7_75t_L g557 ( 
.A(n_550),
.B(n_389),
.C(n_367),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_446),
.B(n_389),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_536),
.B(n_386),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_L g560 ( 
.A(n_520),
.B(n_386),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_478),
.Y(n_561)
);

NOR3xp33_ASAP7_75t_L g562 ( 
.A(n_445),
.B(n_407),
.C(n_368),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_L g563 ( 
.A(n_516),
.B(n_416),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_448),
.B(n_351),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_450),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_461),
.Y(n_566)
);

NAND2x1p5_ASAP7_75t_L g567 ( 
.A(n_459),
.B(n_431),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_492),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_491),
.B(n_240),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_L g570 ( 
.A(n_520),
.B(n_244),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_507),
.B(n_246),
.Y(n_571)
);

NOR3xp33_ASAP7_75t_L g572 ( 
.A(n_489),
.B(n_412),
.C(n_402),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_490),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_516),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_508),
.B(n_251),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_525),
.B(n_260),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_534),
.B(n_263),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_493),
.B(n_268),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_493),
.B(n_270),
.Y(n_579)
);

INVx6_ASAP7_75t_L g580 ( 
.A(n_529),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_472),
.B(n_394),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_475),
.B(n_476),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_459),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_523),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_537),
.B(n_275),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_537),
.B(n_276),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_524),
.B(n_279),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_512),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_479),
.A2(n_283),
.B1(n_285),
.B2(n_293),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_529),
.B(n_339),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_546),
.B(n_296),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_551),
.B(n_304),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_551),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_483),
.B(n_312),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_506),
.B(n_314),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_501),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_460),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_506),
.B(n_317),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_547),
.B(n_485),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_523),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_460),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_498),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_532),
.B(n_318),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_547),
.Y(n_604)
);

AND2x2_ASAP7_75t_SL g605 ( 
.A(n_453),
.B(n_424),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_519),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_519),
.B(n_333),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_466),
.B(n_427),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_456),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_488),
.Y(n_610)
);

AND2x6_ASAP7_75t_SL g611 ( 
.A(n_509),
.B(n_424),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_465),
.B(n_394),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_548),
.B(n_444),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_455),
.B(n_408),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_479),
.A2(n_390),
.B1(n_373),
.B2(n_403),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_547),
.B(n_387),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_496),
.B(n_388),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_494),
.Y(n_618)
);

INVxp67_ASAP7_75t_SL g619 ( 
.A(n_440),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_482),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_496),
.B(n_388),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_480),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_527),
.B(n_469),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_480),
.B(n_378),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_527),
.B(n_345),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_531),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_481),
.B(n_345),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_503),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_510),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_499),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_503),
.B(n_511),
.Y(n_631)
);

BUFx5_ASAP7_75t_L g632 ( 
.A(n_527),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_469),
.B(n_511),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_515),
.B(n_53),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_517),
.B(n_406),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_518),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_522),
.B(n_406),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_SL g638 ( 
.A(n_509),
.B(n_401),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_470),
.B(n_400),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_609),
.B(n_462),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_628),
.B(n_470),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_631),
.B(n_486),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_593),
.B(n_555),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_554),
.A2(n_440),
.B(n_442),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_620),
.B(n_442),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_619),
.A2(n_581),
.B(n_612),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_574),
.B(n_545),
.Y(n_647)
);

O2A1O1Ixp33_ASAP7_75t_L g648 ( 
.A1(n_562),
.A2(n_572),
.B(n_564),
.C(n_633),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_588),
.B(n_545),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_561),
.B(n_509),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_584),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_558),
.A2(n_545),
.B1(n_457),
.B2(n_467),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_563),
.B(n_497),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_560),
.A2(n_458),
.B(n_447),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_556),
.A2(n_458),
.B(n_447),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_556),
.A2(n_452),
.B(n_443),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_599),
.B(n_521),
.Y(n_657)
);

A2O1A1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_582),
.A2(n_540),
.B(n_526),
.C(n_528),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_633),
.B(n_530),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_559),
.A2(n_449),
.B(n_443),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_583),
.Y(n_661)
);

INVx1_ASAP7_75t_SL g662 ( 
.A(n_580),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_559),
.A2(n_449),
.B(n_452),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_582),
.A2(n_539),
.B(n_543),
.C(n_542),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_566),
.B(n_457),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_600),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_610),
.B(n_521),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_597),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_567),
.B(n_541),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_613),
.B(n_457),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_618),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_601),
.Y(n_672)
);

AO21x1_ASAP7_75t_L g673 ( 
.A1(n_634),
.A2(n_451),
.B(n_454),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_629),
.A2(n_484),
.B(n_487),
.C(n_454),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_567),
.B(n_451),
.Y(n_675)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_636),
.A2(n_463),
.B(n_397),
.C(n_553),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_580),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_622),
.B(n_463),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_580),
.B(n_590),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_557),
.A2(n_549),
.B1(n_544),
.B2(n_538),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_630),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_569),
.B(n_59),
.Y(n_682)
);

NOR2xp67_ASAP7_75t_L g683 ( 
.A(n_602),
.B(n_61),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_616),
.B(n_62),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_565),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_596),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_565),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_604),
.B(n_585),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_632),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_623),
.A2(n_533),
.B1(n_464),
.B2(n_514),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_605),
.B(n_73),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_571),
.A2(n_477),
.B(n_513),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_568),
.B(n_77),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_568),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_575),
.A2(n_474),
.B(n_505),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_576),
.A2(n_474),
.B(n_504),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_611),
.Y(n_697)
);

INVx5_ASAP7_75t_L g698 ( 
.A(n_606),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_608),
.A2(n_577),
.B(n_614),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_586),
.B(n_85),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_603),
.B(n_88),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_594),
.B(n_107),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_591),
.B(n_592),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_589),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_638),
.B(n_108),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_635),
.A2(n_473),
.B1(n_502),
.B2(n_500),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_578),
.B(n_114),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_579),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_573),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_570),
.A2(n_471),
.B1(n_468),
.B2(n_495),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_626),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_626),
.Y(n_712)
);

AOI21x1_ASAP7_75t_L g713 ( 
.A1(n_654),
.A2(n_673),
.B(n_655),
.Y(n_713)
);

NAND2x1_ASAP7_75t_L g714 ( 
.A(n_693),
.B(n_639),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_697),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_644),
.A2(n_637),
.B(n_639),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_L g717 ( 
.A1(n_646),
.A2(n_615),
.B(n_625),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_643),
.B(n_624),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_703),
.A2(n_617),
.B(n_621),
.C(n_627),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_645),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_645),
.A2(n_587),
.B(n_598),
.Y(n_721)
);

AOI21x1_ASAP7_75t_L g722 ( 
.A1(n_682),
.A2(n_607),
.B(n_595),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_647),
.B(n_133),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_669),
.A2(n_134),
.B(n_140),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_658),
.A2(n_664),
.B1(n_642),
.B2(n_684),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_698),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_686),
.B(n_142),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_641),
.B(n_148),
.Y(n_728)
);

NOR2x1_ASAP7_75t_SL g729 ( 
.A(n_689),
.B(n_698),
.Y(n_729)
);

OAI22x1_ASAP7_75t_L g730 ( 
.A1(n_652),
.A2(n_159),
.B1(n_163),
.B2(n_164),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_649),
.B(n_168),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_656),
.A2(n_175),
.B(n_659),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_660),
.A2(n_663),
.B(n_699),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_684),
.A2(n_708),
.B1(n_704),
.B2(n_693),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_698),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_650),
.A2(n_665),
.B1(n_688),
.B2(n_657),
.Y(n_736)
);

AOI21xp33_ASAP7_75t_L g737 ( 
.A1(n_667),
.A2(n_675),
.B(n_640),
.Y(n_737)
);

O2A1O1Ixp5_ASAP7_75t_L g738 ( 
.A1(n_700),
.A2(n_702),
.B(n_701),
.C(n_707),
.Y(n_738)
);

O2A1O1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_670),
.A2(n_672),
.B(n_661),
.C(n_668),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_709),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_689),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_662),
.B(n_640),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_662),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_692),
.A2(n_696),
.B(n_695),
.Y(n_744)
);

AO31x2_ASAP7_75t_L g745 ( 
.A1(n_676),
.A2(n_674),
.A3(n_690),
.B(n_706),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_657),
.B(n_679),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_680),
.B(n_706),
.C(n_690),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_694),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_677),
.B(n_681),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_691),
.B(n_653),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_671),
.A2(n_651),
.B(n_666),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_653),
.B(n_694),
.Y(n_752)
);

NAND2x1p5_ASAP7_75t_L g753 ( 
.A(n_685),
.B(n_687),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_711),
.B(n_683),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_711),
.B(n_712),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_678),
.B(n_705),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_687),
.B(n_710),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_686),
.Y(n_758)
);

NAND2x1p5_ASAP7_75t_L g759 ( 
.A(n_698),
.B(n_662),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_643),
.B(n_648),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_643),
.B(n_648),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_644),
.A2(n_646),
.B(n_669),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_709),
.Y(n_763)
);

OAI21xp5_ASAP7_75t_L g764 ( 
.A1(n_644),
.A2(n_646),
.B(n_669),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_709),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_645),
.Y(n_766)
);

OAI21xp5_ASAP7_75t_L g767 ( 
.A1(n_644),
.A2(n_646),
.B(n_669),
.Y(n_767)
);

BUFx2_ASAP7_75t_SL g768 ( 
.A(n_662),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_643),
.B(n_389),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_686),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_644),
.A2(n_646),
.B(n_669),
.Y(n_771)
);

AOI21xp33_ASAP7_75t_L g772 ( 
.A1(n_643),
.A2(n_649),
.B(n_564),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_643),
.B(n_648),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_643),
.B(n_648),
.C(n_558),
.Y(n_774)
);

BUFx4_ASAP7_75t_SL g775 ( 
.A(n_697),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_643),
.B(n_648),
.Y(n_776)
);

NAND2x1p5_ASAP7_75t_L g777 ( 
.A(n_698),
.B(n_662),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_645),
.Y(n_778)
);

INVxp67_ASAP7_75t_SL g779 ( 
.A(n_645),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_SL g780 ( 
.A(n_652),
.B(n_501),
.C(n_411),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_643),
.B(n_648),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_643),
.B(n_648),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_709),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_643),
.B(n_648),
.Y(n_784)
);

AO31x2_ASAP7_75t_L g785 ( 
.A1(n_673),
.A2(n_669),
.A3(n_654),
.B(n_655),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_686),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_643),
.B(n_648),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_643),
.B(n_648),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_644),
.A2(n_646),
.B(n_669),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_698),
.Y(n_790)
);

NAND2xp33_ASAP7_75t_SL g791 ( 
.A(n_643),
.B(n_198),
.Y(n_791)
);

AND3x4_ASAP7_75t_L g792 ( 
.A(n_657),
.B(n_557),
.C(n_572),
.Y(n_792)
);

OAI22x1_ASAP7_75t_L g793 ( 
.A1(n_652),
.A2(n_411),
.B1(n_367),
.B2(n_402),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_643),
.B(n_648),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_709),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_697),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_709),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_643),
.B(n_574),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_644),
.A2(n_646),
.B(n_669),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_643),
.B(n_648),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_647),
.A2(n_557),
.B1(n_562),
.B2(n_572),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_644),
.A2(n_646),
.B(n_669),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_720),
.A2(n_779),
.B(n_738),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_791),
.Y(n_804)
);

AOI221xp5_ASAP7_75t_L g805 ( 
.A1(n_772),
.A2(n_801),
.B1(n_793),
.B2(n_774),
.C(n_798),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_769),
.B(n_718),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_770),
.B(n_758),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_775),
.Y(n_808)
);

AOI22x1_ASAP7_75t_L g809 ( 
.A1(n_730),
.A2(n_733),
.B1(n_732),
.B2(n_744),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_759),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_715),
.Y(n_811)
);

AO21x2_ASAP7_75t_L g812 ( 
.A1(n_762),
.A2(n_802),
.B(n_767),
.Y(n_812)
);

CKINVDCx11_ASAP7_75t_R g813 ( 
.A(n_786),
.Y(n_813)
);

INVx3_ASAP7_75t_SL g814 ( 
.A(n_735),
.Y(n_814)
);

AO21x2_ASAP7_75t_L g815 ( 
.A1(n_802),
.A2(n_764),
.B(n_799),
.Y(n_815)
);

BUFx2_ASAP7_75t_SL g816 ( 
.A(n_735),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_750),
.B(n_736),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_740),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_760),
.B(n_761),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_734),
.B(n_768),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_743),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_759),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_790),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_763),
.Y(n_824)
);

OAI21x1_ASAP7_75t_SL g825 ( 
.A1(n_729),
.A2(n_724),
.B(n_739),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_765),
.Y(n_826)
);

OA21x2_ASAP7_75t_L g827 ( 
.A1(n_764),
.A2(n_771),
.B(n_789),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_SL g828 ( 
.A(n_796),
.B(n_790),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_726),
.Y(n_829)
);

OAI21x1_ASAP7_75t_SL g830 ( 
.A1(n_724),
.A2(n_800),
.B(n_794),
.Y(n_830)
);

INVx8_ASAP7_75t_L g831 ( 
.A(n_726),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_716),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_783),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_777),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_773),
.B(n_784),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_776),
.B(n_788),
.Y(n_836)
);

BUFx6f_ASAP7_75t_SL g837 ( 
.A(n_795),
.Y(n_837)
);

CKINVDCx6p67_ASAP7_75t_R g838 ( 
.A(n_742),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_781),
.A2(n_782),
.B(n_787),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_777),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_746),
.B(n_792),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_797),
.B(n_749),
.Y(n_842)
);

OAI21x1_ASAP7_75t_SL g843 ( 
.A1(n_725),
.A2(n_751),
.B(n_717),
.Y(n_843)
);

BUFx4f_ASAP7_75t_SL g844 ( 
.A(n_748),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_725),
.A2(n_747),
.B(n_717),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_780),
.A2(n_737),
.B1(n_731),
.B2(n_756),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_755),
.B(n_752),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_727),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_748),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_723),
.A2(n_754),
.B1(n_757),
.B2(n_714),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_719),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_721),
.B(n_728),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_722),
.Y(n_853)
);

BUFx4f_ASAP7_75t_L g854 ( 
.A(n_753),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_741),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_785),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_745),
.Y(n_857)
);

AO21x2_ASAP7_75t_L g858 ( 
.A1(n_713),
.A2(n_764),
.B(n_762),
.Y(n_858)
);

AND2x6_ASAP7_75t_L g859 ( 
.A(n_766),
.B(n_778),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_798),
.B(n_574),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_766),
.B(n_778),
.Y(n_861)
);

NAND2x1p5_ASAP7_75t_L g862 ( 
.A(n_735),
.B(n_790),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_766),
.B(n_778),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_720),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_791),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_766),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_772),
.B(n_769),
.Y(n_867)
);

AO21x2_ASAP7_75t_L g868 ( 
.A1(n_713),
.A2(n_764),
.B(n_762),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_740),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_798),
.B(n_769),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_740),
.Y(n_871)
);

OAI21x1_ASAP7_75t_SL g872 ( 
.A1(n_734),
.A2(n_729),
.B(n_724),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_740),
.Y(n_873)
);

OR2x6_ASAP7_75t_L g874 ( 
.A(n_734),
.B(n_768),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_806),
.B(n_870),
.Y(n_875)
);

INVxp33_ASAP7_75t_L g876 ( 
.A(n_813),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_813),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_832),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_859),
.Y(n_879)
);

NAND2x1_ASAP7_75t_L g880 ( 
.A(n_825),
.B(n_872),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_814),
.Y(n_881)
);

CKINVDCx11_ASAP7_75t_R g882 ( 
.A(n_814),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_841),
.B(n_806),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_841),
.A2(n_805),
.B1(n_867),
.B2(n_817),
.Y(n_884)
);

BUFx10_ASAP7_75t_L g885 ( 
.A(n_808),
.Y(n_885)
);

INVx6_ASAP7_75t_L g886 ( 
.A(n_831),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_864),
.Y(n_887)
);

AO21x2_ASAP7_75t_L g888 ( 
.A1(n_830),
.A2(n_843),
.B(n_845),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_864),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_867),
.A2(n_819),
.B1(n_836),
.B2(n_835),
.Y(n_890)
);

OAI22xp33_ASAP7_75t_L g891 ( 
.A1(n_804),
.A2(n_865),
.B1(n_874),
.B2(n_820),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_820),
.A2(n_874),
.B1(n_866),
.B2(n_846),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_859),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_861),
.A2(n_863),
.B1(n_846),
.B2(n_866),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_861),
.B(n_863),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_861),
.A2(n_863),
.B1(n_860),
.B2(n_839),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_821),
.B(n_820),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_831),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_858),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_807),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_818),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_859),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_831),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_842),
.B(n_824),
.Y(n_904)
);

AOI211xp5_ASAP7_75t_L g905 ( 
.A1(n_848),
.A2(n_828),
.B(n_847),
.C(n_833),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_826),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_869),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_871),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_873),
.B(n_855),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_853),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_816),
.B(n_838),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_837),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_874),
.A2(n_850),
.B1(n_837),
.B2(n_823),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_854),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_854),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_910),
.Y(n_916)
);

NOR2xp67_ASAP7_75t_L g917 ( 
.A(n_913),
.B(n_840),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_893),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_883),
.A2(n_851),
.B1(n_850),
.B2(n_812),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_879),
.B(n_856),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_887),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_893),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_884),
.A2(n_815),
.B1(n_812),
.B2(n_823),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_888),
.B(n_827),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_902),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_888),
.B(n_827),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_875),
.A2(n_890),
.B1(n_892),
.B2(n_896),
.Y(n_927)
);

INVxp67_ASAP7_75t_SL g928 ( 
.A(n_887),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_888),
.B(n_827),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_889),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_889),
.B(n_897),
.Y(n_931)
);

NOR2x1_ASAP7_75t_L g932 ( 
.A(n_891),
.B(n_822),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_878),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_896),
.A2(n_856),
.B1(n_857),
.B2(n_809),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_901),
.B(n_906),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_933),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_916),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_918),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_927),
.B(n_901),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_921),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_927),
.A2(n_895),
.B1(n_876),
.B2(n_897),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_932),
.B(n_879),
.Y(n_942)
);

NOR3xp33_ASAP7_75t_L g943 ( 
.A(n_932),
.B(n_905),
.C(n_911),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_920),
.B(n_899),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_924),
.B(n_856),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_924),
.B(n_868),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_924),
.B(n_868),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_931),
.B(n_921),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_946),
.B(n_947),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_948),
.B(n_931),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_937),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_936),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_940),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_946),
.B(n_926),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_947),
.B(n_926),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_948),
.B(n_931),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_944),
.B(n_926),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_945),
.B(n_929),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_939),
.B(n_930),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_938),
.B(n_928),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_938),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_960),
.B(n_879),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_954),
.B(n_919),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_954),
.B(n_919),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_949),
.B(n_950),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_950),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_956),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_949),
.B(n_945),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_956),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_951),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_955),
.B(n_929),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_952),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_955),
.B(n_929),
.Y(n_973)
);

NAND2xp33_ASAP7_75t_L g974 ( 
.A(n_960),
.B(n_943),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_957),
.B(n_944),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_953),
.Y(n_976)
);

OR2x2_ASAP7_75t_SL g977 ( 
.A(n_961),
.B(n_912),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_959),
.B(n_923),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_L g979 ( 
.A(n_974),
.B(n_978),
.C(n_882),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_972),
.Y(n_980)
);

NOR2x1_ASAP7_75t_L g981 ( 
.A(n_974),
.B(n_917),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_966),
.B(n_953),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_968),
.B(n_958),
.Y(n_983)
);

OAI32xp33_ASAP7_75t_L g984 ( 
.A1(n_965),
.A2(n_942),
.A3(n_881),
.B1(n_922),
.B2(n_925),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_976),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_976),
.B(n_957),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_970),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_965),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_967),
.Y(n_989)
);

OAI22xp33_ASAP7_75t_L g990 ( 
.A1(n_962),
.A2(n_942),
.B1(n_917),
.B2(n_918),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_969),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_963),
.A2(n_957),
.B1(n_941),
.B2(n_958),
.Y(n_992)
);

OAI321xp33_ASAP7_75t_L g993 ( 
.A1(n_992),
.A2(n_964),
.A3(n_962),
.B1(n_942),
.B2(n_923),
.C(n_977),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_980),
.Y(n_994)
);

AO21x1_ASAP7_75t_L g995 ( 
.A1(n_979),
.A2(n_977),
.B(n_962),
.Y(n_995)
);

NAND2x1_ASAP7_75t_L g996 ( 
.A(n_986),
.B(n_975),
.Y(n_996)
);

AOI211x1_ASAP7_75t_L g997 ( 
.A1(n_984),
.A2(n_968),
.B(n_973),
.C(n_971),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_SL g998 ( 
.A1(n_981),
.A2(n_975),
.B(n_894),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_988),
.B(n_971),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_982),
.Y(n_1000)
);

NAND3xp33_ASAP7_75t_L g1001 ( 
.A(n_987),
.B(n_877),
.C(n_907),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_997),
.A2(n_986),
.B1(n_985),
.B2(n_982),
.Y(n_1002)
);

AOI21xp33_ASAP7_75t_SL g1003 ( 
.A1(n_1001),
.A2(n_990),
.B(n_987),
.Y(n_1003)
);

AND4x1_ASAP7_75t_L g1004 ( 
.A(n_1001),
.B(n_885),
.C(n_989),
.D(n_991),
.Y(n_1004)
);

OAI211xp5_ASAP7_75t_L g1005 ( 
.A1(n_998),
.A2(n_894),
.B(n_934),
.C(n_900),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_1000),
.Y(n_1006)
);

AOI221x1_ASAP7_75t_L g1007 ( 
.A1(n_995),
.A2(n_907),
.B1(n_908),
.B2(n_906),
.C(n_975),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_994),
.Y(n_1008)
);

OAI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_996),
.A2(n_973),
.B(n_983),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_999),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_1005),
.A2(n_993),
.B1(n_957),
.B2(n_972),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1006),
.Y(n_1012)
);

NAND4xp25_ASAP7_75t_L g1013 ( 
.A(n_1007),
.B(n_903),
.C(n_898),
.D(n_914),
.Y(n_1013)
);

NAND2xp67_ASAP7_75t_SL g1014 ( 
.A(n_1003),
.B(n_885),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_1002),
.A2(n_903),
.B(n_898),
.C(n_904),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_1008),
.Y(n_1016)
);

NAND2xp67_ASAP7_75t_SL g1017 ( 
.A(n_1004),
.B(n_885),
.Y(n_1017)
);

NOR2x1_ASAP7_75t_SL g1018 ( 
.A(n_1017),
.B(n_898),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_SL g1019 ( 
.A1(n_1016),
.A2(n_1010),
.B1(n_885),
.B2(n_1009),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_L g1020 ( 
.A(n_1015),
.B(n_811),
.C(n_1010),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_1012),
.A2(n_811),
.B(n_880),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_1011),
.B(n_951),
.Y(n_1022)
);

NAND4xp75_ASAP7_75t_L g1023 ( 
.A(n_1014),
.B(n_829),
.C(n_908),
.D(n_803),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1020),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1022),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1021),
.B(n_1013),
.Y(n_1026)
);

NAND4xp75_ASAP7_75t_L g1027 ( 
.A(n_1018),
.B(n_909),
.C(n_886),
.D(n_849),
.Y(n_1027)
);

NOR3xp33_ASAP7_75t_L g1028 ( 
.A(n_1023),
.B(n_840),
.C(n_810),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_1019),
.B(n_886),
.Y(n_1029)
);

NOR3xp33_ASAP7_75t_L g1030 ( 
.A(n_1023),
.B(n_834),
.C(n_915),
.Y(n_1030)
);

NOR2x1_ASAP7_75t_L g1031 ( 
.A(n_1024),
.B(n_903),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1026),
.Y(n_1032)
);

NAND2x1p5_ASAP7_75t_SL g1033 ( 
.A(n_1027),
.B(n_1029),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1025),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1030),
.Y(n_1035)
);

OA21x2_ASAP7_75t_L g1036 ( 
.A1(n_1032),
.A2(n_1028),
.B(n_852),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_1031),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_1037),
.Y(n_1038)
);

XNOR2xp5_ASAP7_75t_L g1039 ( 
.A(n_1036),
.B(n_1033),
.Y(n_1039)
);

INVxp67_ASAP7_75t_SL g1040 ( 
.A(n_1038),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_1039),
.B(n_1032),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_1040),
.A2(n_1041),
.B(n_1034),
.Y(n_1042)
);

AO22x2_ASAP7_75t_L g1043 ( 
.A1(n_1040),
.A2(n_1035),
.B1(n_1036),
.B2(n_915),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1043),
.Y(n_1044)
);

AOI21x1_ASAP7_75t_L g1045 ( 
.A1(n_1042),
.A2(n_935),
.B(n_909),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1043),
.A2(n_886),
.B1(n_914),
.B2(n_915),
.Y(n_1046)
);

AO221x2_ASAP7_75t_L g1047 ( 
.A1(n_1044),
.A2(n_886),
.B1(n_914),
.B2(n_844),
.C(n_935),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_1047),
.A2(n_1046),
.B(n_1045),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_1048),
.B(n_862),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_1049),
.A2(n_822),
.B1(n_844),
.B2(n_862),
.Y(n_1050)
);


endmodule