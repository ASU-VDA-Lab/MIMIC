module fake_jpeg_24890_n_265 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_37),
.B(n_42),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_43),
.B(n_44),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_0),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_17),
.B1(n_33),
.B2(n_32),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_51),
.A2(n_56),
.B1(n_58),
.B2(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_59),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_48),
.B1(n_41),
.B2(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

OA22x2_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_22),
.B1(n_34),
.B2(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_61),
.Y(n_99)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_69),
.Y(n_109)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_25),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_74),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_65),
.Y(n_107)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_28),
.B1(n_26),
.B2(n_32),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_17),
.B1(n_20),
.B2(n_33),
.Y(n_70)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_73),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_19),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_14),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_43),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_80),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_29),
.B1(n_20),
.B2(n_21),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_117)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_110)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_29),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_86),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_42),
.B(n_1),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_21),
.B1(n_18),
.B2(n_23),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_88),
.A2(n_71),
.B1(n_50),
.B2(n_6),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_34),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_35),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_35),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_116),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_52),
.B(n_18),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_54),
.C(n_56),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx6_ASAP7_75t_SL g112 ( 
.A(n_52),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_113),
.Y(n_119)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_1),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_78),
.B1(n_69),
.B2(n_66),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_58),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_120),
.B(n_121),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_53),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_123),
.B(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_92),
.B(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_130),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_84),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_131),
.B(n_134),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_72),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_141),
.B1(n_113),
.B2(n_11),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_63),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_136),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_83),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_106),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_142),
.B1(n_148),
.B2(n_102),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_71),
.B1(n_50),
.B2(n_85),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_143),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_114),
.A2(n_5),
.B(n_7),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_144),
.A2(n_147),
.B(n_108),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_5),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_145),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

CKINVDCx10_ASAP7_75t_R g154 ( 
.A(n_146),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_8),
.B(n_9),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_98),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_149),
.B(n_158),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_172),
.B(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_156),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_144),
.Y(n_178)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_106),
.B1(n_111),
.B2(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_162),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_106),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_164),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_90),
.Y(n_164)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_169),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_111),
.B1(n_100),
.B2(n_95),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_107),
.Y(n_171)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

NOR2x1p5_ASAP7_75t_SL g172 ( 
.A(n_118),
.B(n_100),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_94),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_135),
.B(n_140),
.C(n_127),
.Y(n_182)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_129),
.C(n_125),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_186),
.C(n_187),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_180),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_176),
.B1(n_164),
.B2(n_149),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_184),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_153),
.A2(n_127),
.B(n_120),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_195),
.B(n_162),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_142),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_124),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_128),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_171),
.Y(n_201)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_194),
.Y(n_202)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

AND2x4_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_201),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_154),
.Y(n_200)
);

AO21x1_ASAP7_75t_L g225 ( 
.A1(n_200),
.A2(n_210),
.B(n_214),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_163),
.C(n_158),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_180),
.C(n_195),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_209),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_151),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_208),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_212),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_152),
.B1(n_170),
.B2(n_159),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_216),
.C(n_218),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_157),
.C(n_188),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_186),
.C(n_150),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_178),
.C(n_166),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_227),
.C(n_228),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_203),
.B(n_187),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_200),
.C(n_228),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_225),
.A2(n_205),
.B(n_212),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_181),
.C(n_160),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_185),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_200),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_230),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_207),
.B1(n_211),
.B2(n_182),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_206),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_236),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_182),
.B1(n_201),
.B2(n_200),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_233),
.A2(n_238),
.B1(n_208),
.B2(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_239),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_217),
.A2(n_221),
.B1(n_179),
.B2(n_169),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_202),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_243),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_238),
.B(n_155),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_248),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_154),
.C(n_155),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_165),
.Y(n_251)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_251),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_165),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_252),
.B(n_254),
.Y(n_255)
);

OAI21x1_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_240),
.B(n_230),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_229),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_165),
.Y(n_254)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_256),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_248),
.C(n_234),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_257),
.A2(n_253),
.B1(n_246),
.B2(n_235),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_235),
.C(n_255),
.Y(n_262)
);

AOI21x1_ASAP7_75t_L g261 ( 
.A1(n_258),
.A2(n_247),
.B(n_249),
.Y(n_261)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_247),
.A3(n_156),
.B1(n_182),
.B2(n_100),
.C1(n_143),
.C2(n_12),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_260),
.Y(n_265)
);


endmodule