module fake_jpeg_22363_n_160 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_160);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_46),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_19),
.B1(n_25),
.B2(n_21),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_45),
.B1(n_25),
.B2(n_21),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_25),
.B1(n_21),
.B2(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_43),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_54),
.Y(n_70)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_55),
.A2(n_39),
.B1(n_24),
.B2(n_14),
.Y(n_80)
);

INVxp33_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_39),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_0),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_67),
.C(n_26),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_1),
.Y(n_72)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_39),
.Y(n_81)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_68),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_31),
.B(n_19),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_14),
.B(n_35),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_38),
.B(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_18),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_44),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_67),
.C(n_68),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_72),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_76),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_1),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_85),
.B(n_86),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_20),
.B1(n_46),
.B2(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_81),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_48),
.CON(n_76),
.SN(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_82),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_52),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_2),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_88),
.C(n_91),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_59),
.C(n_58),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_59),
.C(n_56),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_48),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_73),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_105),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_104),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_74),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_107),
.B(n_111),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_76),
.B(n_85),
.Y(n_107)
);

OA21x2_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_71),
.B(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_108),
.B(n_87),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_113),
.B(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_97),
.B1(n_95),
.B2(n_89),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_119),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_123),
.B(n_111),
.CI(n_106),
.CON(n_136),
.SN(n_136)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_127),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_97),
.B1(n_53),
.B2(n_65),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_115),
.C(n_114),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_79),
.B1(n_65),
.B2(n_28),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_128),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_28),
.B1(n_27),
.B2(n_23),
.Y(n_128)
);

BUFx24_ASAP7_75t_SL g129 ( 
.A(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_134),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_137),
.C(n_125),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_120),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_138),
.C(n_12),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_115),
.C(n_109),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_107),
.C(n_13),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_52),
.C(n_24),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_135),
.A2(n_124),
.B1(n_119),
.B2(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_119),
.B1(n_127),
.B2(n_27),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_144),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_132),
.B(n_133),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_145),
.B(n_17),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_23),
.B(n_17),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_143),
.B(n_14),
.CI(n_24),
.CON(n_146),
.SN(n_146)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_52),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_151),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_8),
.C1(n_142),
.C2(n_148),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_150),
.A2(n_141),
.B(n_6),
.C(n_5),
.Y(n_152)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_146),
.A3(n_147),
.B1(n_151),
.B2(n_149),
.C1(n_11),
.C2(n_13),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_146),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_3),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_155),
.A2(n_156),
.B(n_152),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_159),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);


endmodule