module fake_jpeg_30115_n_163 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_20),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx9p33_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_0),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_66),
.B(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_52),
.B(n_71),
.C(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_89),
.B(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_53),
.B(n_63),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_96),
.B(n_2),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_46),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_55),
.C(n_46),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_101),
.C(n_0),
.Y(n_115)
);

OR2x4_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_44),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_27),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_61),
.C(n_48),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_57),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_103),
.A2(n_64),
.B1(n_56),
.B2(n_58),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_64),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_5),
.C(n_8),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_112),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_96),
.B1(n_90),
.B2(n_97),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_126),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_121),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_124),
.B(n_8),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_122),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_2),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_3),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_125),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_28),
.B1(n_42),
.B2(n_39),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_137),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_136),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_143),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_43),
.B(n_30),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_29),
.B(n_37),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_141),
.B1(n_122),
.B2(n_120),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_11),
.B1(n_38),
.B2(n_15),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_14),
.C(n_16),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_139),
.B1(n_142),
.B2(n_137),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_124),
.B(n_23),
.C(n_25),
.D(n_32),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_151),
.C(n_19),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_127),
.C(n_114),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_139),
.B1(n_129),
.B2(n_131),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_153),
.B1(n_151),
.B2(n_146),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_155),
.A2(n_137),
.B(n_149),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_157),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_154),
.B1(n_147),
.B2(n_130),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_134),
.B(n_150),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_143),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_161),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_33),
.Y(n_163)
);


endmodule