module fake_jpeg_13345_n_369 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_369);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_369;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_58),
.Y(n_68)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_33),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_35),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_65),
.B(n_75),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_20),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_38),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_76),
.B(n_78),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_50),
.B1(n_61),
.B2(n_58),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_77),
.A2(n_41),
.B1(n_51),
.B2(n_47),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_25),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_43),
.A2(n_22),
.B1(n_37),
.B2(n_41),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_54),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_35),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_45),
.A2(n_22),
.B1(n_37),
.B2(n_41),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_35),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_29),
.B1(n_22),
.B2(n_37),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_44),
.A2(n_29),
.B1(n_35),
.B2(n_38),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_57),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_92),
.Y(n_135)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_130),
.B1(n_67),
.B2(n_80),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_18),
.B1(n_28),
.B2(n_40),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_122),
.B1(n_127),
.B2(n_41),
.Y(n_139)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_28),
.B(n_40),
.C(n_36),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_98),
.A2(n_99),
.B(n_107),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_36),
.B(n_42),
.C(n_24),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_71),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_110),
.Y(n_140)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_65),
.A2(n_55),
.B(n_23),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_23),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_126),
.C(n_85),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_82),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_118),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_84),
.B(n_56),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_128),
.C(n_60),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_121),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_18),
.B1(n_34),
.B2(n_27),
.Y(n_122)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_64),
.B(n_34),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g148 ( 
.A(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_70),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_69),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_64),
.B(n_70),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_69),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_85),
.B1(n_80),
.B2(n_73),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_91),
.A2(n_77),
.B1(n_87),
.B2(n_81),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_145),
.B1(n_155),
.B2(n_158),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_105),
.B1(n_126),
.B2(n_94),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_117),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_92),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_91),
.A2(n_73),
.B1(n_9),
.B2(n_10),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_95),
.A2(n_73),
.B1(n_9),
.B2(n_10),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_114),
.A2(n_8),
.B1(n_16),
.B2(n_14),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_107),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_171),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_135),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_172),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_120),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_136),
.A2(n_130),
.B1(n_111),
.B2(n_99),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_92),
.B1(n_130),
.B2(n_98),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_141),
.B1(n_139),
.B2(n_155),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_147),
.A2(n_97),
.B(n_129),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_147),
.Y(n_191)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_130),
.B1(n_113),
.B2(n_112),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_180),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_179),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_161),
.B(n_117),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_135),
.A2(n_93),
.B1(n_100),
.B2(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_101),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_189),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_131),
.B(n_119),
.CI(n_116),
.CON(n_184),
.SN(n_184)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_185),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_161),
.B(n_110),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_187),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_144),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_143),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_109),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_191),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_163),
.A2(n_141),
.B(n_102),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_193),
.A2(n_184),
.B(n_189),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_175),
.A2(n_145),
.B(n_149),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_194),
.A2(n_215),
.B(n_167),
.Y(n_232)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_148),
.Y(n_197)
);

A2O1A1O1Ixp25_ASAP7_75t_L g241 ( 
.A1(n_197),
.A2(n_186),
.B(n_151),
.C(n_187),
.D(n_156),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_183),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_210),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

AO21x2_ASAP7_75t_L g208 ( 
.A1(n_173),
.A2(n_159),
.B(n_153),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_218),
.B1(n_210),
.B2(n_214),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_213),
.B(n_133),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_149),
.B(n_151),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_180),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_218),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_132),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_169),
.C(n_168),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_222),
.B(n_224),
.C(n_250),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_162),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_220),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_225),
.B(n_240),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_239),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_228),
.A2(n_229),
.B1(n_212),
.B2(n_194),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_195),
.A2(n_165),
.B1(n_174),
.B2(n_173),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_206),
.A2(n_177),
.B1(n_172),
.B2(n_171),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_233),
.B1(n_236),
.B2(n_238),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_235),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_195),
.A2(n_184),
.B1(n_164),
.B2(n_181),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_200),
.A2(n_166),
.B1(n_176),
.B2(n_182),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_165),
.B1(n_178),
.B2(n_187),
.Y(n_238)
);

INVxp33_ASAP7_75t_SL g239 ( 
.A(n_196),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_241),
.B(n_247),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_143),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_208),
.B1(n_204),
.B2(n_199),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_191),
.A2(n_209),
.B(n_203),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_248),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_196),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_187),
.B(n_133),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_249),
.B(n_207),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_203),
.B(n_13),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_222),
.B(n_197),
.Y(n_255)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_255),
.B(n_275),
.C(n_268),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_227),
.A2(n_212),
.B1(n_201),
.B2(n_216),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_256),
.A2(n_259),
.B1(n_208),
.B2(n_214),
.Y(n_283)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_258),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_230),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_267),
.Y(n_291)
);

OAI32xp33_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_197),
.A3(n_202),
.B1(n_198),
.B2(n_207),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_263),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_245),
.Y(n_264)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_229),
.A2(n_202),
.B1(n_208),
.B2(n_205),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_236),
.B1(n_242),
.B2(n_238),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_198),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_266),
.B(n_270),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_202),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_271),
.Y(n_297)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_273),
.B(n_244),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_224),
.B(n_193),
.C(n_202),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_232),
.C(n_223),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_205),
.C(n_204),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_284),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_223),
.B1(n_242),
.B2(n_221),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_278),
.A2(n_292),
.B1(n_288),
.B2(n_261),
.Y(n_300)
);

AOI21xp33_ASAP7_75t_L g279 ( 
.A1(n_262),
.A2(n_248),
.B(n_250),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_279),
.A2(n_286),
.B(n_290),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_280),
.A2(n_282),
.B1(n_283),
.B2(n_146),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_235),
.C(n_233),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_294),
.C(n_257),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_259),
.A2(n_231),
.B1(n_208),
.B2(n_241),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_199),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_252),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_11),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_257),
.A2(n_261),
.B(n_251),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_208),
.B(n_217),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_295),
.Y(n_301)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_251),
.A2(n_214),
.B(n_132),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_269),
.A2(n_153),
.B1(n_146),
.B2(n_123),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_254),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_298),
.A2(n_297),
.B(n_292),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_300),
.A2(n_280),
.B1(n_297),
.B2(n_278),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_276),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_304),
.C(n_308),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_263),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_277),
.A2(n_296),
.B1(n_253),
.B2(n_264),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_306),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_296),
.A2(n_256),
.B1(n_271),
.B2(n_265),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_307),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_269),
.C(n_272),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_313),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_272),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_314),
.C(n_316),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_312),
.A2(n_106),
.B1(n_103),
.B2(n_9),
.Y(n_325)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_291),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_115),
.C(n_108),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_315),
.A2(n_17),
.B1(n_14),
.B2(n_12),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_282),
.B(n_115),
.C(n_108),
.Y(n_316)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_318),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_319),
.B(n_325),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_297),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_322),
.A2(n_302),
.B(n_308),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_16),
.C(n_14),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_329),
.C(n_314),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_328),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_8),
.C(n_11),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_298),
.A2(n_6),
.B(n_1),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_330),
.B(n_331),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_299),
.B(n_0),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_1),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_1),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_310),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_336),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_311),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_304),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_337),
.B(n_340),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_342),
.Y(n_350)
);

INVx11_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_301),
.C(n_316),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_343),
.B(n_324),
.C(n_328),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_332),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_321),
.Y(n_345)
);

AO21x1_ASAP7_75t_L g354 ( 
.A1(n_345),
.A2(n_334),
.B(n_318),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_348),
.Y(n_359)
);

BUFx24_ASAP7_75t_SL g347 ( 
.A(n_335),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_347),
.B(n_340),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_326),
.C(n_324),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_351),
.B(n_352),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_327),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_357),
.C(n_2),
.Y(n_364)
);

NOR4xp25_ASAP7_75t_L g355 ( 
.A(n_349),
.B(n_338),
.C(n_322),
.D(n_342),
.Y(n_355)
);

O2A1O1Ixp33_ASAP7_75t_SL g362 ( 
.A1(n_355),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_356),
.B(n_358),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_353),
.A2(n_345),
.B(n_350),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_338),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_360),
.A2(n_344),
.B(n_3),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_361),
.A2(n_362),
.B(n_364),
.Y(n_366)
);

AOI321xp33_ASAP7_75t_L g365 ( 
.A1(n_363),
.A2(n_359),
.A3(n_355),
.B1(n_5),
.B2(n_6),
.C(n_4),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_365),
.Y(n_367)
);

OAI321xp33_ASAP7_75t_L g368 ( 
.A1(n_367),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_366),
.C(n_360),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_368),
.B(n_2),
.Y(n_369)
);


endmodule