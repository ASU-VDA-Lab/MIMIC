module real_jpeg_2738_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_0),
.B(n_10),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_0),
.B(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_1),
.Y(n_18)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_1),
.B(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_1),
.B(n_24),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

AO21x2_ASAP7_75t_L g10 ( 
.A1(n_3),
.A2(n_11),
.B(n_12),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_11),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_28),
.Y(n_27)
);

NAND2x1_ASAP7_75t_SL g29 ( 
.A(n_5),
.B(n_28),
.Y(n_29)
);

NOR3xp33_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_21),
.C(n_31),
.Y(n_6)
);

OAI221xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_7)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_8),
.A2(n_15),
.B1(n_22),
.B2(n_30),
.Y(n_21)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_10),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_10),
.A2(n_19),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_25),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_14),
.Y(n_13)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_14),
.B(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_24),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);


endmodule