module fake_jpeg_22278_n_103 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_17),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_26),
.A2(n_29),
.B1(n_24),
.B2(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_19),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_7),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_30),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_17),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_8),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_48),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_65),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_27),
.B1(n_33),
.B2(n_14),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_61),
.B1(n_41),
.B2(n_16),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_22),
.B1(n_13),
.B2(n_18),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_59),
.B1(n_37),
.B2(n_46),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_32),
.C(n_25),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_16),
.B(n_10),
.Y(n_73)
);

AO22x2_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_32),
.B1(n_19),
.B2(n_18),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_13),
.B1(n_18),
.B2(n_12),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_16),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_74),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.Y(n_83)
);

AO21x1_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_37),
.B(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_75),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_10),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_11),
.C(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_76),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_56),
.B1(n_53),
.B2(n_64),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_68),
.B1(n_59),
.B2(n_73),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_67),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_81),
.B1(n_83),
.B2(n_82),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_86),
.C(n_90),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_88),
.B(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_90),
.B1(n_94),
.B2(n_93),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_98),
.A2(n_97),
.B(n_77),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_101),
.A3(n_87),
.B1(n_77),
.B2(n_52),
.C1(n_63),
.C2(n_54),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_87),
.B(n_57),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_61),
.Y(n_103)
);


endmodule