module fake_netlist_6_3557_n_1781 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1781);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1781;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_1),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_5),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_58),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_28),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_21),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_88),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_75),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_2),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_100),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_90),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_34),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_16),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_63),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_34),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_3),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_51),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_54),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_27),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_16),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_55),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_22),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_105),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_20),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_143),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_129),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_7),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_35),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_2),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_85),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_37),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_76),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_96),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_70),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_160),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_127),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_93),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_152),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_91),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_112),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_122),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_11),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_138),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_45),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_87),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_117),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_103),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_1),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_17),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_106),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_113),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_101),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_155),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_48),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_124),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_19),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_42),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_86),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_8),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_119),
.Y(n_234)
);

INVxp67_ASAP7_75t_SL g235 ( 
.A(n_14),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_89),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_116),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_12),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_60),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_110),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_136),
.Y(n_242)
);

BUFx8_ASAP7_75t_SL g243 ( 
.A(n_33),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_74),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_145),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_77),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_94),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_128),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_132),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_163),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_41),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_59),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_82),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_12),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_141),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_24),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_65),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_111),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_159),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_137),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_57),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_134),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_22),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_79),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_72),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_71),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_81),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_83),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_41),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_109),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_157),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_115),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_14),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_130),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_80),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_61),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_29),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_18),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_64),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_108),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_27),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_125),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_98),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_167),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_52),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_149),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_25),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_21),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_131),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_24),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_28),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_156),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_30),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_36),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_69),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_95),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_56),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_51),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_118),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_45),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_29),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_68),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_66),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_150),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_10),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_107),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_140),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_15),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_36),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_135),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_38),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_17),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_37),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_46),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_9),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_151),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_19),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_73),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_120),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_32),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_44),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_148),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_8),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_142),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_11),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_46),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_18),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_4),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_53),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_102),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_23),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_133),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_123),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_43),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_3),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_7),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_223),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_229),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_243),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_229),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_232),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_229),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_171),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_229),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_229),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_181),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_181),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_232),
.B(n_0),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_234),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_290),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_174),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_196),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_290),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_178),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_317),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_253),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_272),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_284),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_182),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_172),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_187),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_172),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_192),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_186),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_170),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_194),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_302),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_285),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_186),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_333),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_195),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_176),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_191),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_200),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_237),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_191),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_230),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_230),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_251),
.Y(n_380)
);

NOR2xp67_ASAP7_75t_L g381 ( 
.A(n_251),
.B(n_0),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_254),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_202),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_206),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_280),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_254),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_285),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_205),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_207),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_170),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_175),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_208),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_256),
.B(n_4),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_210),
.Y(n_394)
);

INVxp33_ASAP7_75t_SL g395 ( 
.A(n_168),
.Y(n_395)
);

INVxp33_ASAP7_75t_SL g396 ( 
.A(n_169),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_256),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_291),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_291),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_211),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_173),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_215),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_301),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_301),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_237),
.Y(n_405)
);

NOR2xp67_ASAP7_75t_L g406 ( 
.A(n_311),
.B(n_5),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_311),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_217),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_321),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_219),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_321),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_222),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_225),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_295),
.B(n_6),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_328),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_295),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_328),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_227),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_334),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_236),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_177),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_320),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_246),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_369),
.Y(n_424)
);

INVx6_ASAP7_75t_L g425 ( 
.A(n_348),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_337),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_349),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_387),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_246),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_338),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_389),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_340),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_395),
.B(n_396),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_340),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_342),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_342),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_357),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_344),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_343),
.B(n_261),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_344),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_358),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_408),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_348),
.B(n_179),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_345),
.B(n_179),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_345),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_351),
.B(n_224),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_376),
.B(n_320),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_390),
.B(n_224),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_413),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_359),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_325),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_R g453 ( 
.A(n_355),
.B(n_360),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_350),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_350),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_362),
.B(n_364),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_366),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_368),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_361),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_401),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_367),
.B(n_231),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_418),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_361),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_346),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_363),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_372),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_346),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_363),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_365),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_365),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_416),
.B(n_325),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_421),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_375),
.B(n_231),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_383),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_347),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_370),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_414),
.B(n_260),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_347),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_370),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_374),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_391),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_353),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_392),
.B(n_394),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_400),
.B(n_247),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_371),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_374),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_377),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_353),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_354),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_402),
.B(n_247),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_384),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_R g494 ( 
.A(n_410),
.B(n_238),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_412),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_377),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_422),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_354),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_378),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_429),
.Y(n_501)
);

BUFx10_ASAP7_75t_L g502 ( 
.A(n_434),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_444),
.B(n_175),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_497),
.B(n_373),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_429),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_479),
.B(n_497),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_483),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_483),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_425),
.Y(n_509)
);

NOR3xp33_ASAP7_75t_L g510 ( 
.A(n_428),
.B(n_341),
.C(n_352),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_447),
.B(n_422),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_462),
.B(n_407),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_483),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_433),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_461),
.A2(n_385),
.B1(n_235),
.B2(n_286),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_429),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_474),
.B(n_242),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_483),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_483),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_460),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_429),
.Y(n_521)
);

NAND3x1_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_335),
.C(n_334),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_426),
.A2(n_201),
.B1(n_309),
.B2(n_188),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_486),
.B(n_248),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_424),
.B(n_339),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_460),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_464),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_464),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_425),
.Y(n_530)
);

OR2x6_ASAP7_75t_L g531 ( 
.A(n_475),
.B(n_331),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_497),
.B(n_266),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_473),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_446),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_446),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_444),
.A2(n_381),
.B1(n_393),
.B2(n_406),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_497),
.B(n_444),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_492),
.B(n_250),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_425),
.B(n_240),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_466),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_497),
.B(n_430),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_497),
.B(n_378),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_L g543 ( 
.A1(n_425),
.A2(n_277),
.B1(n_226),
.B2(n_193),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_430),
.B(n_266),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_440),
.B(n_241),
.Y(n_546)
);

INVx4_ASAP7_75t_SL g547 ( 
.A(n_446),
.Y(n_547)
);

AND2x2_ASAP7_75t_SL g548 ( 
.A(n_457),
.B(n_184),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_448),
.B(n_379),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_446),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_448),
.B(n_244),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_452),
.B(n_252),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_469),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_452),
.B(n_379),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_472),
.B(n_255),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_433),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_453),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_472),
.B(n_257),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_437),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_476),
.B(n_380),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_449),
.B(n_296),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_445),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_431),
.B(n_258),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_445),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_449),
.B(n_296),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_431),
.B(n_435),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_498),
.B(n_380),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_449),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_470),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_R g571 ( 
.A(n_467),
.B(n_180),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_437),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_470),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_435),
.B(n_259),
.Y(n_574)
);

INVx4_ASAP7_75t_SL g575 ( 
.A(n_449),
.Y(n_575)
);

OAI22xp33_ASAP7_75t_L g576 ( 
.A1(n_467),
.A2(n_189),
.B1(n_220),
.B2(n_331),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_491),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_495),
.B(n_296),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_495),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_436),
.B(n_267),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_471),
.A2(n_335),
.B1(n_264),
.B2(n_322),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_494),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_436),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_491),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_491),
.B(n_296),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_439),
.B(n_268),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_491),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_439),
.B(n_274),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_441),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_441),
.B(n_282),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_478),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_491),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_499),
.B(n_296),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_499),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_454),
.B(n_283),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_478),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_481),
.A2(n_276),
.B1(n_190),
.B2(n_199),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_481),
.B(n_382),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_482),
.B(n_382),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_482),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_432),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_488),
.A2(n_249),
.B1(n_322),
.B2(n_319),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_493),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_454),
.B(n_289),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_499),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_458),
.B(n_292),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_499),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_488),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_489),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_SL g610 ( 
.A(n_432),
.B(n_281),
.C(n_336),
.Y(n_610)
);

OR2x6_ASAP7_75t_L g611 ( 
.A(n_489),
.B(n_184),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_496),
.B(n_386),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_499),
.B(n_190),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_458),
.B(n_297),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_496),
.B(n_386),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_500),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_500),
.B(n_303),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_468),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_468),
.B(n_199),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_468),
.B(n_397),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_465),
.B(n_397),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_443),
.A2(n_307),
.B1(n_332),
.B2(n_330),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_465),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_477),
.B(n_398),
.Y(n_624)
);

BUFx10_ASAP7_75t_L g625 ( 
.A(n_443),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_477),
.B(n_480),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_480),
.B(n_203),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_455),
.Y(n_628)
);

INVx6_ASAP7_75t_L g629 ( 
.A(n_455),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_456),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_R g631 ( 
.A(n_450),
.B(n_183),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_484),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_484),
.Y(n_633)
);

AND2x2_ASAP7_75t_SL g634 ( 
.A(n_490),
.B(n_203),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_490),
.B(n_204),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_456),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_450),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_427),
.B(n_204),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_463),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_438),
.B(n_209),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_463),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_442),
.B(n_398),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_451),
.B(n_209),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_459),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_487),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_483),
.Y(n_646)
);

INVx4_ASAP7_75t_SL g647 ( 
.A(n_425),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_494),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_548),
.B(n_304),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_517),
.B(n_212),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_537),
.A2(n_228),
.B(n_212),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_517),
.B(n_214),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_524),
.B(n_214),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_623),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_548),
.B(n_306),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_524),
.B(n_218),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_538),
.B(n_218),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_511),
.B(n_185),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_538),
.B(n_228),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_543),
.A2(n_233),
.B1(n_245),
.B2(n_249),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_597),
.A2(n_233),
.B1(n_319),
.B2(n_318),
.Y(n_661)
);

INVx8_ASAP7_75t_L g662 ( 
.A(n_644),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_512),
.A2(n_324),
.B1(n_316),
.B2(n_262),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_512),
.B(n_245),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_537),
.A2(n_316),
.B(n_264),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_545),
.B(n_262),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_545),
.A2(n_318),
.B1(n_265),
.B2(n_270),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_503),
.B(n_265),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_623),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_511),
.B(n_270),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_561),
.B(n_197),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_642),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_504),
.B(n_271),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_549),
.B(n_271),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_549),
.B(n_275),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_561),
.B(n_213),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_554),
.B(n_275),
.Y(n_677)
);

AND2x6_ASAP7_75t_SL g678 ( 
.A(n_638),
.B(n_399),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_603),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_558),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_568),
.B(n_216),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_589),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_568),
.B(n_198),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_554),
.A2(n_279),
.B1(n_299),
.B2(n_310),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_551),
.B(n_221),
.Y(n_685)
);

OR2x6_ASAP7_75t_L g686 ( 
.A(n_645),
.B(n_276),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_618),
.B(n_279),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_581),
.A2(n_310),
.B(n_299),
.C(n_415),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_618),
.B(n_399),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_582),
.B(n_198),
.Y(n_690)
);

AOI221xp5_ASAP7_75t_L g691 ( 
.A1(n_543),
.A2(n_308),
.B1(n_239),
.B2(n_263),
.C(n_269),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_558),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_542),
.B(n_609),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_506),
.A2(n_260),
.B1(n_313),
.B2(n_273),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_509),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_583),
.B(n_403),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_557),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_583),
.B(n_403),
.Y(n_698)
);

AOI221xp5_ASAP7_75t_SL g699 ( 
.A1(n_597),
.A2(n_419),
.B1(n_417),
.B2(n_415),
.C(n_411),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_541),
.A2(n_356),
.B(n_417),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_552),
.B(n_555),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_559),
.B(n_404),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_563),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_565),
.B(n_260),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_509),
.B(n_404),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_530),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_581),
.A2(n_419),
.B(n_411),
.C(n_409),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_563),
.Y(n_708)
);

O2A1O1Ixp5_ASAP7_75t_L g709 ( 
.A1(n_544),
.A2(n_409),
.B(n_356),
.C(n_260),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_589),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_530),
.B(n_329),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_520),
.B(n_327),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_565),
.B(n_326),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_565),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_616),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_616),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_526),
.B(n_323),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_648),
.B(n_198),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_533),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_602),
.A2(n_198),
.B1(n_314),
.B2(n_312),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_632),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_528),
.B(n_315),
.Y(n_722)
);

NAND3xp33_ASAP7_75t_L g723 ( 
.A(n_536),
.B(n_305),
.C(n_300),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_506),
.A2(n_298),
.B1(n_294),
.B2(n_293),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_529),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_598),
.Y(n_726)
);

AOI22x1_ASAP7_75t_L g727 ( 
.A1(n_540),
.A2(n_288),
.B1(n_287),
.B2(n_278),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_514),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_514),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_578),
.B(n_6),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_553),
.B(n_166),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_569),
.B(n_154),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_570),
.B(n_153),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_598),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_633),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_573),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_503),
.A2(n_146),
.B1(n_144),
.B2(n_126),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_536),
.A2(n_114),
.B1(n_104),
.B2(n_99),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_591),
.B(n_92),
.Y(n_739)
);

AND2x2_ASAP7_75t_SL g740 ( 
.A(n_602),
.B(n_84),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_596),
.B(n_78),
.Y(n_741)
);

NOR2x2_ASAP7_75t_L g742 ( 
.A(n_638),
.B(n_9),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_600),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_633),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_578),
.B(n_10),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_636),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_569),
.B(n_67),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_502),
.B(n_13),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_608),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_631),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_612),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_546),
.B(n_62),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_560),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_544),
.B(n_13),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_612),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_636),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_503),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_560),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_503),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_572),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_539),
.B(n_15),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_541),
.A2(n_23),
.B(n_25),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_617),
.B(n_26),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_572),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_564),
.B(n_26),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_574),
.B(n_30),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_647),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_621),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_626),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_595),
.B(n_31),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_580),
.B(n_31),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_604),
.B(n_53),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_502),
.B(n_32),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_629),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_606),
.B(n_52),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_575),
.B(n_33),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_629),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_624),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_614),
.B(n_50),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_571),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_634),
.B(n_50),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_508),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_571),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_575),
.B(n_40),
.Y(n_784)
);

NOR3xp33_ASAP7_75t_L g785 ( 
.A(n_523),
.B(n_576),
.C(n_610),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_586),
.B(n_43),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_628),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_634),
.B(n_44),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_630),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_556),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_567),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_647),
.B(n_47),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_588),
.B(n_47),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_592),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_620),
.B(n_48),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_525),
.B(n_49),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_620),
.B(n_49),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_644),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_590),
.B(n_550),
.Y(n_799)
);

O2A1O1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_619),
.A2(n_627),
.B(n_599),
.C(n_615),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_592),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_507),
.B(n_513),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_644),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_631),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_611),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_599),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_594),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_SL g808 ( 
.A(n_579),
.B(n_576),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_611),
.A2(n_622),
.B1(n_515),
.B2(n_522),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_508),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_510),
.B(n_611),
.C(n_615),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_501),
.B(n_505),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_735),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_679),
.Y(n_814)
);

OAI21x1_ASAP7_75t_L g815 ( 
.A1(n_812),
.A2(n_807),
.B(n_801),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_740),
.A2(n_619),
.B1(n_635),
.B2(n_566),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_660),
.A2(n_613),
.B(n_566),
.C(n_562),
.Y(n_817)
);

AO21x1_ASAP7_75t_L g818 ( 
.A1(n_730),
.A2(n_613),
.B(n_532),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_799),
.A2(n_518),
.B(n_519),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_740),
.A2(n_635),
.B1(n_562),
.B2(n_627),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_661),
.A2(n_660),
.B1(n_745),
.B2(n_730),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_714),
.A2(n_693),
.B(n_695),
.Y(n_822)
);

AOI21x1_ASAP7_75t_L g823 ( 
.A1(n_802),
.A2(n_532),
.B(n_521),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_714),
.A2(n_646),
.B(n_518),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_701),
.B(n_647),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_695),
.A2(n_646),
.B(n_519),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_658),
.A2(n_637),
.B(n_641),
.C(n_607),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_734),
.B(n_579),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_701),
.A2(n_508),
.B(n_605),
.Y(n_829)
);

NOR3xp33_ASAP7_75t_L g830 ( 
.A(n_658),
.B(n_601),
.C(n_645),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_791),
.B(n_501),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_706),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_672),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_734),
.B(n_639),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_750),
.B(n_531),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_806),
.B(n_505),
.Y(n_836)
);

NOR2x1_ASAP7_75t_L g837 ( 
.A(n_803),
.B(n_531),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_682),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_668),
.A2(n_705),
.B(n_800),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_676),
.B(n_535),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_732),
.A2(n_605),
.B(n_587),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_710),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_673),
.A2(n_607),
.B(n_594),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_732),
.A2(n_587),
.B(n_605),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_681),
.A2(n_584),
.B(n_577),
.C(n_516),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_710),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_747),
.A2(n_527),
.B(n_534),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_744),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_681),
.A2(n_585),
.B(n_593),
.C(n_639),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_747),
.A2(n_534),
.B(n_585),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_650),
.A2(n_593),
.B(n_639),
.C(n_644),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_670),
.A2(n_635),
.B(n_531),
.C(n_638),
.Y(n_852)
);

OAI21xp33_ASAP7_75t_L g853 ( 
.A1(n_664),
.A2(n_640),
.B(n_643),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_746),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_683),
.B(n_639),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_795),
.A2(n_534),
.B(n_575),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_769),
.A2(n_534),
.B(n_547),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_652),
.A2(n_640),
.B(n_643),
.C(n_625),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_719),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_653),
.B(n_547),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_666),
.A2(n_547),
.B(n_640),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_797),
.A2(n_643),
.B(n_625),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_706),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_656),
.B(n_657),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_661),
.A2(n_659),
.B1(n_734),
.B2(n_804),
.Y(n_865)
);

OAI21x1_ASAP7_75t_L g866 ( 
.A1(n_801),
.A2(n_807),
.B(n_756),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_726),
.B(n_755),
.Y(n_867)
);

NOR3xp33_ASAP7_75t_L g868 ( 
.A(n_785),
.B(n_691),
.C(n_809),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_702),
.B(n_685),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_781),
.A2(n_788),
.B(n_745),
.C(n_649),
.Y(n_870)
);

AO32x1_ASAP7_75t_L g871 ( 
.A1(n_738),
.A2(n_736),
.A3(n_749),
.B1(n_725),
.B2(n_743),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_746),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_690),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_756),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_685),
.B(n_674),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_675),
.B(n_677),
.Y(n_876)
);

INVxp33_ASAP7_75t_SL g877 ( 
.A(n_798),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_768),
.B(n_778),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_689),
.B(n_763),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_734),
.A2(n_706),
.B1(n_715),
.B2(n_716),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_706),
.B(n_757),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_787),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_711),
.A2(n_767),
.B(n_752),
.Y(n_883)
);

CKINVDCx8_ASAP7_75t_R g884 ( 
.A(n_678),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_763),
.B(n_765),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_713),
.A2(n_794),
.B(n_696),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_765),
.B(n_766),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_L g888 ( 
.A(n_663),
.B(n_771),
.C(n_793),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_713),
.A2(n_698),
.B(n_774),
.Y(n_889)
);

CKINVDCx8_ASAP7_75t_R g890 ( 
.A(n_662),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_751),
.A2(n_708),
.B1(n_692),
.B2(n_703),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_789),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_649),
.A2(n_655),
.B1(n_766),
.B2(n_771),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_777),
.Y(n_894)
);

OAI21xp33_ASAP7_75t_L g895 ( 
.A1(n_720),
.A2(n_808),
.B(n_684),
.Y(n_895)
);

NAND2x1_ASAP7_75t_L g896 ( 
.A(n_782),
.B(n_810),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_718),
.B(n_811),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_758),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_731),
.A2(n_741),
.B(n_739),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_792),
.B(n_680),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_803),
.B(n_805),
.Y(n_901)
);

NOR3xp33_ASAP7_75t_L g902 ( 
.A(n_723),
.B(n_655),
.C(n_748),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_786),
.B(n_793),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_733),
.A2(n_810),
.B(n_782),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_662),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_728),
.A2(n_753),
.B(n_760),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_757),
.A2(n_759),
.B1(n_786),
.B2(n_770),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_729),
.A2(n_764),
.B(n_777),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_790),
.B(n_772),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_712),
.B(n_717),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_722),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_687),
.A2(n_654),
.B(n_721),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_775),
.B(n_779),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_669),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_805),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_792),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_754),
.B(n_704),
.Y(n_917)
);

NOR3xp33_ASAP7_75t_L g918 ( 
.A(n_773),
.B(n_796),
.C(n_784),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_757),
.A2(n_759),
.B(n_776),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_757),
.A2(n_759),
.B(n_776),
.Y(n_920)
);

AOI21x1_ASAP7_75t_L g921 ( 
.A1(n_700),
.A2(n_651),
.B(n_665),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_686),
.B(n_759),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_686),
.Y(n_923)
);

OAI22xp33_ASAP7_75t_L g924 ( 
.A1(n_780),
.A2(n_783),
.B1(n_784),
.B2(n_694),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_SL g925 ( 
.A1(n_662),
.A2(n_761),
.B1(n_697),
.B2(n_686),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_724),
.B(n_667),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_737),
.B(n_709),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_762),
.A2(n_707),
.B(n_688),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_699),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_707),
.A2(n_688),
.B(n_727),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_720),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_742),
.B(n_750),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_800),
.A2(n_701),
.B(n_791),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_682),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_682),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_735),
.Y(n_936)
);

AOI21xp33_ASAP7_75t_L g937 ( 
.A1(n_658),
.A2(n_676),
.B(n_671),
.Y(n_937)
);

NOR2x1_ASAP7_75t_L g938 ( 
.A(n_803),
.B(n_582),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_740),
.A2(n_701),
.B1(n_791),
.B2(n_806),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_682),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_799),
.A2(n_714),
.B(n_693),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_740),
.B(n_701),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_799),
.A2(n_714),
.B(n_693),
.Y(n_943)
);

INVx4_ASAP7_75t_L g944 ( 
.A(n_706),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_750),
.B(n_804),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_701),
.B(n_791),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_701),
.B(n_791),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_701),
.B(n_791),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_682),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_734),
.B(n_557),
.Y(n_950)
);

AOI21x1_ASAP7_75t_L g951 ( 
.A1(n_812),
.A2(n_802),
.B(n_799),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_679),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_701),
.B(n_791),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_679),
.Y(n_954)
);

O2A1O1Ixp5_ASAP7_75t_SL g955 ( 
.A1(n_670),
.A2(n_650),
.B(n_653),
.C(n_652),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_799),
.A2(n_714),
.B(n_693),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_701),
.B(n_791),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_658),
.A2(n_701),
.B(n_676),
.C(n_681),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_750),
.B(n_804),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_740),
.A2(n_701),
.B1(n_791),
.B2(n_806),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_701),
.B(n_791),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_658),
.A2(n_701),
.B(n_676),
.C(n_681),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_679),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_660),
.A2(n_670),
.B(n_664),
.C(n_781),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_799),
.A2(n_714),
.B(n_693),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_706),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_701),
.A2(n_740),
.B1(n_658),
.B2(n_791),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_672),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_750),
.B(n_804),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_740),
.A2(n_701),
.B1(n_791),
.B2(n_806),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_734),
.B(n_557),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_701),
.B(n_791),
.Y(n_972)
);

NAND3xp33_ASAP7_75t_L g973 ( 
.A(n_658),
.B(n_676),
.C(n_671),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_800),
.A2(n_701),
.B(n_791),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_734),
.B(n_557),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_697),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_734),
.B(n_557),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_735),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_799),
.A2(n_714),
.B(n_693),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_660),
.A2(n_670),
.B(n_664),
.C(n_781),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_660),
.A2(n_670),
.B(n_664),
.C(n_781),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_679),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_701),
.B(n_791),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_740),
.A2(n_701),
.B1(n_791),
.B2(n_806),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_672),
.B(n_642),
.Y(n_985)
);

INVx3_ASAP7_75t_SL g986 ( 
.A(n_976),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_937),
.B(n_973),
.Y(n_987)
);

OAI22x1_ASAP7_75t_L g988 ( 
.A1(n_967),
.A2(n_893),
.B1(n_869),
.B2(n_888),
.Y(n_988)
);

NAND2x1_ASAP7_75t_L g989 ( 
.A(n_944),
.B(n_832),
.Y(n_989)
);

O2A1O1Ixp5_ASAP7_75t_L g990 ( 
.A1(n_958),
.A2(n_962),
.B(n_885),
.C(n_903),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_955),
.A2(n_887),
.B(n_875),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_SL g992 ( 
.A1(n_942),
.A2(n_974),
.B(n_933),
.Y(n_992)
);

AO31x2_ASAP7_75t_L g993 ( 
.A1(n_818),
.A2(n_939),
.A3(n_984),
.B(n_960),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_905),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_882),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_944),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_942),
.A2(n_870),
.B(n_869),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_946),
.B(n_947),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_866),
.A2(n_815),
.B(n_904),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_948),
.A2(n_961),
.B1(n_957),
.B2(n_972),
.Y(n_1000)
);

NAND2xp33_ASAP7_75t_L g1001 ( 
.A(n_821),
.B(n_970),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_823),
.A2(n_844),
.B(n_841),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_892),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_953),
.B(n_983),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_839),
.A2(n_980),
.B(n_964),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_855),
.B(n_873),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_945),
.B(n_959),
.Y(n_1007)
);

AO31x2_ASAP7_75t_L g1008 ( 
.A1(n_930),
.A2(n_928),
.A3(n_845),
.B(n_849),
.Y(n_1008)
);

AOI21x1_ASAP7_75t_L g1009 ( 
.A1(n_840),
.A2(n_951),
.B(n_829),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_945),
.B(n_959),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_956),
.A2(n_965),
.B(n_979),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_981),
.A2(n_876),
.B(n_917),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_910),
.B(n_864),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_910),
.A2(n_865),
.B(n_821),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_911),
.B(n_969),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_847),
.A2(n_843),
.B(n_886),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_915),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_877),
.Y(n_1018)
);

AO31x2_ASAP7_75t_L g1019 ( 
.A1(n_907),
.A2(n_827),
.A3(n_913),
.B(n_851),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_969),
.B(n_932),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_932),
.B(n_911),
.Y(n_1021)
);

NAND3xp33_ASAP7_75t_SL g1022 ( 
.A(n_868),
.B(n_895),
.C(n_830),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_879),
.B(n_931),
.Y(n_1023)
);

NAND3xp33_ASAP7_75t_L g1024 ( 
.A(n_868),
.B(n_926),
.C(n_918),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_SL g1025 ( 
.A(n_830),
.B(n_862),
.C(n_918),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_878),
.B(n_902),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_838),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_SL g1028 ( 
.A(n_902),
.B(n_926),
.C(n_852),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_899),
.A2(n_825),
.B(n_819),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_816),
.A2(n_817),
.B(n_889),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_842),
.Y(n_1031)
);

NAND3xp33_ASAP7_75t_SL g1032 ( 
.A(n_853),
.B(n_858),
.C(n_925),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_836),
.B(n_909),
.Y(n_1033)
);

AO31x2_ASAP7_75t_L g1034 ( 
.A1(n_880),
.A2(n_871),
.A3(n_891),
.B(n_860),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_833),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_846),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_883),
.A2(n_822),
.B(n_881),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_816),
.A2(n_820),
.B(n_920),
.Y(n_1038)
);

AOI21x1_ASAP7_75t_L g1039 ( 
.A1(n_927),
.A2(n_850),
.B(n_881),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_968),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_916),
.B(n_820),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_912),
.A2(n_826),
.B(n_921),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_916),
.B(n_831),
.Y(n_1043)
);

OAI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_985),
.A2(n_897),
.B(n_835),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_824),
.A2(n_906),
.B(n_908),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_915),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_924),
.B(n_935),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_857),
.A2(n_919),
.B(n_896),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_924),
.B(n_940),
.Y(n_1049)
);

NOR2x1_ASAP7_75t_L g1050 ( 
.A(n_905),
.B(n_859),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_934),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_835),
.B(n_954),
.Y(n_1052)
);

AO21x1_ASAP7_75t_L g1053 ( 
.A1(n_856),
.A2(n_861),
.B(n_834),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_854),
.A2(n_874),
.B(n_872),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_952),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_949),
.A2(n_898),
.B(n_936),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_952),
.B(n_954),
.Y(n_1057)
);

CKINVDCx8_ASAP7_75t_R g1058 ( 
.A(n_901),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_848),
.B(n_978),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_929),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_900),
.A2(n_966),
.B(n_863),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_832),
.A2(n_863),
.B(n_966),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_950),
.B(n_977),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_901),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_914),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_814),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_971),
.A2(n_975),
.B(n_894),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_894),
.A2(n_871),
.B(n_828),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_938),
.A2(n_837),
.B(n_929),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_871),
.A2(n_922),
.B(n_867),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_867),
.B(n_922),
.Y(n_1071)
);

AOI21xp33_ASAP7_75t_L g1072 ( 
.A1(n_963),
.A2(n_982),
.B(n_923),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_929),
.A2(n_925),
.B(n_890),
.Y(n_1073)
);

AND3x4_ASAP7_75t_L g1074 ( 
.A(n_884),
.B(n_785),
.C(n_830),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_929),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_958),
.A2(n_962),
.B(n_973),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_946),
.B(n_947),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_916),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_968),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_946),
.B(n_947),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_941),
.A2(n_714),
.B(n_943),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_958),
.A2(n_962),
.B(n_967),
.C(n_937),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_916),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_958),
.A2(n_962),
.B(n_967),
.C(n_937),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_815),
.A2(n_866),
.B(n_823),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_946),
.B(n_947),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_815),
.A2(n_866),
.B(n_823),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_815),
.A2(n_866),
.B(n_823),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_985),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_968),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_968),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_866),
.A2(n_815),
.B(n_904),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_946),
.B(n_947),
.Y(n_1093)
);

AO31x2_ASAP7_75t_L g1094 ( 
.A1(n_818),
.A2(n_962),
.A3(n_958),
.B(n_960),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_958),
.A2(n_962),
.B(n_973),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_946),
.B(n_947),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_944),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_915),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_882),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_958),
.A2(n_962),
.B(n_967),
.C(n_937),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_946),
.B(n_947),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_941),
.A2(n_714),
.B(n_943),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_916),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_813),
.Y(n_1104)
);

NAND2x1_ASAP7_75t_L g1105 ( 
.A(n_944),
.B(n_767),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_946),
.B(n_947),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_SL g1107 ( 
.A1(n_958),
.A2(n_962),
.B(n_942),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_866),
.A2(n_815),
.B(n_904),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_818),
.A2(n_962),
.A3(n_958),
.B(n_960),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_937),
.B(n_973),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_866),
.A2(n_815),
.B(n_904),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_968),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_813),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_SL g1114 ( 
.A(n_976),
.B(n_432),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_958),
.A2(n_962),
.B(n_973),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_869),
.B(n_683),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_882),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_866),
.A2(n_815),
.B(n_904),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_941),
.A2(n_714),
.B(n_943),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_937),
.B(n_958),
.Y(n_1120)
);

O2A1O1Ixp5_ASAP7_75t_L g1121 ( 
.A1(n_937),
.A2(n_962),
.B(n_958),
.C(n_885),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_866),
.A2(n_815),
.B(n_904),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_958),
.A2(n_962),
.B(n_973),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_946),
.B(n_947),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_941),
.A2(n_714),
.B(n_943),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_866),
.A2(n_815),
.B(n_904),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_958),
.A2(n_962),
.B(n_973),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_1035),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1064),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_1046),
.Y(n_1130)
);

BUFx10_ASAP7_75t_L g1131 ( 
.A(n_1018),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1013),
.B(n_998),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_1090),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1000),
.B(n_1077),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_1073),
.B(n_1064),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1080),
.B(n_1086),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_1071),
.B(n_1050),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_987),
.A2(n_1110),
.B1(n_1022),
.B2(n_1024),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1014),
.A2(n_1096),
.B1(n_1124),
.B2(n_1106),
.Y(n_1139)
);

NOR2x1_ASAP7_75t_L g1140 ( 
.A(n_994),
.B(n_1066),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1090),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1082),
.A2(n_1084),
.B(n_1100),
.C(n_987),
.Y(n_1142)
);

NAND2x1p5_ASAP7_75t_L g1143 ( 
.A(n_996),
.B(n_1097),
.Y(n_1143)
);

OR2x2_ASAP7_75t_L g1144 ( 
.A(n_1004),
.B(n_1022),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1015),
.B(n_1093),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1110),
.A2(n_1121),
.B(n_1084),
.C(n_1100),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1101),
.B(n_1010),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_SL g1148 ( 
.A(n_1018),
.B(n_1058),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1006),
.B(n_1091),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1116),
.B(n_1020),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1010),
.B(n_1007),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1021),
.B(n_1089),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1091),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1089),
.B(n_1052),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1052),
.B(n_1017),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1040),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1078),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_986),
.Y(n_1158)
);

INVx8_ASAP7_75t_L g1159 ( 
.A(n_1078),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1003),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_1078),
.Y(n_1161)
);

AO21x2_ASAP7_75t_L g1162 ( 
.A1(n_1005),
.A2(n_1030),
.B(n_991),
.Y(n_1162)
);

BUFx12f_ASAP7_75t_L g1163 ( 
.A(n_1066),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1112),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1028),
.A2(n_1001),
.B1(n_1025),
.B2(n_988),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1099),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_1055),
.B(n_1057),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1017),
.B(n_1098),
.Y(n_1168)
);

CKINVDCx6p67_ASAP7_75t_R g1169 ( 
.A(n_986),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1078),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1079),
.Y(n_1171)
);

BUFx12f_ASAP7_75t_L g1172 ( 
.A(n_1083),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1117),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1023),
.B(n_1012),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_994),
.B(n_1065),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1083),
.Y(n_1176)
);

INVx8_ASAP7_75t_L g1177 ( 
.A(n_1083),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1027),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1098),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_1083),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1026),
.B(n_1001),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1082),
.A2(n_1120),
.B(n_1025),
.C(n_1028),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_1075),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_1060),
.Y(n_1184)
);

BUFx8_ASAP7_75t_SL g1185 ( 
.A(n_1103),
.Y(n_1185)
);

AO21x2_ASAP7_75t_L g1186 ( 
.A1(n_1076),
.A2(n_1127),
.B(n_1123),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1031),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_1060),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1047),
.B(n_1049),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1075),
.Y(n_1190)
);

OR2x2_ASAP7_75t_SL g1191 ( 
.A(n_1032),
.B(n_1074),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1011),
.A2(n_1102),
.B(n_1081),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1103),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_996),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1103),
.Y(n_1195)
);

O2A1O1Ixp5_ASAP7_75t_SL g1196 ( 
.A1(n_1120),
.A2(n_1115),
.B(n_1095),
.C(n_997),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1033),
.B(n_1063),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1063),
.B(n_1044),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1036),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1097),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1032),
.A2(n_1074),
.B1(n_1038),
.B2(n_1041),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1051),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1119),
.A2(n_1125),
.B(n_1107),
.Y(n_1203)
);

AO21x1_ASAP7_75t_L g1204 ( 
.A1(n_1068),
.A2(n_1070),
.B(n_1037),
.Y(n_1204)
);

AOI222xp33_ASAP7_75t_L g1205 ( 
.A1(n_1114),
.A2(n_1043),
.B1(n_1056),
.B2(n_1113),
.C1(n_1104),
.C2(n_1059),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_992),
.A2(n_1113),
.B1(n_1104),
.B2(n_1121),
.Y(n_1206)
);

INVx5_ASAP7_75t_L g1207 ( 
.A(n_1072),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1094),
.B(n_1109),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1085),
.A2(n_1088),
.B(n_1087),
.Y(n_1209)
);

OR2x6_ASAP7_75t_L g1210 ( 
.A(n_1067),
.B(n_1069),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_989),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1054),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1094),
.B(n_1109),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1053),
.A2(n_1061),
.B1(n_1062),
.B2(n_1029),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1105),
.Y(n_1215)
);

CKINVDCx14_ASAP7_75t_R g1216 ( 
.A(n_990),
.Y(n_1216)
);

INVxp67_ASAP7_75t_SL g1217 ( 
.A(n_1039),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1019),
.B(n_1048),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1016),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1094),
.B(n_1109),
.Y(n_1220)
);

OR2x6_ASAP7_75t_L g1221 ( 
.A(n_1085),
.B(n_1088),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1094),
.B(n_1109),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_1019),
.Y(n_1223)
);

NAND2x1p5_ASAP7_75t_L g1224 ( 
.A(n_1087),
.B(n_1045),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_993),
.B(n_1019),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_993),
.B(n_1008),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1008),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1042),
.A2(n_1002),
.B(n_999),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_993),
.B(n_1034),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_993),
.B(n_1034),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1034),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1009),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1034),
.B(n_1092),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1108),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1111),
.B(n_1118),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_1122),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1126),
.A2(n_967),
.B1(n_808),
.B2(n_973),
.Y(n_1237)
);

O2A1O1Ixp5_ASAP7_75t_L g1238 ( 
.A1(n_1120),
.A2(n_937),
.B(n_962),
.C(n_958),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1116),
.B(n_937),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_1046),
.Y(n_1240)
);

AND2x2_ASAP7_75t_SL g1241 ( 
.A(n_1001),
.B(n_740),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1090),
.Y(n_1242)
);

CKINVDCx11_ASAP7_75t_R g1243 ( 
.A(n_986),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1064),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1035),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1064),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1064),
.B(n_1071),
.Y(n_1247)
);

CKINVDCx11_ASAP7_75t_R g1248 ( 
.A(n_986),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1121),
.A2(n_962),
.B(n_958),
.Y(n_1249)
);

CKINVDCx8_ASAP7_75t_R g1250 ( 
.A(n_1018),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1116),
.B(n_937),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1090),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1064),
.B(n_1071),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_995),
.Y(n_1254)
);

BUFx4_ASAP7_75t_SL g1255 ( 
.A(n_1090),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_1046),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1013),
.B(n_1000),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1013),
.B(n_1000),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1013),
.A2(n_967),
.B1(n_821),
.B2(n_1014),
.Y(n_1259)
);

OAI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1013),
.A2(n_967),
.B1(n_808),
.B2(n_973),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1090),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1013),
.B(n_946),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1013),
.B(n_1000),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1090),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1241),
.A2(n_1259),
.B1(n_1239),
.B2(n_1251),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1201),
.A2(n_1138),
.B1(n_1259),
.B2(n_1165),
.Y(n_1266)
);

OR2x6_ASAP7_75t_L g1267 ( 
.A(n_1135),
.B(n_1182),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1128),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1216),
.A2(n_1207),
.B1(n_1249),
.B2(n_1147),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1157),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1160),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1245),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1157),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1138),
.B(n_1144),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1166),
.Y(n_1275)
);

BUFx10_ASAP7_75t_L g1276 ( 
.A(n_1141),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1168),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1181),
.B(n_1197),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_1243),
.Y(n_1279)
);

CKINVDCx11_ASAP7_75t_R g1280 ( 
.A(n_1250),
.Y(n_1280)
);

INVx4_ASAP7_75t_L g1281 ( 
.A(n_1194),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1173),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1254),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1178),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1132),
.A2(n_1136),
.B1(n_1262),
.B2(n_1147),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1260),
.A2(n_1186),
.B1(n_1181),
.B2(n_1249),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1187),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1185),
.Y(n_1288)
);

INVx3_ASAP7_75t_SL g1289 ( 
.A(n_1169),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1199),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1159),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1186),
.A2(n_1207),
.B1(n_1198),
.B2(n_1139),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1157),
.Y(n_1293)
);

INVx6_ASAP7_75t_L g1294 ( 
.A(n_1194),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1141),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1161),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1228),
.A2(n_1203),
.B(n_1192),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1238),
.B(n_1142),
.C(n_1196),
.Y(n_1298)
);

CKINVDCx6p67_ASAP7_75t_R g1299 ( 
.A(n_1248),
.Y(n_1299)
);

AO21x1_ASAP7_75t_L g1300 ( 
.A1(n_1237),
.A2(n_1257),
.B(n_1263),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1151),
.A2(n_1145),
.B1(n_1207),
.B2(n_1148),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1179),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1202),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1224),
.A2(n_1214),
.B(n_1235),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1139),
.A2(n_1150),
.B1(n_1135),
.B2(n_1162),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1245),
.Y(n_1306)
);

INVx3_ASAP7_75t_SL g1307 ( 
.A(n_1158),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1194),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1161),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1255),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1135),
.A2(n_1162),
.B1(n_1134),
.B2(n_1149),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1134),
.A2(n_1149),
.B1(n_1258),
.B2(n_1263),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1183),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1152),
.B(n_1154),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1190),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1184),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1184),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1188),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1247),
.B(n_1253),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1170),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1188),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1171),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1155),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1191),
.A2(n_1167),
.B1(n_1252),
.B2(n_1257),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1180),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1131),
.Y(n_1326)
);

NAND2x1p5_ASAP7_75t_L g1327 ( 
.A(n_1218),
.B(n_1223),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1224),
.A2(n_1209),
.B(n_1206),
.Y(n_1328)
);

AO21x2_ASAP7_75t_L g1329 ( 
.A1(n_1233),
.A2(n_1204),
.B(n_1146),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1247),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1189),
.B(n_1174),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1232),
.Y(n_1332)
);

AOI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1234),
.A2(n_1233),
.B(n_1212),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1167),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1195),
.B(n_1137),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1227),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1222),
.B(n_1213),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1200),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1174),
.Y(n_1339)
);

INVxp33_ASAP7_75t_L g1340 ( 
.A(n_1242),
.Y(n_1340)
);

AO21x2_ASAP7_75t_L g1341 ( 
.A1(n_1217),
.A2(n_1225),
.B(n_1226),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1200),
.Y(n_1342)
);

BUFx8_ASAP7_75t_L g1343 ( 
.A(n_1264),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1206),
.A2(n_1225),
.B(n_1220),
.Y(n_1344)
);

AO21x1_ASAP7_75t_L g1345 ( 
.A1(n_1208),
.A2(n_1230),
.B(n_1229),
.Y(n_1345)
);

NOR2x1_ASAP7_75t_L g1346 ( 
.A(n_1140),
.B(n_1261),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1208),
.B(n_1231),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1219),
.Y(n_1348)
);

CKINVDCx8_ASAP7_75t_R g1349 ( 
.A(n_1141),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1156),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_SL g1351 ( 
.A1(n_1230),
.A2(n_1236),
.B(n_1210),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1176),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1221),
.Y(n_1353)
);

AOI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1148),
.A2(n_1175),
.B1(n_1164),
.B2(n_1205),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1176),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1130),
.A2(n_1256),
.B1(n_1240),
.B2(n_1175),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1205),
.A2(n_1221),
.B(n_1236),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1221),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1193),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1193),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1193),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1210),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1143),
.A2(n_1210),
.B(n_1215),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1133),
.A2(n_1153),
.B1(n_1246),
.B2(n_1129),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1159),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1129),
.B(n_1246),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1244),
.B(n_1246),
.Y(n_1367)
);

BUFx12f_ASAP7_75t_L g1368 ( 
.A(n_1131),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1211),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1177),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1244),
.Y(n_1371)
);

AOI222xp33_ASAP7_75t_L g1372 ( 
.A1(n_1163),
.A2(n_1241),
.B1(n_1001),
.B2(n_895),
.C1(n_973),
.C2(n_1024),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1177),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1211),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1172),
.A2(n_937),
.B1(n_868),
.B2(n_973),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1241),
.A2(n_808),
.B1(n_973),
.B2(n_479),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1185),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1241),
.A2(n_937),
.B1(n_868),
.B2(n_973),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1274),
.B(n_1347),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1278),
.B(n_1339),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1345),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1329),
.B(n_1347),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1362),
.B(n_1353),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1345),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1274),
.B(n_1278),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1265),
.B(n_1277),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1348),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1348),
.Y(n_1388)
);

AO21x2_ASAP7_75t_L g1389 ( 
.A1(n_1297),
.A2(n_1333),
.B(n_1300),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_1280),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1362),
.B(n_1353),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1337),
.B(n_1341),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1267),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1336),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1344),
.A2(n_1300),
.B(n_1328),
.Y(n_1395)
);

INVxp67_ASAP7_75t_L g1396 ( 
.A(n_1302),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1341),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1267),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1334),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1337),
.B(n_1358),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1334),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1277),
.B(n_1286),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1266),
.A2(n_1376),
.B1(n_1378),
.B2(n_1372),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1267),
.B(n_1305),
.Y(n_1404)
);

INVxp67_ASAP7_75t_SL g1405 ( 
.A(n_1298),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1363),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1358),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1267),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1343),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1323),
.B(n_1292),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1351),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1311),
.B(n_1312),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1285),
.A2(n_1375),
.B1(n_1269),
.B2(n_1331),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1343),
.Y(n_1414)
);

OR2x6_ASAP7_75t_L g1415 ( 
.A(n_1327),
.B(n_1304),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1357),
.B(n_1314),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1316),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1294),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1302),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1324),
.A2(n_1354),
.B1(n_1301),
.B2(n_1326),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1317),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1271),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1357),
.B(n_1332),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1350),
.B(n_1340),
.Y(n_1424)
);

BUFx2_ASAP7_75t_SL g1425 ( 
.A(n_1349),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1275),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1282),
.B(n_1283),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1284),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1287),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1290),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1303),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1318),
.B(n_1321),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1272),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1343),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1319),
.B(n_1330),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1306),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1313),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1338),
.A2(n_1342),
.B(n_1315),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1369),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1294),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1319),
.B(n_1335),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1268),
.B(n_1319),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1335),
.B(n_1325),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_1335),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1294),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1349),
.A2(n_1326),
.B1(n_1356),
.B2(n_1322),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1374),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1416),
.B(n_1352),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1438),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1406),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1416),
.B(n_1307),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1379),
.B(n_1340),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1440),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1383),
.B(n_1366),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1382),
.B(n_1355),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1382),
.B(n_1423),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1392),
.B(n_1307),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1423),
.B(n_1359),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1423),
.B(n_1360),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1400),
.B(n_1361),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1400),
.B(n_1320),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1383),
.B(n_1366),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1379),
.B(n_1309),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1433),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1385),
.B(n_1371),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1433),
.Y(n_1466)
);

NAND2x1p5_ASAP7_75t_L g1467 ( 
.A(n_1406),
.B(n_1308),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1385),
.B(n_1380),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1406),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1397),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1392),
.B(n_1367),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1403),
.A2(n_1299),
.B1(n_1368),
.B2(n_1289),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1424),
.B(n_1280),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1383),
.Y(n_1474)
);

AND2x4_ASAP7_75t_SL g1475 ( 
.A(n_1415),
.B(n_1281),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1380),
.B(n_1366),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1419),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1397),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1381),
.B(n_1364),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1417),
.B(n_1273),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1413),
.A2(n_1299),
.B1(n_1368),
.B2(n_1279),
.Y(n_1481)
);

NAND4xp25_ASAP7_75t_L g1482 ( 
.A(n_1413),
.B(n_1346),
.C(n_1310),
.D(n_1377),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1417),
.B(n_1293),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1381),
.B(n_1295),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1482),
.A2(n_1412),
.B1(n_1404),
.B2(n_1393),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1471),
.B(n_1437),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1482),
.A2(n_1412),
.B1(n_1393),
.B2(n_1398),
.Y(n_1487)
);

OAI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1481),
.A2(n_1420),
.B1(n_1446),
.B2(n_1405),
.C(n_1442),
.Y(n_1488)
);

NAND3xp33_ASAP7_75t_L g1489 ( 
.A(n_1481),
.B(n_1420),
.C(n_1405),
.Y(n_1489)
);

OR2x2_ASAP7_75t_SL g1490 ( 
.A(n_1451),
.B(n_1408),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1471),
.B(n_1437),
.Y(n_1491)
);

NOR3xp33_ASAP7_75t_L g1492 ( 
.A(n_1457),
.B(n_1446),
.C(n_1411),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_SL g1493 ( 
.A1(n_1467),
.A2(n_1434),
.B(n_1414),
.Y(n_1493)
);

AOI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1472),
.A2(n_1396),
.B1(n_1436),
.B2(n_1386),
.C(n_1419),
.Y(n_1494)
);

AOI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1464),
.A2(n_1396),
.B1(n_1436),
.B2(n_1386),
.C(n_1410),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1457),
.A2(n_1425),
.B1(n_1398),
.B2(n_1442),
.Y(n_1496)
);

AOI21xp33_ASAP7_75t_L g1497 ( 
.A1(n_1451),
.A2(n_1411),
.B(n_1408),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1468),
.B(n_1410),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1456),
.B(n_1384),
.Y(n_1499)
);

AOI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1464),
.A2(n_1384),
.B1(n_1402),
.B2(n_1407),
.C(n_1429),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1452),
.B(n_1421),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1479),
.B(n_1432),
.C(n_1422),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1452),
.B(n_1440),
.Y(n_1503)
);

NAND3xp33_ASAP7_75t_L g1504 ( 
.A(n_1479),
.B(n_1432),
.C(n_1422),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1473),
.B(n_1445),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1476),
.B(n_1402),
.Y(n_1506)
);

NAND3xp33_ASAP7_75t_L g1507 ( 
.A(n_1466),
.B(n_1407),
.C(n_1406),
.Y(n_1507)
);

AOI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1466),
.A2(n_1431),
.B1(n_1430),
.B2(n_1429),
.C(n_1426),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1476),
.A2(n_1425),
.B1(n_1409),
.B2(n_1434),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1455),
.B(n_1391),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1455),
.B(n_1415),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1475),
.A2(n_1389),
.B(n_1415),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1474),
.B(n_1415),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1474),
.B(n_1415),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1454),
.B(n_1445),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_L g1516 ( 
.A(n_1448),
.B(n_1387),
.C(n_1388),
.Y(n_1516)
);

AOI221xp5_ASAP7_75t_L g1517 ( 
.A1(n_1477),
.A2(n_1431),
.B1(n_1430),
.B2(n_1426),
.C(n_1443),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1454),
.A2(n_1399),
.B1(n_1401),
.B2(n_1441),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1465),
.B(n_1460),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1458),
.B(n_1459),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1458),
.B(n_1415),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1460),
.B(n_1428),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1458),
.B(n_1395),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1460),
.B(n_1428),
.Y(n_1524)
);

NAND4xp25_ASAP7_75t_L g1525 ( 
.A(n_1448),
.B(n_1427),
.C(n_1394),
.D(n_1443),
.Y(n_1525)
);

NAND3xp33_ASAP7_75t_L g1526 ( 
.A(n_1484),
.B(n_1394),
.C(n_1447),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1454),
.B(n_1409),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1477),
.A2(n_1414),
.B1(n_1434),
.B2(n_1444),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1484),
.B(n_1447),
.C(n_1439),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1523),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1502),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1490),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1522),
.Y(n_1533)
);

NOR2x1p5_ASAP7_75t_L g1534 ( 
.A(n_1489),
.B(n_1414),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1521),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1511),
.B(n_1450),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1499),
.B(n_1498),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1520),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1511),
.B(n_1450),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1524),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1490),
.B(n_1449),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1486),
.B(n_1470),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1526),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1516),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1529),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1513),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1526),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1491),
.B(n_1470),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1529),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1513),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1502),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1504),
.B(n_1478),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1504),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1489),
.A2(n_1435),
.B1(n_1441),
.B2(n_1463),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1514),
.Y(n_1555)
);

NAND3xp33_ASAP7_75t_L g1556 ( 
.A(n_1494),
.B(n_1483),
.C(n_1480),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1506),
.B(n_1501),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1514),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1544),
.B(n_1519),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1532),
.B(n_1510),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1532),
.B(n_1510),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1545),
.B(n_1525),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1532),
.B(n_1527),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1538),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1538),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1535),
.B(n_1546),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1544),
.B(n_1492),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1544),
.B(n_1495),
.Y(n_1568)
);

A2O1A1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1534),
.A2(n_1488),
.B(n_1485),
.C(n_1487),
.Y(n_1569)
);

NOR2x1_ASAP7_75t_L g1570 ( 
.A(n_1534),
.B(n_1493),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1538),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1538),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1530),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1551),
.Y(n_1574)
);

INVxp67_ASAP7_75t_L g1575 ( 
.A(n_1551),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1557),
.B(n_1289),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1557),
.B(n_1503),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1530),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1535),
.B(n_1515),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1556),
.B(n_1533),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1545),
.B(n_1480),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1545),
.B(n_1483),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1543),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1535),
.B(n_1469),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1530),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1556),
.B(n_1500),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1543),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1535),
.B(n_1469),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1533),
.B(n_1463),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1547),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1533),
.B(n_1463),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1547),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1535),
.B(n_1469),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1540),
.B(n_1517),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1540),
.B(n_1461),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1549),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1546),
.B(n_1550),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1549),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1573),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1586),
.B(n_1553),
.Y(n_1600)
);

INVxp67_ASAP7_75t_SL g1601 ( 
.A(n_1570),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1596),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1596),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1579),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1573),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1562),
.B(n_1553),
.Y(n_1606)
);

AOI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1569),
.A2(n_1531),
.B1(n_1509),
.B2(n_1554),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1560),
.B(n_1546),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1567),
.B(n_1531),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1570),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1598),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1563),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1598),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1568),
.A2(n_1493),
.B(n_1549),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1563),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1562),
.B(n_1552),
.Y(n_1616)
);

INVxp67_ASAP7_75t_SL g1617 ( 
.A(n_1574),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1560),
.B(n_1546),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1566),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1573),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1577),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1581),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1581),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1561),
.B(n_1550),
.Y(n_1624)
);

XNOR2x2_ASAP7_75t_L g1625 ( 
.A(n_1580),
.B(n_1541),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1594),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1578),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1582),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1566),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1561),
.B(n_1550),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1576),
.A2(n_1554),
.B1(n_1528),
.B2(n_1505),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1579),
.B(n_1550),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1575),
.A2(n_1587),
.B(n_1583),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1578),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1583),
.B(n_1541),
.Y(n_1635)
);

NAND2x1p5_ASAP7_75t_L g1636 ( 
.A(n_1587),
.B(n_1541),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1584),
.B(n_1555),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1582),
.Y(n_1638)
);

CKINVDCx20_ASAP7_75t_R g1639 ( 
.A(n_1559),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1590),
.B(n_1279),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1590),
.B(n_1552),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1612),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1602),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1602),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1626),
.B(n_1592),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1612),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1603),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1603),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1611),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1615),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1613),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1613),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1606),
.B(n_1592),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1601),
.B(n_1597),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1606),
.B(n_1564),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1625),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1600),
.B(n_1621),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1617),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1625),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1616),
.B(n_1564),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1622),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1639),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1622),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1607),
.A2(n_1512),
.B(n_1542),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1635),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1607),
.A2(n_1454),
.B1(n_1462),
.B2(n_1555),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1616),
.B(n_1565),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1609),
.B(n_1555),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1610),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1633),
.B(n_1555),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1623),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1636),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1623),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1614),
.B(n_1558),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1628),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1610),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1659),
.B(n_1640),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1648),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1651),
.Y(n_1680)
);

NAND2x1_ASAP7_75t_L g1681 ( 
.A(n_1660),
.B(n_1635),
.Y(n_1681)
);

OAI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1657),
.A2(n_1631),
.B1(n_1636),
.B2(n_1604),
.C(n_1641),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1648),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1642),
.B(n_1604),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1649),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1649),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1650),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1660),
.A2(n_1631),
.B(n_1641),
.Y(n_1688)
);

OAI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1666),
.A2(n_1628),
.B(n_1638),
.C(n_1619),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_1646),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1654),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1665),
.A2(n_1638),
.B1(n_1630),
.B2(n_1624),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1650),
.Y(n_1693)
);

O2A1O1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1670),
.A2(n_1636),
.B(n_1619),
.C(n_1629),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1655),
.B(n_1632),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1667),
.A2(n_1624),
.B1(n_1608),
.B2(n_1618),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1655),
.B(n_1632),
.Y(n_1697)
);

AOI222xp33_ASAP7_75t_L g1698 ( 
.A1(n_1658),
.A2(n_1608),
.B1(n_1630),
.B2(n_1618),
.C1(n_1629),
.C2(n_1637),
.Y(n_1698)
);

INVxp67_ASAP7_75t_SL g1699 ( 
.A(n_1673),
.Y(n_1699)
);

INVxp67_ASAP7_75t_SL g1700 ( 
.A(n_1673),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1663),
.A2(n_1558),
.B1(n_1589),
.B2(n_1591),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1645),
.B(n_1537),
.Y(n_1702)
);

OAI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1677),
.A2(n_1507),
.B1(n_1496),
.B2(n_1453),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1690),
.B(n_1662),
.Y(n_1704)
);

NAND2xp33_ASAP7_75t_SL g1705 ( 
.A(n_1681),
.B(n_1688),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1684),
.B(n_1675),
.Y(n_1706)
);

OR2x6_ASAP7_75t_L g1707 ( 
.A(n_1680),
.B(n_1288),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1684),
.B(n_1664),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1691),
.Y(n_1709)
);

INVxp33_ASAP7_75t_L g1710 ( 
.A(n_1678),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1691),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1695),
.B(n_1672),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1695),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1692),
.B(n_1654),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1697),
.B(n_1674),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1697),
.B(n_1699),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1679),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1700),
.B(n_1676),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1682),
.B(n_1671),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1689),
.B(n_1643),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1683),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1702),
.B(n_1390),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1685),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1705),
.A2(n_1694),
.B1(n_1703),
.B2(n_1686),
.C(n_1687),
.Y(n_1724)
);

NAND4xp25_ASAP7_75t_L g1725 ( 
.A(n_1719),
.B(n_1698),
.C(n_1693),
.D(n_1696),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1719),
.B(n_1703),
.C(n_1647),
.Y(n_1726)
);

OAI211xp5_ASAP7_75t_L g1727 ( 
.A1(n_1714),
.A2(n_1652),
.B(n_1644),
.C(n_1653),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1714),
.A2(n_1701),
.B(n_1652),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_SL g1729 ( 
.A1(n_1720),
.A2(n_1669),
.B1(n_1656),
.B2(n_1661),
.C(n_1668),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1713),
.A2(n_1656),
.B1(n_1661),
.B2(n_1668),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1706),
.B(n_1637),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1710),
.A2(n_1627),
.B1(n_1620),
.B2(n_1605),
.C(n_1599),
.Y(n_1732)
);

NAND3xp33_ASAP7_75t_L g1733 ( 
.A(n_1716),
.B(n_1634),
.C(n_1605),
.Y(n_1733)
);

OA21x2_ASAP7_75t_L g1734 ( 
.A1(n_1709),
.A2(n_1605),
.B(n_1599),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1722),
.A2(n_1634),
.B1(n_1599),
.B2(n_1627),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1734),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_SL g1737 ( 
.A1(n_1726),
.A2(n_1711),
.B1(n_1704),
.B2(n_1722),
.Y(n_1737)
);

NAND2xp33_ASAP7_75t_SL g1738 ( 
.A(n_1731),
.B(n_1708),
.Y(n_1738)
);

OAI211xp5_ASAP7_75t_L g1739 ( 
.A1(n_1724),
.A2(n_1718),
.B(n_1721),
.C(n_1723),
.Y(n_1739)
);

NOR3xp33_ASAP7_75t_L g1740 ( 
.A(n_1725),
.B(n_1715),
.C(n_1712),
.Y(n_1740)
);

NOR2x1_ASAP7_75t_L g1741 ( 
.A(n_1727),
.B(n_1707),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1733),
.Y(n_1742)
);

NAND3xp33_ASAP7_75t_L g1743 ( 
.A(n_1728),
.B(n_1707),
.C(n_1717),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1730),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1729),
.B(n_1707),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1735),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1732),
.Y(n_1747)
);

AOI211xp5_ASAP7_75t_L g1748 ( 
.A1(n_1739),
.A2(n_1377),
.B(n_1288),
.C(n_1627),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1744),
.B(n_1565),
.Y(n_1749)
);

NOR3xp33_ASAP7_75t_L g1750 ( 
.A(n_1737),
.B(n_1620),
.C(n_1295),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1741),
.B(n_1620),
.Y(n_1751)
);

NOR3xp33_ASAP7_75t_SL g1752 ( 
.A(n_1739),
.B(n_1497),
.C(n_1542),
.Y(n_1752)
);

OAI211xp5_ASAP7_75t_SL g1753 ( 
.A1(n_1745),
.A2(n_1740),
.B(n_1747),
.C(n_1746),
.Y(n_1753)
);

OAI221xp5_ASAP7_75t_SL g1754 ( 
.A1(n_1742),
.A2(n_1578),
.B1(n_1585),
.B2(n_1518),
.C(n_1572),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1751),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1749),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1753),
.A2(n_1738),
.B1(n_1743),
.B2(n_1736),
.Y(n_1757)
);

OAI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1752),
.A2(n_1572),
.B(n_1571),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1750),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1748),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1754),
.A2(n_1584),
.B1(n_1588),
.B2(n_1593),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1755),
.Y(n_1762)
);

NOR2x1p5_ASAP7_75t_L g1763 ( 
.A(n_1759),
.B(n_1760),
.Y(n_1763)
);

NOR3x1_ASAP7_75t_L g1764 ( 
.A(n_1756),
.B(n_1758),
.C(n_1757),
.Y(n_1764)
);

OAI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1761),
.A2(n_1585),
.B1(n_1571),
.B2(n_1548),
.C(n_1558),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1755),
.B(n_1597),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1762),
.B(n_1585),
.Y(n_1767)
);

INVx4_ASAP7_75t_L g1768 ( 
.A(n_1766),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1764),
.B(n_1588),
.Y(n_1769)
);

XNOR2xp5_ASAP7_75t_L g1770 ( 
.A(n_1769),
.B(n_1763),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1768),
.B1(n_1767),
.B2(n_1765),
.C(n_1373),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1771),
.B(n_1276),
.Y(n_1772)
);

OAI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1771),
.A2(n_1593),
.B(n_1595),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1772),
.B(n_1540),
.Y(n_1774)
);

NAND2xp33_ASAP7_75t_L g1775 ( 
.A(n_1773),
.B(n_1291),
.Y(n_1775)
);

OA22x2_ASAP7_75t_L g1776 ( 
.A1(n_1774),
.A2(n_1370),
.B1(n_1365),
.B2(n_1291),
.Y(n_1776)
);

AOI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1775),
.A2(n_1548),
.B1(n_1508),
.B2(n_1365),
.C(n_1281),
.Y(n_1777)
);

INVx2_ASAP7_75t_SL g1778 ( 
.A(n_1776),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1778),
.A2(n_1777),
.B1(n_1276),
.B2(n_1530),
.Y(n_1779)
);

AOI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1779),
.A2(n_1308),
.B1(n_1281),
.B2(n_1536),
.C(n_1539),
.Y(n_1780)
);

AOI211xp5_ASAP7_75t_L g1781 ( 
.A1(n_1780),
.A2(n_1418),
.B(n_1270),
.C(n_1296),
.Y(n_1781)
);


endmodule