module fake_jpeg_18102_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_SL g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_42),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_0),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_20),
.B1(n_25),
.B2(n_15),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_43),
.A2(n_35),
.B1(n_22),
.B2(n_31),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_20),
.B1(n_25),
.B2(n_15),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_48),
.B1(n_55),
.B2(n_35),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_41),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_32),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_17),
.B1(n_21),
.B2(n_23),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_24),
.B(n_19),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_26),
.B(n_24),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_67),
.B1(n_87),
.B2(n_47),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_34),
.C(n_50),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_56),
.B(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_69),
.Y(n_92)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_22),
.B(n_26),
.C(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_17),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_72),
.Y(n_95)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_74),
.Y(n_96)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_54),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_22),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_79),
.Y(n_99)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_18),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_51),
.B1(n_50),
.B2(n_47),
.Y(n_98)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_18),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_31),
.B1(n_37),
.B2(n_36),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_53),
.B1(n_45),
.B2(n_43),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_94),
.B1(n_109),
.B2(n_117),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_45),
.B1(n_51),
.B2(n_53),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_98),
.B1(n_104),
.B2(n_79),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_62),
.A3(n_76),
.B1(n_70),
.B2(n_67),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_112),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_60),
.A2(n_58),
.B1(n_36),
.B2(n_34),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_61),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_40),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_71),
.C(n_65),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_88),
.B(n_74),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_38),
.B1(n_54),
.B2(n_50),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_120),
.B(n_124),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g121 ( 
.A1(n_108),
.A2(n_89),
.B(n_84),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_121),
.A2(n_27),
.B(n_29),
.Y(n_179)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_146),
.C(n_139),
.Y(n_151)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_130),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_94),
.B1(n_124),
.B2(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_136),
.Y(n_169)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_24),
.B(n_27),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_118),
.B(n_91),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_90),
.A2(n_73),
.B1(n_72),
.B2(n_63),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_144),
.B1(n_114),
.B2(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_137),
.B(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_64),
.B1(n_68),
.B2(n_24),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_92),
.B(n_14),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_143),
.Y(n_174)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_68),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_88),
.B1(n_38),
.B2(n_40),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_24),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_59),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_149),
.A2(n_128),
.B1(n_126),
.B2(n_136),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_32),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_116),
.C(n_91),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_153),
.C(n_162),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_107),
.C(n_97),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_175),
.B1(n_29),
.B2(n_28),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_104),
.B1(n_110),
.B2(n_113),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_158),
.B1(n_127),
.B2(n_130),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_101),
.C(n_113),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_101),
.C(n_113),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_177),
.C(n_0),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_27),
.B(n_100),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_29),
.B(n_28),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_129),
.A2(n_138),
.B1(n_125),
.B2(n_122),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_176),
.B1(n_178),
.B2(n_4),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_121),
.A2(n_100),
.B1(n_93),
.B2(n_110),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_93),
.B1(n_114),
.B2(n_117),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_114),
.B1(n_103),
.B2(n_14),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_103),
.C(n_32),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_121),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_179),
.A2(n_29),
.B(n_28),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_186),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_133),
.B1(n_144),
.B2(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_189),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_190),
.B(n_202),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_205),
.B1(n_213),
.B2(n_159),
.Y(n_230)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_13),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_28),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_0),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_196),
.B(n_206),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_149),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_171),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_181),
.B(n_2),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_201),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_2),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_164),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_203),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_3),
.B(n_4),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_204),
.A2(n_212),
.B1(n_178),
.B2(n_166),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_151),
.B(n_4),
.Y(n_206)
);

OAI21x1_ASAP7_75t_R g207 ( 
.A1(n_159),
.A2(n_4),
.B(n_5),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_207),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_155),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_209),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_153),
.B(n_6),
.C(n_7),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_162),
.C(n_165),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_169),
.A2(n_6),
.B(n_7),
.Y(n_211)
);

AOI211xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_179),
.B(n_181),
.C(n_154),
.Y(n_220)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_160),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_230),
.B1(n_185),
.B2(n_204),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_210),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_234),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_177),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_237),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_185),
.B(n_197),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_188),
.C(n_196),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_190),
.C(n_183),
.Y(n_252)
);

FAx1_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_160),
.CI(n_176),
.CON(n_234),
.SN(n_234)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_159),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_242),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_225),
.B(n_199),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_248),
.Y(n_267)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_223),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_246),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_215),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_220),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_211),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_258),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_189),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_240),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_253),
.C(n_216),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_186),
.C(n_168),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_238),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_212),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_257),
.A2(n_228),
.B1(n_231),
.B2(n_224),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_237),
.B(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_227),
.B1(n_233),
.B2(n_234),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_261),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_268),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_264),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_247),
.A2(n_221),
.B(n_228),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_8),
.B(n_10),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_217),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_274),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_217),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_271),
.B(n_249),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_244),
.C(n_252),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_248),
.C(n_258),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_SL g273 ( 
.A1(n_239),
.A2(n_234),
.B(n_235),
.C(n_227),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_198),
.B1(n_207),
.B2(n_11),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_243),
.A2(n_229),
.B1(n_222),
.B2(n_213),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_166),
.B1(n_155),
.B2(n_168),
.Y(n_275)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_281),
.C(n_282),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_250),
.C(n_202),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_203),
.C(n_198),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_285),
.B(n_288),
.Y(n_300)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

XNOR2x1_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_207),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_11),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_8),
.C(n_10),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_290),
.A2(n_12),
.B(n_10),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_262),
.C(n_268),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_8),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_265),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_273),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_278),
.B(n_269),
.Y(n_293)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_283),
.A2(n_273),
.B1(n_276),
.B2(n_263),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_295),
.B1(n_301),
.B2(n_284),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_289),
.A2(n_273),
.B1(n_277),
.B2(n_271),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_302),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_291),
.C(n_284),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_12),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_280),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_307),
.B(n_310),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_282),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_281),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_288),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_312),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_294),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_298),
.C(n_295),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_316),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_310),
.B(n_304),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_318),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_317),
.A2(n_299),
.B(n_305),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_319),
.B(n_322),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

NOR3xp33_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_314),
.C(n_320),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_319),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_307),
.C(n_303),
.Y(n_328)
);


endmodule