module fake_jpeg_28749_n_537 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_537);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_537;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_15),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_53),
.B(n_82),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_54),
.B(n_85),
.Y(n_123)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g153 ( 
.A(n_68),
.Y(n_153)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_18),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_100),
.Y(n_150)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_41),
.Y(n_129)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_51),
.B1(n_25),
.B2(n_27),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_109),
.A2(n_131),
.B1(n_162),
.B2(n_44),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_51),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_63),
.B(n_22),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_128),
.B(n_40),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_135),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_64),
.A2(n_23),
.B1(n_27),
.B2(n_34),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_83),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_87),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_133),
.B(n_48),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_22),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_57),
.B(n_35),
.C(n_44),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_163),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_62),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_60),
.B(n_42),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_58),
.A2(n_43),
.B(n_35),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_165),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_105),
.A2(n_91),
.B1(n_67),
.B2(n_68),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_168),
.A2(n_185),
.B1(n_186),
.B2(n_207),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_73),
.B1(n_58),
.B2(n_24),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_169),
.A2(n_188),
.B1(n_216),
.B2(n_218),
.Y(n_231)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

INVx11_ASAP7_75t_L g260 ( 
.A(n_170),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_172),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_173),
.B(n_175),
.Y(n_229)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_174),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_163),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_176),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_165),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_177),
.B(n_181),
.Y(n_232)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_182),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_126),
.A2(n_75),
.B1(n_76),
.B2(n_97),
.Y(n_185)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_144),
.A2(n_73),
.B1(n_28),
.B2(n_48),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_190),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_123),
.B(n_119),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_191),
.B(n_202),
.Y(n_274)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_192),
.Y(n_270)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_195),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_123),
.A2(n_40),
.B(n_28),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_194),
.A2(n_217),
.B(n_167),
.Y(n_238)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_140),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_197),
.B(n_199),
.Y(n_250)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_201),
.Y(n_255)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_135),
.B(n_103),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_203),
.Y(n_259)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_204),
.B(n_205),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_130),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_206),
.B(n_208),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_105),
.A2(n_88),
.B1(n_89),
.B2(n_114),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_209),
.B(n_210),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_118),
.B(n_28),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_211),
.B(n_212),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_118),
.B(n_28),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_114),
.A2(n_102),
.B1(n_98),
.B2(n_49),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_217),
.B1(n_153),
.B2(n_161),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_134),
.B(n_49),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_223),
.C(n_153),
.Y(n_249)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_215),
.Y(n_261)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_108),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_139),
.A2(n_48),
.B1(n_17),
.B2(n_16),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_138),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_219),
.A2(n_221),
.B1(n_222),
.B2(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_111),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_220),
.Y(n_263)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_136),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

NAND2xp33_ASAP7_75t_SL g223 ( 
.A(n_127),
.B(n_48),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_146),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_138),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_225),
.A2(n_145),
.B1(n_150),
.B2(n_160),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_171),
.B(n_13),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_233),
.B(n_243),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_238),
.A2(n_267),
.B(n_214),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_173),
.B(n_161),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_239),
.B(n_266),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_194),
.B(n_13),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_177),
.B(n_184),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_244),
.B(n_9),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_249),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_167),
.B(n_13),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_273),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_179),
.A2(n_116),
.B1(n_106),
.B2(n_152),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_251),
.A2(n_253),
.B1(n_264),
.B2(n_268),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_179),
.A2(n_106),
.B1(n_150),
.B2(n_113),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_185),
.A2(n_160),
.B1(n_16),
.B2(n_15),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_202),
.B(n_0),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_223),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_188),
.A2(n_14),
.B1(n_5),
.B2(n_6),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_191),
.B(n_4),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_7),
.Y(n_310)
);

NOR4xp25_ASAP7_75t_SL g272 ( 
.A(n_169),
.B(n_14),
.C(n_6),
.D(n_7),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_272),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_221),
.B(n_14),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_255),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_302),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_276),
.B(n_283),
.Y(n_333)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_242),
.Y(n_278)
);

INVx4_ASAP7_75t_SL g320 ( 
.A(n_278),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_239),
.B(n_198),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_281),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_229),
.B(n_178),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_187),
.C(n_195),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_274),
.C(n_271),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_229),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_233),
.B(n_216),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_285),
.B(n_300),
.Y(n_341)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_238),
.A2(n_166),
.B(n_218),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_288),
.A2(n_289),
.B(n_301),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_243),
.A2(n_203),
.B(n_170),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_290),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_232),
.A2(n_176),
.B(n_192),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_291),
.A2(n_303),
.B(n_309),
.Y(n_355)
);

NAND2xp33_ASAP7_75t_SL g293 ( 
.A(n_249),
.B(n_225),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_298),
.Y(n_340)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_257),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_294),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_226),
.A2(n_168),
.B1(n_174),
.B2(n_172),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_295),
.A2(n_284),
.B1(n_264),
.B2(n_303),
.Y(n_319)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_297),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_219),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_250),
.B(n_5),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_307),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_232),
.Y(n_300)
);

NOR2x1_ASAP7_75t_L g301 ( 
.A(n_244),
.B(n_6),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_262),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_253),
.A2(n_244),
.B(n_251),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_304),
.B(n_263),
.Y(n_358)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

INVx3_ASAP7_75t_SL g306 ( 
.A(n_242),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_306),
.Y(n_348)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_227),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_262),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_315),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_246),
.A2(n_189),
.B(n_8),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_311),
.Y(n_338)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_227),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_313),
.Y(n_342)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_274),
.B(n_189),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_235),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_317),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_250),
.B(n_9),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_266),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_319),
.A2(n_325),
.B1(n_349),
.B2(n_279),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_322),
.B(n_314),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_281),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_324),
.B(n_353),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_283),
.A2(n_226),
.B1(n_245),
.B2(n_231),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_286),
.A2(n_254),
.B1(n_241),
.B2(n_259),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_326),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_288),
.A2(n_272),
.B1(n_265),
.B2(n_271),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_301),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_284),
.A2(n_279),
.B1(n_295),
.B2(n_280),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_332),
.A2(n_334),
.B1(n_293),
.B2(n_298),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_279),
.A2(n_274),
.B1(n_268),
.B2(n_265),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_335),
.B(n_337),
.C(n_343),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_282),
.B(n_269),
.C(n_247),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_247),
.C(n_261),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_302),
.B(n_273),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_345),
.B(n_356),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_290),
.A2(n_294),
.B1(n_287),
.B2(n_316),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_312),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_350),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_296),
.B(n_241),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_357),
.C(n_276),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_291),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_289),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_292),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_263),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_267),
.Y(n_357)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_358),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_298),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_374),
.C(n_379),
.Y(n_401)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_342),
.Y(n_360)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_361),
.A2(n_334),
.B1(n_339),
.B2(n_324),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_321),
.B(n_275),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_367),
.Y(n_398)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_365),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_301),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_369),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_370),
.A2(n_372),
.B1(n_325),
.B2(n_355),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_371),
.B(n_373),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_314),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_310),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_375),
.B(n_344),
.Y(n_394)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

OA21x2_ASAP7_75t_L g377 ( 
.A1(n_355),
.A2(n_315),
.B(n_267),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g421 ( 
.A1(n_377),
.A2(n_367),
.B(n_364),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_321),
.B(n_299),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_378),
.B(n_384),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_337),
.B(n_311),
.C(n_307),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_347),
.Y(n_380)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_380),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_343),
.B(n_317),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_389),
.C(n_346),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_347),
.B(n_305),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_387),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_386),
.Y(n_422)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_323),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_390),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_322),
.B(n_313),
.C(n_297),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_277),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_341),
.B(n_277),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_391),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_340),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_392),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_393),
.A2(n_292),
.B(n_329),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_394),
.B(n_400),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_366),
.B(n_371),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_396),
.B(n_397),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_340),
.Y(n_397)
);

MAJx2_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_340),
.C(n_323),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_415),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_363),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_403),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_407),
.B(n_421),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_372),
.A2(n_354),
.B1(n_331),
.B2(n_353),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_384),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_360),
.A2(n_319),
.B1(n_332),
.B2(n_339),
.Y(n_410)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_410),
.Y(n_447)
);

OAI22x1_ASAP7_75t_L g413 ( 
.A1(n_377),
.A2(n_381),
.B1(n_368),
.B2(n_339),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_413),
.A2(n_414),
.B(n_377),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_392),
.A2(n_327),
.B(n_336),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_374),
.B(n_357),
.Y(n_415)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_417),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_381),
.A2(n_327),
.B(n_336),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_418),
.A2(n_361),
.B(n_378),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_362),
.A2(n_346),
.B1(n_329),
.B2(n_338),
.Y(n_423)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_423),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_424),
.B(n_379),
.C(n_389),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_426),
.A2(n_428),
.B(n_434),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_422),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_432),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_359),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_395),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_375),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_437),
.C(n_442),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_413),
.A2(n_365),
.B(n_388),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_382),
.C(n_373),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_403),
.B(n_386),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_439),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_398),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_445),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_401),
.B(n_338),
.C(n_376),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_422),
.Y(n_443)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_443),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_406),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_401),
.B(n_369),
.C(n_352),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_450),
.C(n_394),
.Y(n_466)
);

FAx1_ASAP7_75t_SL g448 ( 
.A(n_411),
.B(n_309),
.CI(n_352),
.CON(n_448),
.SN(n_448)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_448),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_383),
.Y(n_449)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_449),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_395),
.B(n_259),
.C(n_236),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_424),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_462),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_466),
.C(n_429),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_431),
.A2(n_417),
.B1(n_407),
.B2(n_409),
.Y(n_457)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_457),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_447),
.A2(n_404),
.B1(n_408),
.B2(n_410),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_458),
.A2(n_465),
.B1(n_468),
.B2(n_425),
.Y(n_481)
);

NAND2x1_ASAP7_75t_SL g460 ( 
.A(n_428),
.B(n_418),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_397),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_448),
.B(n_421),
.Y(n_464)
);

CKINVDCx14_ASAP7_75t_R g480 ( 
.A(n_464),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_447),
.A2(n_421),
.B1(n_416),
.B2(n_402),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_444),
.A2(n_414),
.B1(n_420),
.B2(n_419),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_412),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_471),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_430),
.A2(n_434),
.B1(n_426),
.B2(n_439),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_470),
.A2(n_472),
.B1(n_443),
.B2(n_320),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_320),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_430),
.A2(n_320),
.B1(n_306),
.B2(n_278),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_473),
.B(n_230),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_466),
.C(n_442),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_483),
.C(n_489),
.Y(n_490)
);

AOI211xp5_ASAP7_75t_L g477 ( 
.A1(n_461),
.A2(n_430),
.B(n_448),
.C(n_435),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_477),
.A2(n_453),
.B1(n_463),
.B2(n_465),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_460),
.A2(n_449),
.B(n_450),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_478),
.A2(n_260),
.B(n_252),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_479),
.A2(n_237),
.B1(n_234),
.B2(n_248),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_469),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_446),
.C(n_433),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_454),
.B(n_437),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_485),
.Y(n_495)
);

FAx1_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_425),
.CI(n_348),
.CON(n_485),
.SN(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_458),
.A2(n_306),
.B1(n_254),
.B2(n_260),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_487),
.Y(n_499)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_459),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_261),
.C(n_242),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_462),
.C(n_471),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_491),
.B(n_497),
.C(n_500),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_492),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_498),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_477),
.A2(n_467),
.B(n_468),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_494),
.A2(n_481),
.B(n_482),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_482),
.A2(n_455),
.B(n_472),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_496),
.A2(n_486),
.B(n_485),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_452),
.C(n_254),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_236),
.C(n_228),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_501),
.B(n_502),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_480),
.B(n_234),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_478),
.B(n_260),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_503),
.B(n_485),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_504),
.B(n_488),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_476),
.Y(n_505)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_505),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_493),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_509),
.A2(n_506),
.B(n_510),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_514),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_513),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_474),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_495),
.B(n_473),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_515),
.B(n_491),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_519),
.B(n_522),
.Y(n_525)
);

AOI21x1_ASAP7_75t_L g524 ( 
.A1(n_520),
.A2(n_521),
.B(n_499),
.Y(n_524)
);

OAI221xp5_ASAP7_75t_L g521 ( 
.A1(n_509),
.A2(n_498),
.B1(n_494),
.B2(n_497),
.C(n_503),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_517),
.A2(n_508),
.B(n_511),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_523),
.B(n_518),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_524),
.B(n_526),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_516),
.B(n_508),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_527),
.A2(n_529),
.B(n_507),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_518),
.Y(n_529)
);

AOI21xp33_ASAP7_75t_L g530 ( 
.A1(n_528),
.A2(n_507),
.B(n_513),
.Y(n_530)
);

AOI21x1_ASAP7_75t_L g532 ( 
.A1(n_530),
.A2(n_531),
.B(n_500),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_237),
.B(n_248),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_237),
.C(n_240),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_534),
.A2(n_10),
.B(n_11),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_12),
.B(n_10),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_11),
.B(n_12),
.Y(n_537)
);


endmodule