module fake_jpeg_502_n_316 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_11),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_51),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_11),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_53),
.B(n_68),
.Y(n_132)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_55),
.A2(n_69),
.B1(n_28),
.B2(n_47),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_57),
.Y(n_117)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_10),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_64),
.Y(n_98)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_12),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_79),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_25),
.A2(n_12),
.B(n_1),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_19),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_70),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_33),
.B(n_9),
.Y(n_79)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_33),
.B(n_9),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_82),
.B(n_84),
.Y(n_137)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_35),
.B(n_13),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_86),
.B(n_88),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_42),
.B(n_14),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_91),
.Y(n_122)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_93),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_52),
.A2(n_28),
.B1(n_26),
.B2(n_36),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_96),
.A2(n_103),
.B1(n_106),
.B2(n_123),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_101),
.A2(n_118),
.B1(n_100),
.B2(n_97),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_125),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_36),
.B1(n_43),
.B2(n_47),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_23),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_114),
.B(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_39),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_74),
.A2(n_88),
.B1(n_86),
.B2(n_62),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_77),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_48),
.B(n_39),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_136),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_56),
.A2(n_40),
.B1(n_45),
.B2(n_0),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_130),
.A2(n_131),
.B1(n_117),
.B2(n_111),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_63),
.A2(n_15),
.B1(n_16),
.B2(n_71),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_51),
.B(n_55),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_87),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_72),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_70),
.A2(n_55),
.B1(n_69),
.B2(n_92),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_116),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_145),
.B(n_147),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_131),
.B1(n_130),
.B2(n_96),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_146),
.A2(n_157),
.B1(n_171),
.B2(n_162),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_110),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_152),
.Y(n_198)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_141),
.A2(n_124),
.B1(n_98),
.B2(n_104),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_159),
.A2(n_177),
.B1(n_178),
.B2(n_181),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_160),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_162),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_170),
.Y(n_192)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_168),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_127),
.C(n_94),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_99),
.C(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_95),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_173),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_121),
.B(n_142),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_172),
.B(n_179),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_113),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_128),
.B(n_144),
.C(n_106),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_180),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_97),
.A2(n_108),
.B1(n_109),
.B2(n_118),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_133),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_100),
.A2(n_142),
.B1(n_107),
.B2(n_115),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_184),
.B1(n_178),
.B2(n_183),
.Y(n_190)
);

CKINVDCx6p67_ASAP7_75t_R g183 ( 
.A(n_117),
.Y(n_183)
);

BUFx8_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_115),
.A2(n_103),
.B1(n_111),
.B2(n_109),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_99),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_145),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_201),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_159),
.B(n_185),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_209),
.B(n_191),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_200),
.B(n_212),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_170),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_155),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_205),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_157),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_169),
.B(n_154),
.CI(n_147),
.CON(n_211),
.SN(n_211)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_211),
.B(n_192),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_177),
.A2(n_152),
.B1(n_161),
.B2(n_173),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_213),
.B1(n_176),
.B2(n_183),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_229),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_158),
.C(n_149),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_235),
.C(n_217),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_192),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_222),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_180),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_SL g249 ( 
.A1(n_223),
.A2(n_228),
.A3(n_194),
.B1(n_199),
.B2(n_214),
.C1(n_203),
.C2(n_208),
.Y(n_249)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_190),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_156),
.B1(n_164),
.B2(n_167),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_226),
.A2(n_231),
.B1(n_186),
.B2(n_206),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_232),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_189),
.A2(n_150),
.B1(n_183),
.B2(n_165),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_166),
.B(n_195),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_233),
.A2(n_237),
.B(n_191),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_204),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_208),
.Y(n_256)
);

OA21x2_ASAP7_75t_SL g238 ( 
.A1(n_217),
.A2(n_211),
.B(n_210),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_238),
.B(n_242),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_244),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_243),
.B(n_241),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_190),
.B1(n_211),
.B2(n_186),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_241),
.A2(n_234),
.B1(n_222),
.B2(n_221),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_233),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_190),
.B(n_199),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_236),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_250),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_229),
.B1(n_215),
.B2(n_226),
.Y(n_264)
);

AOI221xp5_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_256),
.B1(n_231),
.B2(n_216),
.C(n_232),
.Y(n_262)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

NAND2xp33_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_235),
.Y(n_257)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_259),
.B(n_268),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_225),
.C(n_220),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_263),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_230),
.C(n_227),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_265),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_214),
.B1(n_227),
.B2(n_245),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_253),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_238),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_274),
.A2(n_248),
.B1(n_271),
.B2(n_267),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_247),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_261),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_247),
.B(n_243),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_265),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_259),
.A2(n_252),
.B(n_256),
.Y(n_281)
);

AO21x1_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_252),
.B(n_255),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_286),
.C(n_290),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_289),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_261),
.C(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_269),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_258),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_291),
.A2(n_281),
.B(n_279),
.Y(n_294)
);

OAI22x1_ASAP7_75t_L g292 ( 
.A1(n_283),
.A2(n_252),
.B1(n_264),
.B2(n_251),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_292),
.A2(n_291),
.B1(n_251),
.B2(n_246),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_280),
.Y(n_296)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_280),
.B1(n_255),
.B2(n_251),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_299),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_295),
.B(n_286),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_302),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_290),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_294),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_306),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_298),
.C(n_284),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_297),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_304),
.B1(n_276),
.B2(n_282),
.Y(n_310)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_307),
.B(n_276),
.CI(n_298),
.CON(n_309),
.SN(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_299),
.B(n_278),
.C(n_270),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_310),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_310),
.B(n_311),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_313),
.C(n_309),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_309),
.Y(n_316)
);


endmodule