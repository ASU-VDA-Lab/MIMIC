module fake_jpeg_30558_n_91 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_91);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_91;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx2_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_6),
.B(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx8_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_25),
.Y(n_32)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_0),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_19),
.B1(n_22),
.B2(n_11),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_12),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_10),
.C(n_11),
.Y(n_33)
);

AND2x6_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_38),
.Y(n_44)
);

AND2x6_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_27),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_22),
.B1(n_24),
.B2(n_23),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_23),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_46),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_48),
.B(n_50),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_33),
.C(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_57),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_39),
.B1(n_29),
.B2(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_28),
.B1(n_18),
.B2(n_16),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_21),
.B(n_17),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_49),
.B(n_11),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_67),
.B(n_54),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_46),
.B1(n_43),
.B2(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_58),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_28),
.C(n_18),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_56),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_18),
.B1(n_28),
.B2(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_52),
.C(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_13),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_72),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_15),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_74),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_60),
.B1(n_65),
.B2(n_63),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_68),
.Y(n_81)
);

AOI31xp33_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_69),
.A3(n_76),
.B(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_80),
.B(n_83),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_1),
.Y(n_86)
);

AOI31xp67_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_13),
.A3(n_14),
.B(n_9),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_75),
.B1(n_14),
.B2(n_3),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_1),
.B(n_2),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_87),
.A2(n_88),
.B1(n_85),
.B2(n_84),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.C1(n_8),
.C2(n_80),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_4),
.Y(n_91)
);


endmodule