module fake_netlist_5_2573_n_1832 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1832);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1832;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g179 ( 
.A(n_20),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_45),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_69),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_100),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_78),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_136),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_141),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_77),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_67),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_3),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_114),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_13),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_87),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_156),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_170),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_112),
.Y(n_201)
);

BUFx8_ASAP7_75t_SL g202 ( 
.A(n_166),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_80),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_10),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_145),
.Y(n_205)
);

BUFx8_ASAP7_75t_SL g206 ( 
.A(n_176),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_94),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_23),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_54),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_46),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_99),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_116),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_107),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_39),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_51),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_10),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_150),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_22),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_56),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_35),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_31),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_2),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_40),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_92),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_82),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_1),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_2),
.Y(n_229)
);

BUFx2_ASAP7_75t_SL g230 ( 
.A(n_70),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_132),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_20),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_146),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_124),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_76),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_134),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_163),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_143),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_153),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_5),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_67),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_88),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_14),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_34),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_120),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_121),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_177),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_97),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_125),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_149),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_65),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_157),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_38),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_73),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_102),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_35),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_65),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_36),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_56),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_30),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_135),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_155),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_60),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_18),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_57),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_41),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_41),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_37),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_75),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_165),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_25),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_91),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_162),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_21),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_110),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_148),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_106),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_115),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_51),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_12),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_53),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_32),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_15),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_59),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_98),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_86),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_74),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_53),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_93),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_44),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_101),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_72),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_18),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_130),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_21),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_66),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_129),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_152),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_140),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_104),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_0),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_34),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_164),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_58),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_174),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_81),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_24),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_113),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_142),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_127),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_84),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_123),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_42),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_168),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_117),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_55),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_154),
.Y(n_317)
);

BUFx2_ASAP7_75t_SL g318 ( 
.A(n_4),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_147),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_138),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_26),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_68),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_60),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_137),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_28),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_47),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_161),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_16),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_13),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_4),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_96),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_105),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_1),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_33),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_90),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_7),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_109),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_172),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_89),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_61),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_46),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_159),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_30),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_126),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_118),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_95),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_175),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_85),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_160),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_173),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_14),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_37),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_11),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_48),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_169),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_274),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_202),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_206),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_197),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_274),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_325),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_274),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_310),
.B(n_0),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_346),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_274),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_352),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_200),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_274),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_288),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_182),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_352),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_3),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_288),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_245),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_185),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_186),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_288),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_288),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_297),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_288),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_188),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_241),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_339),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_346),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_317),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_189),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_342),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_193),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_199),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_310),
.B(n_5),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_241),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_201),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_203),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_183),
.B(n_6),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_260),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_205),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_260),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_267),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_287),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_207),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_267),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_211),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_277),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_212),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_217),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_225),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_277),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_179),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_233),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_234),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_215),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_179),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_235),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_287),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_242),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_247),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_248),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_249),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_252),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_261),
.Y(n_420)
);

INVxp33_ASAP7_75t_L g421 ( 
.A(n_221),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_204),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_183),
.B(n_184),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_270),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_277),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_273),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_275),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_278),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_204),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_224),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_215),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_224),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_258),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_258),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_184),
.B(n_6),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_244),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_286),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_244),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_289),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_291),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_294),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_298),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_253),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_180),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_253),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_187),
.B(n_8),
.Y(n_446)
);

NAND2xp33_ASAP7_75t_R g447 ( 
.A(n_219),
.B(n_8),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_237),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_257),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_361),
.B(n_219),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_356),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_380),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_361),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_L g454 ( 
.A(n_363),
.B(n_284),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_388),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_366),
.B(n_187),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_433),
.B(n_191),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_389),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_399),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_356),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_360),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_360),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_380),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_362),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_392),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_384),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_R g467 ( 
.A(n_357),
.B(n_299),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_191),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_396),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_402),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_423),
.B(n_300),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_362),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_414),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_414),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_365),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_371),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_359),
.Y(n_479)
);

AND2x2_ASAP7_75t_SL g480 ( 
.A(n_390),
.B(n_239),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_384),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_404),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_405),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_407),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_365),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_368),
.B(n_355),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_431),
.B(n_213),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_413),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_368),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_369),
.B(n_303),
.Y(n_490)
);

OA21x2_ASAP7_75t_L g491 ( 
.A1(n_369),
.A2(n_263),
.B(n_257),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_407),
.B(n_192),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_367),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_374),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_373),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_373),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_377),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_417),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_419),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_447),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_377),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_364),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_424),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_421),
.B(n_231),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_378),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_378),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_408),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_437),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_371),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_364),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_444),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_444),
.B(n_196),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_439),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_444),
.B(n_196),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_382),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_384),
.B(n_198),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_382),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_391),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_448),
.B(n_198),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_448),
.B(n_220),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_412),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_412),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_440),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_R g525 ( 
.A(n_358),
.B(n_370),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_391),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_422),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_375),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_395),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_478),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_526),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_480),
.A2(n_491),
.B1(n_456),
.B2(n_435),
.Y(n_532)
);

OR2x6_ASAP7_75t_L g533 ( 
.A(n_492),
.B(n_318),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_455),
.Y(n_534)
);

BUFx10_ASAP7_75t_L g535 ( 
.A(n_504),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_511),
.B(n_376),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_511),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_511),
.B(n_381),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_478),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_480),
.B(n_385),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_479),
.Y(n_541)
);

AND2x6_ASAP7_75t_L g542 ( 
.A(n_456),
.B(n_220),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_500),
.B(n_385),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_500),
.B(n_425),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_504),
.B(n_386),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_491),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_491),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_471),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_502),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_509),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_491),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_471),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_511),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_L g554 ( 
.A(n_472),
.B(n_287),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_466),
.B(n_393),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_492),
.B(n_318),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_480),
.A2(n_400),
.B1(n_409),
.B2(n_406),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_459),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_502),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_526),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_459),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_473),
.B(n_403),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_466),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_480),
.A2(n_446),
.B1(n_394),
.B2(n_372),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_459),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_491),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_473),
.B(n_403),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_459),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_491),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_526),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_526),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_466),
.B(n_410),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_459),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_501),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_471),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_501),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_510),
.B(n_415),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_471),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_487),
.B(n_239),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_510),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_475),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_481),
.B(n_308),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_481),
.B(n_416),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_507),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_481),
.B(n_418),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_456),
.B(n_420),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_516),
.Y(n_587)
);

NAND3x1_ASAP7_75t_L g588 ( 
.A(n_457),
.B(n_265),
.C(n_263),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_518),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_457),
.A2(n_468),
.B1(n_372),
.B2(n_284),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_486),
.B(n_426),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_475),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_475),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_486),
.B(n_427),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_518),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_475),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_476),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_501),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_516),
.B(n_226),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_450),
.A2(n_428),
.B1(n_442),
.B2(n_441),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_522),
.Y(n_601)
);

BUFx6f_ASAP7_75t_SL g602 ( 
.A(n_522),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_501),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_457),
.B(n_422),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_523),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_490),
.B(n_236),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_476),
.Y(n_607)
);

OAI21xp33_ASAP7_75t_SL g608 ( 
.A1(n_468),
.A2(n_227),
.B(n_226),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_454),
.A2(n_279),
.B1(n_354),
.B2(n_353),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_512),
.B(n_308),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_454),
.A2(n_279),
.B1(n_354),
.B2(n_353),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_523),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_520),
.B(n_227),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_476),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_512),
.B(n_314),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_527),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_476),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_520),
.B(n_429),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_501),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_512),
.B(n_314),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_514),
.B(n_306),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_479),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_521),
.B(n_238),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_514),
.B(n_238),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_485),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_450),
.B(n_429),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_485),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_485),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_528),
.Y(n_629)
);

INVxp33_ASAP7_75t_SL g630 ( 
.A(n_467),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_517),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_527),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_451),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_521),
.B(n_246),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_521),
.B(n_430),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_528),
.B(n_194),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_451),
.B(n_430),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_460),
.B(n_309),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_485),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_517),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_453),
.B(n_432),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_460),
.B(n_311),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_461),
.B(n_432),
.Y(n_643)
);

AND2x2_ASAP7_75t_SL g644 ( 
.A(n_453),
.B(n_246),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_461),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_462),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_495),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_L g648 ( 
.A(n_462),
.B(n_287),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_464),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_464),
.B(n_436),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_474),
.B(n_477),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_484),
.B(n_194),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_517),
.Y(n_653)
);

INVxp33_ASAP7_75t_L g654 ( 
.A(n_525),
.Y(n_654)
);

INVx5_ASAP7_75t_L g655 ( 
.A(n_517),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_474),
.B(n_312),
.Y(n_656)
);

NAND2x1p5_ASAP7_75t_L g657 ( 
.A(n_517),
.B(n_250),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_477),
.B(n_250),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_484),
.B(n_436),
.Y(n_659)
);

INVx5_ASAP7_75t_L g660 ( 
.A(n_495),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_489),
.B(n_315),
.Y(n_661)
);

BUFx10_ASAP7_75t_L g662 ( 
.A(n_455),
.Y(n_662)
);

INVx11_ASAP7_75t_L g663 ( 
.A(n_458),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_495),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_529),
.B(n_254),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_458),
.A2(n_379),
.B1(n_387),
.B2(n_383),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_452),
.Y(n_667)
);

AND2x6_ASAP7_75t_L g668 ( 
.A(n_496),
.B(n_254),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_496),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_497),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_586),
.B(n_190),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_564),
.A2(n_280),
.B(n_265),
.C(n_321),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_606),
.B(n_497),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g674 ( 
.A(n_630),
.B(n_465),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_587),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_544),
.B(n_195),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_591),
.B(n_505),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_564),
.A2(n_608),
.B(n_594),
.C(n_591),
.Y(n_678)
);

AO22x1_ASAP7_75t_L g679 ( 
.A1(n_585),
.A2(n_321),
.B1(n_351),
.B2(n_280),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_546),
.B(n_194),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_587),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_562),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_594),
.B(n_506),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_532),
.B(n_506),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_532),
.A2(n_276),
.B1(n_255),
.B2(n_262),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_542),
.B(n_255),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_540),
.B(n_208),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_542),
.A2(n_320),
.B1(n_262),
.B2(n_269),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_546),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_542),
.B(n_269),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_540),
.B(n_209),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_567),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_542),
.B(n_272),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_542),
.B(n_272),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_543),
.B(n_210),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_584),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_604),
.B(n_276),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_626),
.B(n_214),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_546),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_546),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_R g701 ( 
.A(n_534),
.B(n_465),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_537),
.B(n_285),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_547),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_547),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_547),
.B(n_194),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_531),
.B(n_285),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_641),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_545),
.B(n_525),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_557),
.A2(n_344),
.B1(n_319),
.B2(n_322),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_589),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_547),
.B(n_287),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_531),
.B(n_292),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_595),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_551),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_551),
.B(n_287),
.Y(n_715)
);

OAI21xp33_ASAP7_75t_L g716 ( 
.A1(n_590),
.A2(n_330),
.B(n_326),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_537),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_659),
.B(n_469),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_551),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_551),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_566),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_566),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_530),
.B(n_292),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_539),
.B(n_320),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_536),
.A2(n_463),
.B(n_452),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_579),
.B(n_218),
.C(n_216),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_550),
.B(n_324),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_566),
.B(n_287),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_644),
.A2(n_349),
.B1(n_335),
.B2(n_347),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_601),
.Y(n_730)
);

INVxp67_ASAP7_75t_R g731 ( 
.A(n_555),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_566),
.B(n_287),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_605),
.Y(n_733)
);

NAND3xp33_ASAP7_75t_L g734 ( 
.A(n_579),
.B(n_228),
.C(n_222),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_569),
.B(n_337),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_612),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_616),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_632),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_569),
.B(n_305),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_538),
.A2(n_463),
.B(n_452),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_563),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_569),
.Y(n_742)
);

BUFx2_ASAP7_75t_L g743 ( 
.A(n_563),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_569),
.B(n_327),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_548),
.Y(n_745)
);

NOR2xp67_ASAP7_75t_SL g746 ( 
.A(n_631),
.B(n_230),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_549),
.B(n_470),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_SL g748 ( 
.A1(n_533),
.A2(n_493),
.B1(n_494),
.B2(n_296),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_559),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_631),
.B(n_331),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_621),
.A2(n_463),
.B(n_452),
.Y(n_751)
);

O2A1O1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_582),
.A2(n_334),
.B(n_351),
.C(n_326),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_560),
.B(n_337),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_570),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_618),
.B(n_338),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_631),
.B(n_332),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_580),
.B(n_240),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_552),
.Y(n_758)
);

NOR2xp67_ASAP7_75t_L g759 ( 
.A(n_600),
.B(n_470),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_624),
.A2(n_338),
.B1(n_345),
.B2(n_350),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_624),
.B(n_348),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_635),
.Y(n_762)
);

NAND2x1_ASAP7_75t_L g763 ( 
.A(n_561),
.B(n_515),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_666),
.B(n_482),
.Y(n_764)
);

INVx5_ASAP7_75t_L g765 ( 
.A(n_658),
.Y(n_765)
);

OAI22x1_ASAP7_75t_L g766 ( 
.A1(n_534),
.A2(n_482),
.B1(n_524),
.B2(n_513),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_577),
.Y(n_767)
);

NOR2xp67_ASAP7_75t_L g768 ( 
.A(n_585),
.B(n_483),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_640),
.B(n_653),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_633),
.B(n_515),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_553),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_535),
.B(n_483),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_645),
.B(n_519),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_640),
.B(n_653),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_535),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_553),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_646),
.B(n_519),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_L g778 ( 
.A(n_652),
.B(n_488),
.C(n_513),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_572),
.B(n_243),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_571),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_669),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_610),
.A2(n_519),
.B(n_529),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_670),
.B(n_519),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_571),
.Y(n_784)
);

NAND3xp33_ASAP7_75t_SL g785 ( 
.A(n_590),
.B(n_498),
.C(n_508),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_575),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_571),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_624),
.A2(n_498),
.B1(n_508),
.B2(n_503),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_575),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_651),
.B(n_529),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_624),
.A2(n_301),
.B1(n_229),
.B2(n_232),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_651),
.B(n_438),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_578),
.Y(n_793)
);

BUFx6f_ASAP7_75t_SL g794 ( 
.A(n_629),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_535),
.Y(n_795)
);

NOR3xp33_ASAP7_75t_L g796 ( 
.A(n_652),
.B(n_503),
.C(n_499),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_624),
.A2(n_499),
.B1(n_181),
.B2(n_223),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_599),
.B(n_438),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_640),
.B(n_251),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_665),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_613),
.A2(n_323),
.B1(n_329),
.B2(n_494),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_554),
.A2(n_330),
.B1(n_334),
.B2(n_341),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_578),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_581),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_653),
.B(n_256),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_571),
.B(n_259),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_613),
.B(n_443),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_654),
.B(n_192),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_576),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_623),
.A2(n_493),
.B1(n_304),
.B2(n_302),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_561),
.B(n_264),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_L g812 ( 
.A(n_658),
.B(n_266),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_623),
.A2(n_313),
.B1(n_268),
.B2(n_271),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_583),
.B(n_316),
.C(n_281),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_634),
.B(n_445),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_554),
.A2(n_341),
.B1(n_343),
.B2(n_192),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_665),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_581),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_634),
.A2(n_343),
.B(n_449),
.C(n_398),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_592),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_665),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_634),
.B(n_449),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_649),
.B(n_282),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_707),
.B(n_654),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_675),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_681),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_743),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_704),
.A2(n_573),
.B(n_561),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_677),
.B(n_582),
.Y(n_829)
);

AOI21x1_ASAP7_75t_L g830 ( 
.A1(n_680),
.A2(n_642),
.B(n_638),
.Y(n_830)
);

AOI21x1_ASAP7_75t_L g831 ( 
.A1(n_705),
.A2(n_661),
.B(n_656),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_767),
.B(n_630),
.Y(n_832)
);

OAI321xp33_ASAP7_75t_L g833 ( 
.A1(n_687),
.A2(n_533),
.A3(n_556),
.B1(n_609),
.B2(n_611),
.C(n_636),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_L g834 ( 
.A(n_678),
.B(n_533),
.C(n_556),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_692),
.B(n_556),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_771),
.Y(n_836)
);

OAI21xp5_ASAP7_75t_L g837 ( 
.A1(n_711),
.A2(n_620),
.B(n_615),
.Y(n_837)
);

INVx11_ASAP7_75t_L g838 ( 
.A(n_731),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_704),
.A2(n_573),
.B(n_598),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_711),
.A2(n_620),
.B(n_598),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_683),
.B(n_636),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_671),
.B(n_629),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_699),
.Y(n_843)
);

OR2x2_ASAP7_75t_SL g844 ( 
.A(n_785),
.B(n_541),
.Y(n_844)
);

AO21x1_ASAP7_75t_L g845 ( 
.A1(n_687),
.A2(n_657),
.B(n_648),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_800),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_715),
.A2(n_619),
.B(n_603),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_704),
.B(n_598),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_673),
.B(n_649),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_699),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_704),
.A2(n_573),
.B(n_603),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_769),
.A2(n_619),
.B(n_603),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_685),
.A2(n_609),
.B1(n_611),
.B2(n_668),
.Y(n_853)
);

AND2x2_ASAP7_75t_SL g854 ( 
.A(n_691),
.B(n_648),
.Y(n_854)
);

NAND2x1p5_ASAP7_75t_L g855 ( 
.A(n_699),
.B(n_558),
.Y(n_855)
);

NAND3xp33_ASAP7_75t_SL g856 ( 
.A(n_797),
.B(n_622),
.C(n_283),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_741),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_701),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_749),
.Y(n_859)
);

AOI33xp33_ASAP7_75t_L g860 ( 
.A1(n_762),
.A2(n_395),
.A3(n_397),
.B1(n_398),
.B2(n_401),
.B3(n_588),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_769),
.A2(n_619),
.B(n_657),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_817),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_684),
.A2(n_588),
.B1(n_558),
.B2(n_565),
.Y(n_863)
);

BUFx4f_ASAP7_75t_L g864 ( 
.A(n_775),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_671),
.B(n_695),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_808),
.B(n_629),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_774),
.A2(n_667),
.B(n_568),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_682),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_821),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_754),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_696),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_747),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_745),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_699),
.B(n_576),
.Y(n_874)
);

CKINVDCx10_ASAP7_75t_R g875 ( 
.A(n_794),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_751),
.A2(n_565),
.B(n_607),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_701),
.Y(n_877)
);

O2A1O1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_672),
.A2(n_637),
.B(n_643),
.C(n_650),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_698),
.B(n_662),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_720),
.A2(n_667),
.B(n_655),
.Y(n_880)
);

BUFx4f_ASAP7_75t_L g881 ( 
.A(n_795),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_698),
.B(n_637),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_739),
.A2(n_735),
.B(n_744),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_790),
.B(n_643),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_744),
.A2(n_655),
.B(n_597),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_779),
.B(n_650),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_695),
.B(n_708),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_717),
.Y(n_888)
);

CKINVDCx10_ASAP7_75t_R g889 ( 
.A(n_794),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_689),
.B(n_576),
.Y(n_890)
);

AOI21x1_ASAP7_75t_L g891 ( 
.A1(n_728),
.A2(n_732),
.B(n_746),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_716),
.A2(n_668),
.B1(n_658),
.B2(n_593),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_732),
.A2(n_593),
.B(n_596),
.Y(n_893)
);

OAI21x1_ASAP7_75t_L g894 ( 
.A1(n_725),
.A2(n_614),
.B(n_617),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_779),
.B(n_658),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_765),
.A2(n_596),
.B(n_614),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_792),
.B(n_658),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_765),
.A2(n_574),
.B(n_664),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_700),
.A2(n_714),
.B(n_703),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_676),
.B(n_662),
.Y(n_900)
);

NAND2xp33_ASAP7_75t_L g901 ( 
.A(n_787),
.B(n_814),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_719),
.A2(n_574),
.B(n_628),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_763),
.A2(n_647),
.B(n_639),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_799),
.A2(n_668),
.B1(n_602),
.B2(n_625),
.Y(n_904)
);

O2A1O1Ixp5_ASAP7_75t_L g905 ( 
.A1(n_686),
.A2(n_647),
.B(n_639),
.C(n_627),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_799),
.A2(n_805),
.B1(n_676),
.B2(n_811),
.Y(n_906)
);

NAND2x1p5_ASAP7_75t_L g907 ( 
.A(n_780),
.B(n_627),
.Y(n_907)
);

NOR3xp33_ASAP7_75t_L g908 ( 
.A(n_748),
.B(n_307),
.C(n_290),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_719),
.B(n_668),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_721),
.A2(n_660),
.B(n_668),
.Y(n_910)
);

AND2x2_ASAP7_75t_SL g911 ( 
.A(n_688),
.B(n_602),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_721),
.B(n_660),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_722),
.B(n_660),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_697),
.A2(n_822),
.B(n_815),
.C(n_807),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_798),
.A2(n_340),
.B(n_336),
.C(n_333),
.Y(n_915)
);

AOI21x1_ASAP7_75t_L g916 ( 
.A1(n_750),
.A2(n_660),
.B(n_133),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_742),
.A2(n_293),
.B(n_295),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_742),
.B(n_328),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_750),
.A2(n_756),
.B(n_784),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_710),
.B(n_9),
.Y(n_920)
);

BUFx4f_ASAP7_75t_L g921 ( 
.A(n_718),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_787),
.B(n_662),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_713),
.B(n_730),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_787),
.B(n_690),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_809),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_693),
.A2(n_694),
.B(n_805),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_733),
.B(n_11),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_757),
.A2(n_663),
.B(n_15),
.C(n_16),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_702),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_761),
.A2(n_171),
.B(n_158),
.Y(n_930)
);

AOI21x1_ASAP7_75t_L g931 ( 
.A1(n_706),
.A2(n_151),
.B(n_139),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_717),
.Y(n_932)
);

AO21x1_ASAP7_75t_L g933 ( 
.A1(n_811),
.A2(n_12),
.B(n_17),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_SL g934 ( 
.A(n_674),
.B(n_119),
.Y(n_934)
);

AOI21xp33_ASAP7_75t_L g935 ( 
.A1(n_729),
.A2(n_757),
.B(n_709),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_776),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_758),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_768),
.B(n_108),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_823),
.B(n_103),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_702),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_770),
.A2(n_71),
.B(n_19),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_736),
.B(n_737),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_738),
.B(n_17),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_773),
.A2(n_19),
.B(n_22),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_777),
.A2(n_23),
.B(n_25),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_783),
.A2(n_26),
.B(n_27),
.Y(n_946)
);

AOI21x1_ASAP7_75t_L g947 ( 
.A1(n_712),
.A2(n_27),
.B(n_29),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_782),
.A2(n_29),
.B(n_31),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_755),
.A2(n_32),
.B(n_33),
.C(n_36),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_781),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_L g951 ( 
.A(n_760),
.B(n_40),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_776),
.A2(n_66),
.B1(n_43),
.B2(n_44),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_740),
.A2(n_809),
.B(n_724),
.Y(n_953)
);

OAI321xp33_ASAP7_75t_L g954 ( 
.A1(n_816),
.A2(n_42),
.A3(n_43),
.B1(n_47),
.B2(n_48),
.C(n_49),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_702),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_806),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_758),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_753),
.Y(n_958)
);

OAI321xp33_ASAP7_75t_L g959 ( 
.A1(n_726),
.A2(n_50),
.A3(n_54),
.B1(n_55),
.B2(n_57),
.C(n_59),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_723),
.A2(n_61),
.B(n_62),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_727),
.A2(n_62),
.B(n_63),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_786),
.B(n_789),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_791),
.A2(n_64),
.B1(n_802),
.B2(n_759),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_786),
.B(n_793),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_734),
.B(n_813),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_810),
.B(n_801),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_772),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_SL g968 ( 
.A1(n_679),
.A2(n_812),
.B1(n_796),
.B2(n_778),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_793),
.A2(n_820),
.B(n_818),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_803),
.A2(n_818),
.B(n_804),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_803),
.A2(n_820),
.B(n_804),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_788),
.A2(n_819),
.B1(n_764),
.B2(n_752),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_766),
.A2(n_704),
.B(n_769),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_678),
.A2(n_685),
.B1(n_671),
.B2(n_594),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_677),
.B(n_683),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_675),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_677),
.B(n_683),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_675),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_751),
.A2(n_740),
.B(n_725),
.Y(n_979)
);

O2A1O1Ixp5_ASAP7_75t_SL g980 ( 
.A1(n_806),
.A2(n_579),
.B(n_636),
.C(n_540),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_707),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_979),
.A2(n_905),
.B(n_883),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_861),
.A2(n_848),
.B(n_852),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_905),
.A2(n_891),
.B(n_903),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_974),
.A2(n_980),
.B(n_865),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_865),
.A2(n_977),
.B(n_975),
.C(n_833),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_916),
.A2(n_894),
.B(n_876),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_873),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_827),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_850),
.Y(n_990)
);

NOR2x1_ASAP7_75t_SL g991 ( 
.A(n_850),
.B(n_843),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_935),
.A2(n_853),
.B(n_834),
.C(n_948),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_871),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_953),
.A2(n_893),
.B(n_971),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_955),
.B(n_929),
.Y(n_995)
);

AND2x2_ASAP7_75t_SL g996 ( 
.A(n_854),
.B(n_853),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_859),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_882),
.A2(n_886),
.B(n_878),
.C(n_854),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_848),
.A2(n_847),
.B(n_839),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_884),
.B(n_887),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_SL g1001 ( 
.A1(n_850),
.A2(n_895),
.B(n_843),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_841),
.B(n_958),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_919),
.A2(n_885),
.B(n_899),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_906),
.A2(n_837),
.B(n_926),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_842),
.A2(n_966),
.B(n_954),
.C(n_959),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_830),
.A2(n_831),
.B(n_924),
.Y(n_1006)
);

BUFx12f_ASAP7_75t_SL g1007 ( 
.A(n_866),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_840),
.A2(n_897),
.B(n_863),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_850),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_824),
.B(n_879),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_851),
.A2(n_828),
.B(n_849),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_867),
.A2(n_880),
.B(n_909),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_874),
.A2(n_914),
.B(n_924),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_969),
.A2(n_970),
.B(n_910),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_872),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_900),
.A2(n_965),
.B1(n_967),
.B2(n_856),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_981),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_955),
.B(n_940),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_874),
.A2(n_829),
.B(n_913),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_958),
.B(n_923),
.Y(n_1020)
);

AO22x1_ASAP7_75t_L g1021 ( 
.A1(n_908),
.A2(n_832),
.B1(n_965),
.B2(n_835),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_912),
.A2(n_890),
.B(n_962),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_955),
.B(n_911),
.Y(n_1023)
);

BUFx12f_ASAP7_75t_L g1024 ( 
.A(n_858),
.Y(n_1024)
);

NOR2x1_ASAP7_75t_SL g1025 ( 
.A(n_938),
.B(n_955),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_942),
.B(n_950),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_921),
.B(n_981),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_870),
.B(n_846),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_836),
.A2(n_901),
.B(n_939),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_928),
.A2(n_956),
.B(n_949),
.C(n_951),
.Y(n_1030)
);

AOI221x1_ASAP7_75t_L g1031 ( 
.A1(n_972),
.A2(n_915),
.B1(n_949),
.B2(n_973),
.C(n_945),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_868),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_931),
.A2(n_930),
.B(n_902),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_862),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_836),
.A2(n_964),
.B(n_855),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_855),
.A2(n_918),
.B(n_896),
.Y(n_1036)
);

BUFx2_ASAP7_75t_SL g1037 ( 
.A(n_888),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_907),
.A2(n_898),
.B(n_925),
.Y(n_1038)
);

O2A1O1Ixp5_ASAP7_75t_L g1039 ( 
.A1(n_941),
.A2(n_927),
.B(n_943),
.C(n_920),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_892),
.A2(n_915),
.B(n_957),
.Y(n_1040)
);

AO31x2_ASAP7_75t_L g1041 ( 
.A1(n_963),
.A2(n_946),
.A3(n_944),
.B(n_961),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_967),
.A2(n_968),
.B1(n_932),
.B2(n_888),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_921),
.B(n_857),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_857),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_907),
.A2(n_892),
.B(n_925),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_869),
.B(n_825),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_936),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_877),
.B(n_936),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_937),
.A2(n_922),
.B(n_904),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_826),
.Y(n_1050)
);

OAI22x1_ASAP7_75t_L g1051 ( 
.A1(n_976),
.A2(n_978),
.B1(n_922),
.B2(n_844),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_947),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_838),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_911),
.B(n_888),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_888),
.B(n_932),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_860),
.B(n_932),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_932),
.A2(n_864),
.B1(n_881),
.B2(n_917),
.Y(n_1057)
);

OR2x6_ASAP7_75t_L g1058 ( 
.A(n_960),
.B(n_952),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_875),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_934),
.B(n_864),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_881),
.B(n_889),
.Y(n_1061)
);

AO21x1_ASAP7_75t_L g1062 ( 
.A1(n_865),
.A2(n_974),
.B(n_906),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_861),
.A2(n_704),
.B(n_769),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_865),
.B(n_500),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_861),
.A2(n_704),
.B(n_769),
.Y(n_1065)
);

AO21x1_ASAP7_75t_L g1066 ( 
.A1(n_865),
.A2(n_974),
.B(n_906),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_871),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_981),
.Y(n_1068)
);

CKINVDCx16_ASAP7_75t_R g1069 ( 
.A(n_827),
.Y(n_1069)
);

O2A1O1Ixp5_ASAP7_75t_L g1070 ( 
.A1(n_865),
.A2(n_678),
.B(n_886),
.C(n_845),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_871),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_974),
.A2(n_678),
.B(n_980),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_979),
.A2(n_905),
.B(n_883),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_L g1074 ( 
.A1(n_865),
.A2(n_678),
.B(n_886),
.C(n_845),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_975),
.B(n_977),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_865),
.B(n_500),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_974),
.A2(n_678),
.B(n_980),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_859),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_871),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_850),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_975),
.B(n_977),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_975),
.B(n_977),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_866),
.B(n_500),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_845),
.A2(n_678),
.A3(n_672),
.B(n_933),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_979),
.A2(n_905),
.B(n_883),
.Y(n_1085)
);

AOI21x1_ASAP7_75t_L g1086 ( 
.A1(n_924),
.A2(n_744),
.B(n_919),
.Y(n_1086)
);

AO31x2_ASAP7_75t_L g1087 ( 
.A1(n_845),
.A2(n_678),
.A3(n_672),
.B(n_933),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_974),
.A2(n_678),
.B(n_980),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_974),
.A2(n_678),
.B(n_980),
.Y(n_1089)
);

AOI21x1_ASAP7_75t_L g1090 ( 
.A1(n_924),
.A2(n_744),
.B(n_919),
.Y(n_1090)
);

AOI21xp33_ASAP7_75t_L g1091 ( 
.A1(n_865),
.A2(n_974),
.B(n_966),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_861),
.A2(n_704),
.B(n_769),
.Y(n_1092)
);

INVx8_ASAP7_75t_L g1093 ( 
.A(n_850),
.Y(n_1093)
);

NAND2x1_ASAP7_75t_L g1094 ( 
.A(n_843),
.B(n_699),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_850),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_979),
.A2(n_905),
.B(n_883),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_871),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_SL g1098 ( 
.A1(n_933),
.A2(n_948),
.B(n_973),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_894),
.A2(n_903),
.B(n_876),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_861),
.A2(n_704),
.B(n_769),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_979),
.A2(n_905),
.B(n_883),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_975),
.B(n_977),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_865),
.B(n_500),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_974),
.A2(n_678),
.B(n_980),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_871),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_975),
.B(n_977),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_894),
.A2(n_903),
.B(n_876),
.Y(n_1107)
);

O2A1O1Ixp5_ASAP7_75t_L g1108 ( 
.A1(n_865),
.A2(n_678),
.B(n_886),
.C(n_845),
.Y(n_1108)
);

AOI21xp33_ASAP7_75t_L g1109 ( 
.A1(n_865),
.A2(n_974),
.B(n_966),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_873),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_894),
.A2(n_903),
.B(n_876),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_866),
.B(n_500),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_845),
.A2(n_678),
.A3(n_672),
.B(n_933),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_975),
.B(n_977),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_871),
.Y(n_1115)
);

OAI22x1_ASAP7_75t_L g1116 ( 
.A1(n_966),
.A2(n_865),
.B1(n_797),
.B2(n_801),
.Y(n_1116)
);

BUFx10_ASAP7_75t_L g1117 ( 
.A(n_1060),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1083),
.B(n_1112),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1017),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_996),
.A2(n_1102),
.B1(n_1106),
.B2(n_1114),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_1093),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_989),
.Y(n_1122)
);

CKINVDCx6p67_ASAP7_75t_R g1123 ( 
.A(n_1069),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_1017),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_989),
.Y(n_1125)
);

AO21x2_ASAP7_75t_L g1126 ( 
.A1(n_985),
.A2(n_1077),
.B(n_1072),
.Y(n_1126)
);

INVx5_ASAP7_75t_L g1127 ( 
.A(n_1093),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_993),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1060),
.B(n_1053),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1010),
.B(n_1064),
.Y(n_1130)
);

OR2x2_ASAP7_75t_L g1131 ( 
.A(n_1000),
.B(n_1020),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1067),
.Y(n_1132)
);

CKINVDCx8_ASAP7_75t_R g1133 ( 
.A(n_1037),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_1032),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_SL g1135 ( 
.A(n_996),
.B(n_1005),
.Y(n_1135)
);

BUFx10_ASAP7_75t_L g1136 ( 
.A(n_1060),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_1054),
.B(n_995),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1095),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_997),
.B(n_1078),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_1095),
.B(n_995),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_995),
.B(n_1018),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_983),
.A2(n_1065),
.B(n_1063),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1095),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1064),
.B(n_1076),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1076),
.B(n_1103),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_1093),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_SL g1147 ( 
.A1(n_992),
.A2(n_998),
.B(n_986),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1024),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1092),
.A2(n_1100),
.B(n_999),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1018),
.B(n_1015),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_1018),
.B(n_1043),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1002),
.B(n_1026),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1027),
.B(n_1048),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1005),
.A2(n_1030),
.B1(n_1023),
.B2(n_1028),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_1047),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1016),
.A2(n_1021),
.B1(n_1023),
.B2(n_1042),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1011),
.A2(n_1008),
.B(n_1029),
.Y(n_1157)
);

AOI222xp33_ASAP7_75t_L g1158 ( 
.A1(n_1030),
.A2(n_1079),
.B1(n_1071),
.B2(n_1105),
.C1(n_1097),
.C2(n_1115),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1034),
.B(n_1046),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1050),
.B(n_1051),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1068),
.B(n_1044),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1068),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1044),
.B(n_1056),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1012),
.A2(n_1013),
.B(n_1001),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1088),
.A2(n_1089),
.B1(n_1104),
.B2(n_1058),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_988),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_1007),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1019),
.A2(n_1025),
.B(n_1108),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_1024),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1110),
.B(n_1058),
.Y(n_1170)
);

INVx5_ASAP7_75t_L g1171 ( 
.A(n_990),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1057),
.B(n_1055),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1058),
.A2(n_1040),
.B1(n_1045),
.B2(n_1052),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_R g1174 ( 
.A(n_1061),
.B(n_1080),
.Y(n_1174)
);

BUFx4f_ASAP7_75t_SL g1175 ( 
.A(n_1059),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_990),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1084),
.B(n_1087),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1055),
.Y(n_1178)
);

AO21x2_ASAP7_75t_L g1179 ( 
.A1(n_1098),
.A2(n_982),
.B(n_1101),
.Y(n_1179)
);

AND2x6_ASAP7_75t_L g1180 ( 
.A(n_1009),
.B(n_1080),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1070),
.A2(n_1108),
.B(n_1074),
.Y(n_1181)
);

BUFx4_ASAP7_75t_SL g1182 ( 
.A(n_991),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1084),
.B(n_1113),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1084),
.B(n_1113),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1084),
.B(n_1113),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1031),
.B(n_1035),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1087),
.B(n_1113),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_1094),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1087),
.B(n_1041),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1038),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1006),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1022),
.B(n_1036),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_984),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_994),
.A2(n_1039),
.B(n_1101),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1003),
.B(n_1014),
.Y(n_1195)
);

BUFx12f_ASAP7_75t_L g1196 ( 
.A(n_1033),
.Y(n_1196)
);

OR2x2_ASAP7_75t_SL g1197 ( 
.A(n_1033),
.B(n_982),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1073),
.A2(n_1085),
.B(n_1096),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1014),
.A2(n_1085),
.B1(n_1096),
.B2(n_987),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1064),
.B(n_1076),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1075),
.B(n_1081),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1004),
.A2(n_704),
.B(n_699),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_989),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_SL g1204 ( 
.A1(n_992),
.A2(n_678),
.B(n_1005),
.C(n_986),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1075),
.B(n_1081),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1064),
.B(n_1076),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1060),
.B(n_1053),
.Y(n_1207)
);

AOI21xp33_ASAP7_75t_L g1208 ( 
.A1(n_1091),
.A2(n_865),
.B(n_1109),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_989),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1017),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1083),
.B(n_1112),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1091),
.A2(n_865),
.B1(n_1109),
.B2(n_1116),
.Y(n_1212)
);

INVxp67_ASAP7_75t_L g1213 ( 
.A(n_1017),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1017),
.Y(n_1214)
);

CKINVDCx11_ASAP7_75t_R g1215 ( 
.A(n_1059),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1075),
.B(n_1081),
.Y(n_1216)
);

NOR2x1p5_ASAP7_75t_SL g1217 ( 
.A(n_1086),
.B(n_830),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_SL g1218 ( 
.A1(n_985),
.A2(n_865),
.B(n_842),
.C(n_832),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_993),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_989),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_989),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1062),
.A2(n_1066),
.A3(n_992),
.B(n_1031),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1091),
.A2(n_865),
.B1(n_1109),
.B2(n_1116),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_996),
.A2(n_1075),
.B1(n_1082),
.B2(n_1081),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_996),
.A2(n_1075),
.B1(n_1082),
.B2(n_1081),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1004),
.A2(n_704),
.B(n_699),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1075),
.B(n_1081),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_993),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_993),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1075),
.B(n_1081),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1004),
.A2(n_704),
.B(n_699),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_989),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1049),
.A2(n_1090),
.B(n_1086),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1095),
.Y(n_1234)
);

INVx1_ASAP7_75t_SL g1235 ( 
.A(n_997),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_989),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1083),
.B(n_1112),
.Y(n_1237)
);

BUFx12f_ASAP7_75t_L g1238 ( 
.A(n_1024),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1099),
.A2(n_1111),
.B(n_1107),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1017),
.Y(n_1240)
);

CKINVDCx6p67_ASAP7_75t_R g1241 ( 
.A(n_1069),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_SL g1242 ( 
.A(n_989),
.Y(n_1242)
);

CKINVDCx8_ASAP7_75t_R g1243 ( 
.A(n_1069),
.Y(n_1243)
);

INVx2_ASAP7_75t_SL g1244 ( 
.A(n_989),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_993),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1137),
.B(n_1141),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1139),
.Y(n_1247)
);

AOI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1233),
.A2(n_1198),
.B(n_1194),
.Y(n_1248)
);

CKINVDCx11_ASAP7_75t_R g1249 ( 
.A(n_1215),
.Y(n_1249)
);

CKINVDCx11_ASAP7_75t_R g1250 ( 
.A(n_1243),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_SL g1251 ( 
.A(n_1220),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1200),
.A2(n_1206),
.B1(n_1208),
.B2(n_1212),
.Y(n_1252)
);

CKINVDCx6p67_ASAP7_75t_R g1253 ( 
.A(n_1242),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1239),
.A2(n_1164),
.B(n_1149),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_1227),
.Y(n_1255)
);

NAND2x1p5_ASAP7_75t_L g1256 ( 
.A(n_1170),
.B(n_1172),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1166),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1230),
.B(n_1201),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_1235),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1235),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1221),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1130),
.B(n_1135),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1201),
.A2(n_1205),
.B1(n_1216),
.B2(n_1144),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1205),
.B(n_1216),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1128),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1208),
.A2(n_1223),
.B1(n_1145),
.B2(n_1135),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1132),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1162),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1196),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1161),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1120),
.B(n_1224),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1219),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1228),
.Y(n_1273)
);

OA21x2_ASAP7_75t_L g1274 ( 
.A1(n_1157),
.A2(n_1181),
.B(n_1192),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1119),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1236),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1229),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1193),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1124),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1168),
.A2(n_1142),
.B(n_1199),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1156),
.A2(n_1152),
.B1(n_1131),
.B2(n_1120),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1210),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1224),
.B(n_1225),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1245),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1122),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1214),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1141),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1159),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_1240),
.Y(n_1289)
);

BUFx2_ASAP7_75t_R g1290 ( 
.A(n_1148),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1238),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1225),
.B(n_1137),
.Y(n_1292)
);

BUFx4f_ASAP7_75t_SL g1293 ( 
.A(n_1123),
.Y(n_1293)
);

NAND2x1p5_ASAP7_75t_L g1294 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1163),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1118),
.A2(n_1211),
.B1(n_1237),
.B2(n_1165),
.Y(n_1296)
);

OAI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1160),
.A2(n_1241),
.B1(n_1154),
.B2(n_1167),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1180),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1154),
.A2(n_1165),
.B1(n_1153),
.B2(n_1173),
.Y(n_1299)
);

BUFx8_ASAP7_75t_L g1300 ( 
.A(n_1242),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1151),
.B(n_1213),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1155),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1209),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1173),
.A2(n_1117),
.B1(n_1136),
.B2(n_1151),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1178),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1127),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1222),
.B(n_1189),
.Y(n_1307)
);

INVxp33_ASAP7_75t_L g1308 ( 
.A(n_1155),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1129),
.B(n_1207),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1175),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1176),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1158),
.B(n_1183),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1127),
.Y(n_1313)
);

AO21x1_ASAP7_75t_SL g1314 ( 
.A1(n_1189),
.A2(n_1184),
.B(n_1187),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1158),
.B(n_1126),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1129),
.B(n_1207),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1179),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1179),
.Y(n_1318)
);

AO21x1_ASAP7_75t_L g1319 ( 
.A1(n_1186),
.A2(n_1184),
.B(n_1177),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1155),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1232),
.Y(n_1321)
);

BUFx4_ASAP7_75t_R g1322 ( 
.A(n_1136),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1186),
.A2(n_1150),
.B1(n_1134),
.B2(n_1174),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_1125),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1218),
.A2(n_1147),
.B(n_1204),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1222),
.Y(n_1326)
);

CKINVDCx11_ASAP7_75t_R g1327 ( 
.A(n_1169),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1202),
.A2(n_1226),
.B(n_1231),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1138),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1222),
.B(n_1187),
.Y(n_1330)
);

OR2x6_ASAP7_75t_L g1331 ( 
.A(n_1190),
.B(n_1217),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1197),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1195),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1150),
.A2(n_1185),
.B1(n_1140),
.B2(n_1244),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1138),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1140),
.B(n_1171),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1133),
.A2(n_1203),
.B1(n_1188),
.B2(n_1127),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1143),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1182),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1143),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1140),
.A2(n_1188),
.B1(n_1127),
.B2(n_1180),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1143),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1234),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1180),
.A2(n_1140),
.B(n_1171),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1146),
.Y(n_1345)
);

CKINVDCx11_ASAP7_75t_R g1346 ( 
.A(n_1146),
.Y(n_1346)
);

AO21x1_ASAP7_75t_L g1347 ( 
.A1(n_1121),
.A2(n_1171),
.B(n_1234),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1234),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1171),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1146),
.B(n_1227),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1170),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1200),
.A2(n_865),
.B(n_1091),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1139),
.Y(n_1353)
);

AOI222xp33_ASAP7_75t_L g1354 ( 
.A1(n_1200),
.A2(n_1206),
.B1(n_966),
.B2(n_1116),
.C1(n_865),
.C2(n_748),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1137),
.B(n_1141),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1200),
.A2(n_865),
.B1(n_1206),
.B2(n_1109),
.Y(n_1356)
);

AOI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1233),
.A2(n_1198),
.B(n_1194),
.Y(n_1357)
);

INVx4_ASAP7_75t_L g1358 ( 
.A(n_1127),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1141),
.Y(n_1359)
);

BUFx2_ASAP7_75t_R g1360 ( 
.A(n_1243),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1222),
.B(n_1189),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1128),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1128),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1200),
.A2(n_1206),
.B1(n_865),
.B2(n_842),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1170),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1128),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1200),
.A2(n_1206),
.B1(n_1230),
.B2(n_1227),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1128),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1227),
.B(n_1230),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1200),
.A2(n_865),
.B1(n_1206),
.B2(n_1109),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1141),
.Y(n_1371)
);

BUFx12f_ASAP7_75t_L g1372 ( 
.A(n_1215),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1312),
.B(n_1271),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1268),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1328),
.B(n_1256),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1278),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1312),
.B(n_1271),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1269),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1248),
.A2(n_1357),
.B(n_1254),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1268),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1283),
.B(n_1315),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1286),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1319),
.A2(n_1326),
.A3(n_1318),
.B(n_1317),
.Y(n_1383)
);

OAI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1352),
.A2(n_1367),
.B1(n_1369),
.B2(n_1258),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1319),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1307),
.B(n_1361),
.Y(n_1386)
);

INVx4_ASAP7_75t_SL g1387 ( 
.A(n_1331),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1286),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1275),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1307),
.B(n_1361),
.Y(n_1390)
);

AO21x1_ASAP7_75t_L g1391 ( 
.A1(n_1297),
.A2(n_1325),
.B(n_1281),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1285),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1333),
.B(n_1332),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1279),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1255),
.B(n_1263),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1330),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1330),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1256),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1331),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1256),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1283),
.B(n_1315),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1294),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1285),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1351),
.B(n_1365),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1264),
.B(n_1356),
.Y(n_1405)
);

AOI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1274),
.A2(n_1331),
.B(n_1280),
.Y(n_1406)
);

BUFx8_ASAP7_75t_L g1407 ( 
.A(n_1372),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1370),
.B(n_1364),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1252),
.A2(n_1354),
.B(n_1266),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1292),
.B(n_1351),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1365),
.B(n_1292),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1294),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1269),
.B(n_1257),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1247),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1282),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1270),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1262),
.B(n_1296),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1269),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1259),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1265),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1311),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1262),
.B(n_1299),
.Y(n_1422)
);

AO21x1_ASAP7_75t_SL g1423 ( 
.A1(n_1334),
.A2(n_1323),
.B(n_1295),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1344),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1267),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1272),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1273),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_SL g1428 ( 
.A(n_1313),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1277),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1284),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1362),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1363),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1347),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1366),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1336),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1368),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1353),
.B(n_1288),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1305),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1314),
.B(n_1316),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1321),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1349),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1314),
.B(n_1316),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1260),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1289),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1298),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1350),
.A2(n_1335),
.B(n_1329),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1301),
.B(n_1302),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1298),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1321),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1309),
.B(n_1316),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1298),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1303),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1309),
.B(n_1359),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1304),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1405),
.B(n_1360),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1386),
.B(n_1320),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1386),
.B(n_1337),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1409),
.A2(n_1309),
.B1(n_1371),
.B2(n_1287),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1384),
.B(n_1308),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1399),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1381),
.B(n_1308),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1399),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1395),
.B(n_1324),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1382),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1382),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1407),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1391),
.A2(n_1287),
.B1(n_1371),
.B2(n_1359),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1391),
.A2(n_1287),
.B1(n_1371),
.B2(n_1359),
.Y(n_1468)
);

NOR2x1_ASAP7_75t_L g1469 ( 
.A(n_1433),
.B(n_1313),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1388),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1424),
.B(n_1393),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1390),
.B(n_1340),
.Y(n_1472)
);

INVx1_ASAP7_75t_SL g1473 ( 
.A(n_1443),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1414),
.B(n_1348),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1376),
.Y(n_1475)
);

NAND2x1p5_ASAP7_75t_L g1476 ( 
.A(n_1433),
.B(n_1336),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1381),
.B(n_1371),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1401),
.B(n_1371),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1376),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1424),
.B(n_1306),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1401),
.B(n_1359),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1388),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1374),
.Y(n_1483)
);

NOR2x2_ASAP7_75t_L g1484 ( 
.A(n_1438),
.B(n_1407),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1389),
.B(n_1394),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1408),
.A2(n_1253),
.B1(n_1303),
.B2(n_1287),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1390),
.B(n_1338),
.Y(n_1487)
);

INVx3_ASAP7_75t_SL g1488 ( 
.A(n_1387),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1396),
.B(n_1342),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1397),
.B(n_1343),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1397),
.B(n_1246),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1379),
.A2(n_1306),
.B(n_1345),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1373),
.B(n_1246),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1402),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1373),
.B(n_1246),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1377),
.B(n_1355),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1377),
.B(n_1355),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1415),
.B(n_1355),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1385),
.B(n_1253),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1407),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1433),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1424),
.B(n_1358),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1420),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1411),
.B(n_1341),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1420),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1380),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1437),
.B(n_1261),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1385),
.B(n_1276),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1411),
.B(n_1358),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1437),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1510),
.B(n_1416),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_L g1512 ( 
.A(n_1459),
.B(n_1454),
.C(n_1419),
.Y(n_1512)
);

NAND4xp25_ASAP7_75t_L g1513 ( 
.A(n_1463),
.B(n_1454),
.C(n_1447),
.D(n_1438),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1486),
.B(n_1413),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1485),
.B(n_1421),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1458),
.A2(n_1417),
.B1(n_1422),
.B2(n_1403),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1467),
.A2(n_1468),
.B1(n_1455),
.B2(n_1499),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1483),
.B(n_1404),
.Y(n_1518)
);

NAND3xp33_ASAP7_75t_L g1519 ( 
.A(n_1499),
.B(n_1444),
.C(n_1447),
.Y(n_1519)
);

NAND4xp25_ASAP7_75t_SL g1520 ( 
.A(n_1504),
.B(n_1422),
.C(n_1339),
.D(n_1417),
.Y(n_1520)
);

OAI21xp33_ASAP7_75t_L g1521 ( 
.A1(n_1507),
.A2(n_1434),
.B(n_1430),
.Y(n_1521)
);

NAND4xp25_ASAP7_75t_L g1522 ( 
.A(n_1474),
.B(n_1431),
.C(n_1430),
.D(n_1429),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1461),
.A2(n_1423),
.B1(n_1398),
.B2(n_1400),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1471),
.B(n_1410),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1506),
.B(n_1456),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1456),
.B(n_1404),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1471),
.B(n_1477),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1508),
.B(n_1413),
.C(n_1441),
.Y(n_1528)
);

AOI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1473),
.A2(n_1413),
.B1(n_1434),
.B2(n_1425),
.C(n_1427),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1461),
.B(n_1436),
.Y(n_1530)
);

OAI21xp33_ASAP7_75t_L g1531 ( 
.A1(n_1457),
.A2(n_1432),
.B(n_1431),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1471),
.B(n_1410),
.Y(n_1532)
);

OAI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1498),
.A2(n_1452),
.B1(n_1403),
.B2(n_1449),
.C(n_1392),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1501),
.A2(n_1423),
.B1(n_1398),
.B2(n_1400),
.Y(n_1534)
);

NAND3xp33_ASAP7_75t_L g1535 ( 
.A(n_1508),
.B(n_1413),
.C(n_1451),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1472),
.B(n_1436),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1466),
.B(n_1452),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1471),
.B(n_1410),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1472),
.B(n_1425),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1478),
.B(n_1439),
.Y(n_1540)
);

OAI21xp33_ASAP7_75t_L g1541 ( 
.A1(n_1457),
.A2(n_1429),
.B(n_1427),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1487),
.B(n_1426),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1478),
.B(n_1439),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1481),
.B(n_1442),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1487),
.B(n_1426),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1464),
.B(n_1432),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1465),
.B(n_1446),
.Y(n_1547)
);

NAND3xp33_ASAP7_75t_L g1548 ( 
.A(n_1469),
.B(n_1445),
.C(n_1448),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1501),
.A2(n_1442),
.B1(n_1504),
.B2(n_1450),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1494),
.B(n_1383),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1501),
.A2(n_1407),
.B1(n_1428),
.B2(n_1450),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1475),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1500),
.A2(n_1392),
.B1(n_1449),
.B2(n_1440),
.Y(n_1553)
);

NOR3xp33_ASAP7_75t_SL g1554 ( 
.A(n_1503),
.B(n_1310),
.C(n_1412),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1470),
.B(n_1446),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1481),
.A2(n_1453),
.B1(n_1375),
.B2(n_1435),
.Y(n_1556)
);

NOR3xp33_ASAP7_75t_L g1557 ( 
.A(n_1469),
.B(n_1440),
.C(n_1327),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1482),
.B(n_1446),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1490),
.B(n_1446),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1490),
.B(n_1393),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1491),
.B(n_1509),
.Y(n_1561)
);

OAI221xp5_ASAP7_75t_L g1562 ( 
.A1(n_1476),
.A2(n_1378),
.B1(n_1418),
.B2(n_1375),
.C(n_1261),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1491),
.B(n_1393),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1493),
.B(n_1250),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1480),
.A2(n_1451),
.B(n_1448),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1559),
.B(n_1494),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1552),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1562),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1547),
.B(n_1475),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1552),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1550),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1527),
.B(n_1561),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1550),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1555),
.Y(n_1574)
);

INVxp67_ASAP7_75t_L g1575 ( 
.A(n_1558),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1539),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1525),
.B(n_1479),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1542),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1512),
.B(n_1519),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1545),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1536),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1540),
.B(n_1492),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1543),
.B(n_1492),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1546),
.B(n_1479),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1565),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1512),
.A2(n_1497),
.B1(n_1495),
.B2(n_1496),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1530),
.Y(n_1587)
);

INVxp67_ASAP7_75t_SL g1588 ( 
.A(n_1519),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1544),
.B(n_1406),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1528),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1528),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1524),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1548),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1532),
.B(n_1502),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1521),
.B(n_1503),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1538),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1544),
.B(n_1406),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1518),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_SL g1599 ( 
.A(n_1557),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1535),
.B(n_1502),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1588),
.B(n_1526),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1588),
.B(n_1515),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1599),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1599),
.A2(n_1534),
.B1(n_1523),
.B2(n_1554),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1593),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1594),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1577),
.Y(n_1607)
);

INVx4_ASAP7_75t_L g1608 ( 
.A(n_1568),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1577),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1577),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1592),
.B(n_1556),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1576),
.B(n_1511),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1598),
.B(n_1560),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1590),
.B(n_1522),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1590),
.B(n_1563),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1590),
.B(n_1591),
.Y(n_1616)
);

NOR2x1_ASAP7_75t_L g1617 ( 
.A(n_1579),
.B(n_1513),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1570),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1591),
.B(n_1531),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1584),
.Y(n_1620)
);

NAND2x1p5_ASAP7_75t_SL g1621 ( 
.A(n_1579),
.B(n_1514),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1591),
.B(n_1531),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1584),
.Y(n_1623)
);

INVxp67_ASAP7_75t_SL g1624 ( 
.A(n_1593),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1566),
.B(n_1541),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1570),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1584),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1585),
.A2(n_1520),
.B(n_1517),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1592),
.B(n_1460),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1568),
.B(n_1551),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1576),
.B(n_1529),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1567),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1592),
.B(n_1596),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1566),
.B(n_1541),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1567),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1566),
.B(n_1489),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1570),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1592),
.B(n_1460),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1596),
.B(n_1460),
.Y(n_1639)
);

NAND4xp25_ASAP7_75t_L g1640 ( 
.A(n_1568),
.B(n_1533),
.C(n_1549),
.D(n_1516),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1567),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1596),
.B(n_1462),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1596),
.B(n_1462),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1576),
.B(n_1505),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1632),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1619),
.B(n_1593),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1611),
.B(n_1606),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1605),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1619),
.B(n_1575),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_1603),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1635),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1641),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1644),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1636),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1636),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1623),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1617),
.B(n_1585),
.Y(n_1657)
);

INVxp67_ASAP7_75t_SL g1658 ( 
.A(n_1624),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1618),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1627),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1631),
.B(n_1585),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1606),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1614),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1611),
.B(n_1582),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1628),
.A2(n_1586),
.B(n_1564),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1620),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1620),
.Y(n_1667)
);

AND3x1_ASAP7_75t_L g1668 ( 
.A(n_1602),
.B(n_1537),
.C(n_1586),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1614),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1607),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1616),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1608),
.B(n_1568),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1606),
.B(n_1582),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1608),
.B(n_1598),
.Y(n_1674)
);

NOR2xp67_ASAP7_75t_L g1675 ( 
.A(n_1608),
.B(n_1575),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1609),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1618),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1629),
.B(n_1582),
.Y(n_1678)
);

OAI21xp33_ASAP7_75t_L g1679 ( 
.A1(n_1640),
.A2(n_1586),
.B(n_1574),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1630),
.Y(n_1680)
);

NOR4xp25_ASAP7_75t_L g1681 ( 
.A(n_1630),
.B(n_1574),
.C(n_1578),
.D(n_1580),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1622),
.B(n_1574),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_1622),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1610),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1629),
.B(n_1583),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1626),
.Y(n_1686)
);

NAND2xp33_ASAP7_75t_SL g1687 ( 
.A(n_1621),
.B(n_1488),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1616),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1625),
.B(n_1634),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1638),
.B(n_1583),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1671),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1650),
.B(n_1372),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_SL g1693 ( 
.A(n_1680),
.B(n_1290),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1651),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1673),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1689),
.B(n_1621),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1679),
.A2(n_1604),
.B1(n_1601),
.B2(n_1615),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1651),
.Y(n_1698)
);

NOR3xp33_ASAP7_75t_SL g1699 ( 
.A(n_1687),
.B(n_1310),
.C(n_1553),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1669),
.B(n_1615),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1665),
.A2(n_1634),
.B(n_1625),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1647),
.B(n_1638),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1663),
.B(n_1612),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1672),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1647),
.B(n_1639),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1664),
.B(n_1639),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1661),
.B(n_1571),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1683),
.B(n_1571),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1673),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1648),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1658),
.Y(n_1711)
);

AOI222xp33_ASAP7_75t_L g1712 ( 
.A1(n_1657),
.A2(n_1300),
.B1(n_1293),
.B2(n_1250),
.C1(n_1327),
.C2(n_1249),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1652),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1664),
.B(n_1642),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1689),
.B(n_1613),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1675),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1688),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1646),
.B(n_1569),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1681),
.B(n_1572),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1652),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1645),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1646),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1668),
.B(n_1626),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1654),
.B(n_1642),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1654),
.B(n_1643),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1656),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1656),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1717),
.B(n_1674),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_SL g1729 ( 
.A1(n_1723),
.A2(n_1251),
.B(n_1249),
.Y(n_1729)
);

AND2x2_ASAP7_75t_SL g1730 ( 
.A(n_1723),
.B(n_1649),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1717),
.Y(n_1731)
);

AOI321xp33_ASAP7_75t_L g1732 ( 
.A1(n_1723),
.A2(n_1697),
.A3(n_1696),
.B1(n_1719),
.B2(n_1703),
.C(n_1700),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1723),
.B(n_1649),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1696),
.B(n_1655),
.Y(n_1734)
);

OAI211xp5_ASAP7_75t_L g1735 ( 
.A1(n_1701),
.A2(n_1667),
.B(n_1666),
.C(n_1655),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1715),
.B(n_1682),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1710),
.B(n_1653),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1701),
.A2(n_1682),
.B1(n_1667),
.B2(n_1666),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1691),
.Y(n_1739)
);

AOI21xp33_ASAP7_75t_L g1740 ( 
.A1(n_1711),
.A2(n_1670),
.B(n_1660),
.Y(n_1740)
);

OAI21xp33_ASAP7_75t_L g1741 ( 
.A1(n_1704),
.A2(n_1653),
.B(n_1660),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1704),
.B(n_1670),
.Y(n_1742)
);

AOI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1722),
.A2(n_1684),
.B1(n_1676),
.B2(n_1686),
.C(n_1662),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1699),
.A2(n_1600),
.B1(n_1676),
.B2(n_1684),
.Y(n_1744)
);

O2A1O1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1716),
.A2(n_1662),
.B(n_1686),
.C(n_1659),
.Y(n_1745)
);

OAI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1693),
.A2(n_1677),
.B1(n_1659),
.B2(n_1685),
.C(n_1678),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1694),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1702),
.B(n_1678),
.Y(n_1748)
);

AO22x1_ASAP7_75t_L g1749 ( 
.A1(n_1722),
.A2(n_1300),
.B1(n_1685),
.B2(n_1690),
.Y(n_1749)
);

OAI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1693),
.A2(n_1677),
.B(n_1595),
.Y(n_1750)
);

O2A1O1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1704),
.A2(n_1712),
.B(n_1692),
.C(n_1721),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1712),
.B(n_1690),
.Y(n_1752)
);

AOI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1721),
.A2(n_1580),
.B1(n_1578),
.B2(n_1581),
.C(n_1587),
.Y(n_1753)
);

AOI211xp5_ASAP7_75t_SL g1754 ( 
.A1(n_1715),
.A2(n_1600),
.B(n_1595),
.C(n_1643),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1730),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1730),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1747),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1731),
.B(n_1702),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1739),
.B(n_1705),
.Y(n_1759)
);

NAND2x1_ASAP7_75t_L g1760 ( 
.A(n_1729),
.B(n_1726),
.Y(n_1760)
);

NAND2xp33_ASAP7_75t_L g1761 ( 
.A(n_1733),
.B(n_1726),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1752),
.B(n_1705),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1751),
.B(n_1291),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1736),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1733),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1734),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1728),
.B(n_1724),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1742),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1737),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1741),
.B(n_1724),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1748),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1738),
.B(n_1725),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1750),
.B(n_1725),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1729),
.B(n_1727),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1754),
.B(n_1706),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1756),
.B(n_1743),
.Y(n_1776)
);

AOI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1761),
.A2(n_1740),
.B1(n_1735),
.B2(n_1745),
.C(n_1732),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1766),
.Y(n_1778)
);

AOI211x1_ASAP7_75t_SL g1779 ( 
.A1(n_1762),
.A2(n_1744),
.B(n_1709),
.C(n_1695),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_R g1780 ( 
.A(n_1756),
.B(n_1291),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_1774),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1763),
.B(n_1760),
.Y(n_1782)
);

NAND4xp75_ASAP7_75t_SL g1783 ( 
.A(n_1775),
.B(n_1749),
.C(n_1706),
.D(n_1714),
.Y(n_1783)
);

AOI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1761),
.A2(n_1746),
.B1(n_1727),
.B2(n_1698),
.C(n_1720),
.Y(n_1784)
);

AOI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1760),
.A2(n_1708),
.B(n_1698),
.Y(n_1785)
);

AOI21xp33_ASAP7_75t_L g1786 ( 
.A1(n_1755),
.A2(n_1713),
.B(n_1694),
.Y(n_1786)
);

OAI21xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1755),
.A2(n_1708),
.B(n_1714),
.Y(n_1787)
);

AOI211xp5_ASAP7_75t_L g1788 ( 
.A1(n_1765),
.A2(n_1720),
.B(n_1713),
.C(n_1707),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1777),
.B(n_1765),
.Y(n_1789)
);

NOR3xp33_ASAP7_75t_L g1790 ( 
.A(n_1782),
.B(n_1769),
.C(n_1768),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1778),
.Y(n_1791)
);

NOR2x1_ASAP7_75t_L g1792 ( 
.A(n_1783),
.B(n_1758),
.Y(n_1792)
);

NOR2x1_ASAP7_75t_L g1793 ( 
.A(n_1776),
.B(n_1757),
.Y(n_1793)
);

O2A1O1Ixp33_ASAP7_75t_L g1794 ( 
.A1(n_1781),
.A2(n_1772),
.B(n_1770),
.C(n_1764),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1784),
.B(n_1759),
.C(n_1775),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1785),
.B(n_1771),
.Y(n_1796)
);

NOR3xp33_ASAP7_75t_SL g1797 ( 
.A(n_1787),
.B(n_1767),
.C(n_1707),
.Y(n_1797)
);

INVx4_ASAP7_75t_L g1798 ( 
.A(n_1780),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1788),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1786),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1796),
.B(n_1779),
.Y(n_1801)
);

NOR3xp33_ASAP7_75t_L g1802 ( 
.A(n_1798),
.B(n_1773),
.C(n_1709),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1796),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1789),
.A2(n_1773),
.B(n_1753),
.Y(n_1804)
);

NOR2x1_ASAP7_75t_L g1805 ( 
.A(n_1793),
.B(n_1276),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1795),
.B(n_1300),
.C(n_1695),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1803),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1805),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1801),
.Y(n_1809)
);

NOR2x1_ASAP7_75t_L g1810 ( 
.A(n_1806),
.B(n_1791),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1802),
.A2(n_1792),
.B1(n_1799),
.B2(n_1790),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1804),
.A2(n_1800),
.B1(n_1797),
.B2(n_1709),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1807),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1810),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1808),
.B(n_1695),
.Y(n_1815)
);

INVxp67_ASAP7_75t_L g1816 ( 
.A(n_1811),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1812),
.B(n_1794),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1814),
.B(n_1809),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1815),
.Y(n_1819)
);

NAND4xp75_ASAP7_75t_L g1820 ( 
.A(n_1817),
.B(n_1346),
.C(n_1251),
.D(n_1589),
.Y(n_1820)
);

AOI22x1_ASAP7_75t_L g1821 ( 
.A1(n_1819),
.A2(n_1813),
.B1(n_1816),
.B2(n_1815),
.Y(n_1821)
);

NOR2x1p5_ASAP7_75t_L g1822 ( 
.A(n_1821),
.B(n_1820),
.Y(n_1822)
);

AO22x2_ASAP7_75t_L g1823 ( 
.A1(n_1822),
.A2(n_1818),
.B1(n_1718),
.B2(n_1637),
.Y(n_1823)
);

OAI21xp33_ASAP7_75t_L g1824 ( 
.A1(n_1822),
.A2(n_1718),
.B(n_1418),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1823),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1824),
.B(n_1637),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_SL g1827 ( 
.A(n_1825),
.B(n_1251),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1826),
.A2(n_1633),
.B1(n_1418),
.B2(n_1378),
.Y(n_1828)
);

OAI222xp33_ASAP7_75t_L g1829 ( 
.A1(n_1828),
.A2(n_1346),
.B1(n_1573),
.B2(n_1571),
.C1(n_1633),
.C2(n_1569),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1829),
.Y(n_1830)
);

OAI221xp5_ASAP7_75t_R g1831 ( 
.A1(n_1830),
.A2(n_1827),
.B1(n_1322),
.B2(n_1484),
.C(n_1573),
.Y(n_1831)
);

AOI211xp5_ASAP7_75t_L g1832 ( 
.A1(n_1831),
.A2(n_1488),
.B(n_1569),
.C(n_1597),
.Y(n_1832)
);


endmodule