module real_jpeg_13511_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_1),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_1),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_84)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_3),
.A2(n_29),
.B1(n_36),
.B2(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_3),
.A2(n_53),
.B1(n_60),
.B2(n_63),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_5),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_5),
.A2(n_60),
.B1(n_63),
.B2(n_68),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_68),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_5),
.A2(n_29),
.B1(n_36),
.B2(n_68),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_7),
.A2(n_29),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_7),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_8),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_8),
.A2(n_60),
.B1(n_63),
.B2(n_101),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_101),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_8),
.A2(n_29),
.B1(n_36),
.B2(n_101),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_9),
.A2(n_65),
.B(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_9),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_9),
.B(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_9),
.B(n_63),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_135),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_9),
.A2(n_44),
.B(n_49),
.C(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_9),
.B(n_109),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_9),
.B(n_33),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_9),
.B(n_54),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g240 ( 
.A1(n_9),
.A2(n_63),
.B(n_190),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_10),
.A2(n_65),
.B1(n_66),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_10),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_10),
.A2(n_60),
.B1(n_63),
.B2(n_137),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_137),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_10),
.A2(n_29),
.B1(n_36),
.B2(n_137),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_14),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_14),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_14),
.A2(n_60),
.B1(n_63),
.B2(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_70),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_14),
.A2(n_29),
.B1(n_36),
.B2(n_70),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_15),
.A2(n_60),
.B1(n_63),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_15),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_78),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_15),
.A2(n_29),
.B1(n_36),
.B2(n_78),
.Y(n_161)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_17),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_17),
.A2(n_46),
.B1(n_60),
.B2(n_63),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_17),
.A2(n_29),
.B1(n_36),
.B2(n_46),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_125),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_124),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_102),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_22),
.B(n_102),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_80),
.C(n_86),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_23),
.B(n_80),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_55),
.B2(n_56),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_24),
.B(n_57),
.C(n_71),
.Y(n_123)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_41),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_28),
.A2(n_33),
.B(n_38),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_28),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_28),
.A2(n_33),
.B1(n_92),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_28),
.A2(n_33),
.B1(n_149),
.B2(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_28),
.A2(n_33),
.B1(n_161),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_28),
.A2(n_33),
.B1(n_193),
.B2(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_28),
.A2(n_33),
.B1(n_135),
.B2(n_226),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_28),
.A2(n_33),
.B1(n_219),
.B2(n_226),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_29),
.B(n_228),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_32),
.A2(n_35),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_32),
.A2(n_90),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_36),
.A2(n_50),
.B(n_135),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_43),
.A2(n_51),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_45),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_44),
.B(n_75),
.Y(n_191)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_45),
.A2(n_63),
.A3(n_74),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_84),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_47),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_47),
.A2(n_54),
.B1(n_84),
.B2(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_47),
.A2(n_54),
.B1(n_95),
.B2(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_47),
.A2(n_54),
.B1(n_143),
.B2(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_47),
.A2(n_54),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_47),
.A2(n_54),
.B1(n_205),
.B2(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_51),
.A2(n_96),
.B1(n_184),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_71),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_67),
.B2(n_69),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_59),
.B1(n_67),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_58),
.A2(n_59),
.B1(n_69),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_58),
.A2(n_59),
.B1(n_132),
.B2(n_136),
.Y(n_131)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_58),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_59),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_63),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g151 ( 
.A1(n_60),
.A2(n_62),
.A3(n_65),
.B1(n_134),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_61),
.B(n_63),
.Y(n_152)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_66),
.B(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_72),
.A2(n_76),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_72),
.A2(n_76),
.B1(n_156),
.B2(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_85),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_82),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_86),
.B(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_97),
.C(n_99),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_87),
.A2(n_88),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_89),
.B(n_93),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_97),
.B(n_99),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_123),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_113),
.B1(n_114),
.B2(n_122),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_110),
.B(n_112),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_110),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_107),
.A2(n_109),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_107),
.A2(n_109),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_266),
.B(n_270),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_176),
.B(n_254),
.C(n_265),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_162),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_128),
.B(n_162),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_146),
.C(n_153),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_129),
.A2(n_130),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_138),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_139),
.C(n_145),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_146),
.B(n_153),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_147),
.B(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.C(n_160),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_154),
.B(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_160),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_164),
.B(n_165),
.C(n_166),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_175),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_168),
.B(n_171),
.C(n_175),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_253),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_197),
.B(n_252),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_194),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_179),
.B(n_194),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_185),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_180),
.B(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_182),
.A2(n_185),
.B1(n_186),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_192),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_246),
.B(n_251),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_235),
.B(n_245),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_215),
.B(n_234),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_208),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_201),
.B(n_208),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_202),
.A2(n_203),
.B1(n_206),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_211),
.C(n_213),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_214),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_223),
.B(n_233),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_217),
.B(n_221),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_229),
.B(n_232),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_230),
.B(n_231),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_236),
.B(n_237),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_241),
.C(n_243),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_247),
.B(n_248),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_256),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_264),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_262),
.B2(n_263),
.Y(n_257)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_258),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_263),
.C(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_259),
.Y(n_263)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);


endmodule