module real_aes_10414_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_1929;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1893;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_1926;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1853;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_1159;
wire n_474;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_1102;
wire n_661;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1855;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_1192;
wire n_518;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1889;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1823;
wire n_1547;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1925;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1842;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1280;
wire n_394;
wire n_1352;
wire n_1323;
wire n_729;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1528 ( .A1(n_0), .A2(n_166), .B1(n_557), .B2(n_580), .Y(n_1528) );
AOI22xp33_ASAP7_75t_L g1535 ( .A1(n_0), .A2(n_166), .B1(n_517), .B2(n_1133), .Y(n_1535) );
INVxp67_ASAP7_75t_SL g786 ( .A(n_1), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_1), .A2(n_7), .B1(n_528), .B2(n_815), .Y(n_814) );
INVxp33_ASAP7_75t_L g988 ( .A(n_2), .Y(n_988) );
AOI21xp5_ASAP7_75t_L g1027 ( .A1(n_2), .A2(n_1028), .B(n_1030), .Y(n_1027) );
INVx1_ASAP7_75t_L g1066 ( .A(n_3), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_4), .A2(n_247), .B1(n_568), .B2(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_4), .A2(n_247), .B1(n_550), .B2(n_826), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g1898 ( .A1(n_5), .A2(n_16), .B1(n_719), .B2(n_1899), .Y(n_1898) );
INVxp67_ASAP7_75t_SL g1921 ( .A(n_5), .Y(n_1921) );
INVx1_ASAP7_75t_L g777 ( .A(n_6), .Y(n_777) );
INVx1_ASAP7_75t_L g785 ( .A(n_7), .Y(n_785) );
INVx1_ASAP7_75t_L g1787 ( .A(n_8), .Y(n_1787) );
INVxp67_ASAP7_75t_SL g1352 ( .A(n_9), .Y(n_1352) );
AOI22xp33_ASAP7_75t_L g1372 ( .A1(n_9), .A2(n_67), .B1(n_717), .B2(n_1056), .Y(n_1372) );
INVxp33_ASAP7_75t_SL g1893 ( .A(n_10), .Y(n_1893) );
AOI22xp33_ASAP7_75t_L g1905 ( .A1(n_10), .A2(n_332), .B1(n_1906), .B2(n_1907), .Y(n_1905) );
CKINVDCx5p33_ASAP7_75t_R g1465 ( .A(n_11), .Y(n_1465) );
INVx1_ASAP7_75t_L g1299 ( .A(n_12), .Y(n_1299) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_12), .A2(n_217), .B1(n_1048), .B2(n_1224), .Y(n_1315) );
INVx1_ASAP7_75t_L g1618 ( .A(n_13), .Y(n_1618) );
AOI22xp33_ASAP7_75t_SL g1533 ( .A1(n_14), .A2(n_314), .B1(n_730), .B2(n_831), .Y(n_1533) );
INVxp67_ASAP7_75t_L g1542 ( .A(n_14), .Y(n_1542) );
INVxp67_ASAP7_75t_SL g1889 ( .A(n_15), .Y(n_1889) );
OAI22xp5_ASAP7_75t_L g1917 ( .A1(n_15), .A2(n_233), .B1(n_492), .B2(n_795), .Y(n_1917) );
INVxp67_ASAP7_75t_SL g1922 ( .A(n_16), .Y(n_1922) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_17), .A2(n_262), .B1(n_521), .B2(n_571), .Y(n_666) );
AOI221xp5_ASAP7_75t_SL g684 ( .A1(n_17), .A2(n_685), .B1(n_686), .B2(n_694), .C(n_696), .Y(n_684) );
INVx1_ASAP7_75t_L g774 ( .A(n_18), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_18), .A2(n_65), .B1(n_792), .B2(n_810), .Y(n_817) );
INVxp33_ASAP7_75t_L g1387 ( .A(n_19), .Y(n_1387) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_19), .A2(n_33), .B1(n_579), .B2(n_1101), .Y(n_1409) );
INVx1_ASAP7_75t_L g894 ( .A(n_20), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_20), .A2(n_338), .B1(n_448), .B2(n_453), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g1607 ( .A1(n_21), .A2(n_128), .B1(n_1556), .B2(n_1564), .Y(n_1607) );
INVx1_ASAP7_75t_L g937 ( .A(n_22), .Y(n_937) );
INVxp67_ASAP7_75t_SL g1082 ( .A(n_23), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_23), .A2(n_228), .B1(n_719), .B2(n_1048), .Y(n_1105) );
OAI211xp5_ASAP7_75t_L g1423 ( .A1(n_24), .A2(n_443), .B(n_1054), .C(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1441 ( .A(n_24), .Y(n_1441) );
OAI222xp33_ASAP7_75t_L g1287 ( .A1(n_25), .A2(n_82), .B1(n_239), .B2(n_782), .C1(n_783), .C2(n_1288), .Y(n_1287) );
AOI22xp33_ASAP7_75t_SL g1321 ( .A1(n_25), .A2(n_191), .B1(n_1204), .B2(n_1205), .Y(n_1321) );
INVxp33_ASAP7_75t_L g1797 ( .A(n_26), .Y(n_1797) );
AOI221xp5_ASAP7_75t_L g1845 ( .A1(n_26), .A2(n_78), .B1(n_517), .B2(n_1189), .C(n_1846), .Y(n_1845) );
INVx1_ASAP7_75t_L g857 ( .A(n_27), .Y(n_857) );
AOI22xp33_ASAP7_75t_SL g871 ( .A1(n_27), .A2(n_207), .B1(n_831), .B2(n_832), .Y(n_871) );
CKINVDCx5p33_ASAP7_75t_R g1503 ( .A(n_28), .Y(n_1503) );
INVx1_ASAP7_75t_L g1520 ( .A(n_29), .Y(n_1520) );
OAI22xp5_ASAP7_75t_L g1539 ( .A1(n_29), .A2(n_32), .B1(n_794), .B2(n_1165), .Y(n_1539) );
AOI22xp33_ASAP7_75t_SL g1199 ( .A1(n_30), .A2(n_92), .B1(n_1200), .B2(n_1201), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_30), .A2(n_92), .B1(n_1048), .B2(n_1056), .Y(n_1219) );
CKINVDCx5p33_ASAP7_75t_R g1448 ( .A(n_31), .Y(n_1448) );
INVx1_ASAP7_75t_L g1521 ( .A(n_32), .Y(n_1521) );
INVx1_ASAP7_75t_L g1383 ( .A(n_33), .Y(n_1383) );
INVx1_ASAP7_75t_L g931 ( .A(n_34), .Y(n_931) );
INVx1_ASAP7_75t_L g1295 ( .A(n_35), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_35), .A2(n_185), .B1(n_1200), .B2(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g750 ( .A(n_36), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_36), .A2(n_232), .B1(n_448), .B2(n_630), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g1504 ( .A(n_37), .Y(n_1504) );
AOI22xp33_ASAP7_75t_L g1819 ( .A1(n_38), .A2(n_353), .B1(n_1820), .B2(n_1821), .Y(n_1819) );
INVxp67_ASAP7_75t_SL g1857 ( .A(n_38), .Y(n_1857) );
INVx1_ASAP7_75t_L g1473 ( .A(n_39), .Y(n_1473) );
OAI22xp5_ASAP7_75t_L g1505 ( .A1(n_39), .A2(n_188), .B1(n_463), .B2(n_471), .Y(n_1505) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_40), .A2(n_139), .B1(n_717), .B2(n_719), .Y(n_716) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_40), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_41), .A2(n_87), .B1(n_528), .B2(n_529), .Y(n_1399) );
AOI22xp33_ASAP7_75t_L g1407 ( .A1(n_41), .A2(n_87), .B1(n_548), .B2(n_1366), .Y(n_1407) );
OAI211xp5_ASAP7_75t_L g635 ( .A1(n_42), .A2(n_483), .B(n_636), .C(n_639), .Y(n_635) );
INVx1_ASAP7_75t_L g679 ( .A(n_42), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_43), .A2(n_122), .B1(n_509), .B2(n_514), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_43), .A2(n_122), .B1(n_719), .B2(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g381 ( .A(n_44), .Y(n_381) );
XNOR2xp5_ASAP7_75t_L g1459 ( .A(n_45), .B(n_1460), .Y(n_1459) );
AOI22xp5_ASAP7_75t_L g1628 ( .A1(n_45), .A2(n_120), .B1(n_1556), .B2(n_1564), .Y(n_1628) );
OAI211xp5_ASAP7_75t_L g705 ( .A1(n_46), .A2(n_483), .B(n_706), .C(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g728 ( .A(n_46), .Y(n_728) );
INVx1_ASAP7_75t_L g1590 ( .A(n_47), .Y(n_1590) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_48), .A2(n_63), .B1(n_390), .B2(n_500), .Y(n_602) );
OAI22xp33_ASAP7_75t_L g613 ( .A1(n_48), .A2(n_356), .B1(n_448), .B2(n_453), .Y(n_613) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_49), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_49), .A2(n_199), .B1(n_528), .B2(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g1523 ( .A(n_50), .Y(n_1523) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_51), .A2(n_240), .B1(n_1201), .B2(n_1208), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1365 ( .A1(n_51), .A2(n_240), .B1(n_1048), .B2(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1804 ( .A(n_52), .Y(n_1804) );
INVxp33_ASAP7_75t_L g1196 ( .A(n_53), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g1221 ( .A1(n_53), .A2(n_301), .B1(n_544), .B2(n_967), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_54), .A2(n_323), .B1(n_568), .B2(n_569), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_54), .A2(n_323), .B1(n_548), .B2(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_55), .A2(n_203), .B1(n_571), .B2(n_792), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_55), .A2(n_203), .B1(n_557), .B2(n_580), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g1608 ( .A1(n_56), .A2(n_76), .B1(n_1572), .B2(n_1586), .Y(n_1608) );
INVxp33_ASAP7_75t_SL g1067 ( .A(n_57), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_57), .A2(n_206), .B1(n_528), .B2(n_529), .Y(n_1087) );
INVxp33_ASAP7_75t_SL g1084 ( .A(n_58), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_58), .A2(n_73), .B1(n_1099), .B2(n_1101), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1825 ( .A1(n_59), .A2(n_202), .B1(n_1158), .B2(n_1826), .Y(n_1825) );
OAI22xp5_ASAP7_75t_L g1865 ( .A1(n_59), .A2(n_202), .B1(n_1866), .B2(n_1867), .Y(n_1865) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_60), .A2(n_86), .B1(n_463), .B2(n_471), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_60), .A2(n_86), .B1(n_548), .B2(n_549), .Y(n_559) );
INVxp67_ASAP7_75t_SL g1117 ( .A(n_61), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_61), .A2(n_225), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_62), .A2(n_368), .B1(n_463), .B2(n_471), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_62), .A2(n_368), .B1(n_681), .B2(n_682), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_63), .A2(n_184), .B1(n_589), .B2(n_591), .Y(n_588) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_64), .A2(n_142), .B1(n_390), .B2(n_500), .Y(n_642) );
INVx1_ASAP7_75t_L g675 ( .A(n_64), .Y(n_675) );
INVx1_ASAP7_75t_L g780 ( .A(n_65), .Y(n_780) );
INVx1_ASAP7_75t_L g790 ( .A(n_66), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_66), .A2(n_266), .B1(n_544), .B2(n_829), .Y(n_828) );
INVxp33_ASAP7_75t_SL g1353 ( .A(n_67), .Y(n_1353) );
AO22x2_ASAP7_75t_L g1332 ( .A1(n_68), .A2(n_1333), .B1(n_1373), .B2(n_1374), .Y(n_1332) );
CKINVDCx14_ASAP7_75t_R g1373 ( .A(n_68), .Y(n_1373) );
AOI22xp33_ASAP7_75t_L g1580 ( .A1(n_69), .A2(n_213), .B1(n_1556), .B2(n_1564), .Y(n_1580) );
CKINVDCx5p33_ASAP7_75t_R g1294 ( .A(n_70), .Y(n_1294) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_71), .A2(n_617), .B1(n_698), .B2(n_699), .Y(n_616) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_71), .Y(n_699) );
AO22x1_ASAP7_75t_SL g1598 ( .A1(n_71), .A2(n_129), .B1(n_1556), .B2(n_1564), .Y(n_1598) );
INVx1_ASAP7_75t_L g1340 ( .A(n_72), .Y(n_1340) );
INVxp67_ASAP7_75t_SL g1077 ( .A(n_73), .Y(n_1077) );
INVx1_ASAP7_75t_L g928 ( .A(n_74), .Y(n_928) );
INVx1_ASAP7_75t_L g1243 ( .A(n_75), .Y(n_1243) );
XOR2x2_ASAP7_75t_L g1782 ( .A(n_76), .B(n_1783), .Y(n_1782) );
AOI22xp33_ASAP7_75t_L g1875 ( .A1(n_76), .A2(n_1876), .B1(n_1923), .B2(n_1927), .Y(n_1875) );
INVx1_ASAP7_75t_L g600 ( .A(n_77), .Y(n_600) );
INVxp33_ASAP7_75t_L g1799 ( .A(n_78), .Y(n_1799) );
CKINVDCx5p33_ASAP7_75t_R g914 ( .A(n_79), .Y(n_914) );
AOI22xp5_ASAP7_75t_L g1581 ( .A1(n_80), .A2(n_227), .B1(n_1568), .B2(n_1572), .Y(n_1581) );
INVxp67_ASAP7_75t_SL g1344 ( .A(n_81), .Y(n_1344) );
AOI22xp33_ASAP7_75t_L g1361 ( .A1(n_81), .A2(n_310), .B1(n_1362), .B2(n_1363), .Y(n_1361) );
INVx1_ASAP7_75t_L g1304 ( .A(n_82), .Y(n_1304) );
INVxp67_ASAP7_75t_SL g1000 ( .A(n_83), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_83), .A2(n_287), .B1(n_1048), .B2(n_1056), .Y(n_1055) );
INVxp67_ASAP7_75t_SL g662 ( .A(n_84), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_84), .A2(n_102), .B1(n_689), .B2(n_692), .Y(n_688) );
INVx1_ASAP7_75t_L g714 ( .A(n_85), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g1444 ( .A1(n_88), .A2(n_271), .B1(n_1362), .B2(n_1445), .C(n_1446), .Y(n_1444) );
AOI22xp33_ASAP7_75t_L g1453 ( .A1(n_88), .A2(n_271), .B1(n_832), .B2(n_945), .Y(n_1453) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_89), .A2(n_98), .B1(n_533), .B2(n_1094), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_89), .A2(n_98), .B1(n_1099), .B2(n_1101), .Y(n_1098) );
AOI22xp5_ASAP7_75t_L g1567 ( .A1(n_90), .A2(n_113), .B1(n_1568), .B2(n_1572), .Y(n_1567) );
OAI22xp5_ASAP7_75t_L g1434 ( .A1(n_91), .A2(n_259), .B1(n_463), .B2(n_471), .Y(n_1434) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_91), .A2(n_259), .B1(n_550), .B2(n_945), .Y(n_1456) );
BUFx2_ASAP7_75t_L g460 ( .A(n_93), .Y(n_460) );
BUFx2_ASAP7_75t_L g503 ( .A(n_93), .Y(n_503) );
INVx1_ASAP7_75t_L g539 ( .A(n_93), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_94), .A2(n_188), .B1(n_823), .B2(n_1475), .Y(n_1474) );
OAI211xp5_ASAP7_75t_L g1500 ( .A1(n_94), .A2(n_483), .B(n_1501), .C(n_1502), .Y(n_1500) );
AOI22xp33_ASAP7_75t_L g1897 ( .A1(n_95), .A2(n_263), .B1(n_1070), .B2(n_1216), .Y(n_1897) );
INVxp67_ASAP7_75t_SL g1916 ( .A(n_95), .Y(n_1916) );
INVx1_ASAP7_75t_L g1069 ( .A(n_96), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_96), .A2(n_119), .B1(n_521), .B2(n_810), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1902 ( .A1(n_97), .A2(n_362), .B1(n_1048), .B2(n_1903), .Y(n_1902) );
AOI22xp33_ASAP7_75t_L g1910 ( .A1(n_97), .A2(n_362), .B1(n_1906), .B2(n_1911), .Y(n_1910) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_99), .A2(n_336), .B1(n_521), .B2(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_99), .A2(n_336), .B1(n_579), .B2(n_580), .Y(n_578) );
INVxp67_ASAP7_75t_SL g1337 ( .A(n_100), .Y(n_1337) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_100), .A2(n_318), .B1(n_641), .B2(n_795), .Y(n_1350) );
AO22x2_ASAP7_75t_L g1282 ( .A1(n_101), .A2(n_1283), .B1(n_1284), .B2(n_1329), .Y(n_1282) );
INVx1_ASAP7_75t_L g1329 ( .A(n_101), .Y(n_1329) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_102), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g1901 ( .A1(n_103), .A2(n_297), .B1(n_1070), .B2(n_1276), .Y(n_1901) );
AOI22xp33_ASAP7_75t_L g1913 ( .A1(n_103), .A2(n_297), .B1(n_1189), .B2(n_1265), .Y(n_1913) );
INVx1_ASAP7_75t_L g842 ( .A(n_104), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_104), .A2(n_365), .B1(n_808), .B2(n_864), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_105), .A2(n_293), .B1(n_528), .B2(n_1091), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_105), .A2(n_293), .B1(n_587), .B2(n_681), .Y(n_1102) );
XNOR2xp5_ASAP7_75t_L g404 ( .A(n_106), .B(n_405), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g1576 ( .A1(n_106), .A2(n_313), .B1(n_1556), .B2(n_1564), .Y(n_1576) );
CKINVDCx5p33_ASAP7_75t_R g1432 ( .A(n_107), .Y(n_1432) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_108), .A2(n_364), .B1(n_579), .B2(n_591), .Y(n_1532) );
INVxp33_ASAP7_75t_L g1544 ( .A(n_108), .Y(n_1544) );
AOI22xp33_ASAP7_75t_L g1629 ( .A1(n_109), .A2(n_274), .B1(n_1572), .B2(n_1586), .Y(n_1629) );
INVx1_ASAP7_75t_L g1496 ( .A(n_110), .Y(n_1496) );
OAI211xp5_ASAP7_75t_SL g1509 ( .A1(n_110), .A2(n_676), .B(n_787), .C(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g968 ( .A(n_111), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_112), .A2(n_114), .B1(n_463), .B2(n_471), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_112), .A2(n_114), .B1(n_548), .B2(n_730), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_115), .A2(n_123), .B1(n_783), .B2(n_847), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_115), .A2(n_123), .B1(n_492), .B2(n_795), .Y(n_852) );
INVxp67_ASAP7_75t_SL g1237 ( .A(n_116), .Y(n_1237) );
AOI22xp33_ASAP7_75t_SL g1261 ( .A1(n_116), .A2(n_251), .B1(n_1200), .B2(n_1262), .Y(n_1261) );
INVx1_ASAP7_75t_L g614 ( .A(n_117), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_118), .A2(n_276), .B1(n_967), .B2(n_1312), .Y(n_1316) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_118), .A2(n_276), .B1(n_1213), .B2(n_1327), .Y(n_1326) );
INVxp33_ASAP7_75t_SL g1063 ( .A(n_119), .Y(n_1063) );
INVx1_ASAP7_75t_L g961 ( .A(n_121), .Y(n_961) );
INVx1_ASAP7_75t_L g1601 ( .A(n_124), .Y(n_1601) );
CKINVDCx5p33_ASAP7_75t_R g1447 ( .A(n_125), .Y(n_1447) );
INVx1_ASAP7_75t_L g941 ( .A(n_126), .Y(n_941) );
OAI22xp33_ASAP7_75t_SL g974 ( .A1(n_126), .A2(n_230), .B1(n_390), .B2(n_463), .Y(n_974) );
AO22x2_ASAP7_75t_L g1512 ( .A1(n_127), .A2(n_1513), .B1(n_1545), .B2(n_1546), .Y(n_1512) );
INVx1_ASAP7_75t_L g1545 ( .A(n_127), .Y(n_1545) );
INVxp33_ASAP7_75t_SL g1193 ( .A(n_130), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_130), .A2(n_229), .B1(n_1223), .B2(n_1224), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_131), .A2(n_268), .B1(n_1070), .B2(n_1155), .Y(n_1154) );
INVxp67_ASAP7_75t_SL g1163 ( .A(n_131), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_132), .A2(n_214), .B1(n_1149), .B2(n_1224), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g1322 ( .A1(n_132), .A2(n_214), .B1(n_1208), .B2(n_1323), .Y(n_1322) );
XOR2xp5_ASAP7_75t_L g873 ( .A(n_133), .B(n_874), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_134), .A2(n_322), .B1(n_832), .B2(n_945), .Y(n_1527) );
AOI22xp33_ASAP7_75t_SL g1534 ( .A1(n_134), .A2(n_322), .B1(n_568), .B2(n_808), .Y(n_1534) );
INVx1_ASAP7_75t_L g1388 ( .A(n_135), .Y(n_1388) );
INVx1_ASAP7_75t_L g1121 ( .A(n_136), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_136), .A2(n_315), .B1(n_794), .B2(n_1165), .Y(n_1164) );
AOI22xp33_ASAP7_75t_SL g1203 ( .A1(n_137), .A2(n_307), .B1(n_1204), .B2(n_1205), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_137), .A2(n_307), .B1(n_967), .B2(n_1216), .Y(n_1215) );
INVxp33_ASAP7_75t_SL g1179 ( .A(n_138), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_138), .A2(n_354), .B1(n_1208), .B2(n_1210), .Y(n_1207) );
INVxp67_ASAP7_75t_SL g739 ( .A(n_139), .Y(n_739) );
INVxp67_ASAP7_75t_SL g1519 ( .A(n_140), .Y(n_1519) );
AOI22xp33_ASAP7_75t_L g1530 ( .A1(n_140), .A2(n_224), .B1(n_571), .B2(n_1133), .Y(n_1530) );
INVx1_ASAP7_75t_L g957 ( .A(n_141), .Y(n_957) );
OAI22xp33_ASAP7_75t_L g963 ( .A1(n_141), .A2(n_146), .B1(n_448), .B2(n_630), .Y(n_963) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_142), .A2(n_357), .B1(n_453), .B2(n_620), .Y(n_619) );
INVxp33_ASAP7_75t_L g1396 ( .A(n_143), .Y(n_1396) );
AOI22xp33_ASAP7_75t_L g1403 ( .A1(n_143), .A2(n_334), .B1(n_517), .B2(n_521), .Y(n_1403) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_144), .A2(n_220), .B1(n_1279), .B2(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1485 ( .A(n_144), .Y(n_1485) );
INVx1_ASAP7_75t_L g891 ( .A(n_145), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_145), .A2(n_302), .B1(n_620), .B2(n_630), .Y(n_916) );
INVx1_ASAP7_75t_L g960 ( .A(n_146), .Y(n_960) );
INVxp33_ASAP7_75t_SL g1517 ( .A(n_147), .Y(n_1517) );
AOI22xp33_ASAP7_75t_SL g1529 ( .A1(n_147), .A2(n_329), .B1(n_568), .B2(n_808), .Y(n_1529) );
INVx1_ASAP7_75t_L g1560 ( .A(n_148), .Y(n_1560) );
OAI211xp5_ASAP7_75t_L g477 ( .A1(n_149), .A2(n_478), .B(n_483), .C(n_490), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_149), .A2(n_270), .B1(n_545), .B2(n_557), .Y(n_556) );
INVxp33_ASAP7_75t_SL g1233 ( .A(n_150), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_150), .A2(n_304), .B1(n_1259), .B2(n_1265), .Y(n_1264) );
INVxp33_ASAP7_75t_SL g1113 ( .A(n_151), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_151), .A2(n_195), .B1(n_1129), .B2(n_1143), .Y(n_1142) );
CKINVDCx5p33_ASAP7_75t_R g840 ( .A(n_152), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_153), .A2(n_371), .B1(n_390), .B2(n_500), .Y(n_704) );
INVx1_ASAP7_75t_L g725 ( .A(n_153), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_154), .A2(n_244), .B1(n_507), .B2(n_512), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_154), .A2(n_244), .B1(n_548), .B2(n_549), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_155), .A2(n_258), .B1(n_810), .B2(n_811), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_155), .A2(n_258), .B1(n_822), .B2(n_823), .Y(n_821) );
XNOR2xp5_ASAP7_75t_L g984 ( .A(n_156), .B(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g1185 ( .A(n_157), .Y(n_1185) );
OAI22xp5_ASAP7_75t_L g1191 ( .A1(n_157), .A2(n_299), .B1(n_641), .B2(n_1165), .Y(n_1191) );
INVx1_ASAP7_75t_L g895 ( .A(n_158), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g1584 ( .A1(n_159), .A2(n_254), .B1(n_1585), .B2(n_1587), .C(n_1589), .Y(n_1584) );
AO22x2_ASAP7_75t_SL g1108 ( .A1(n_160), .A2(n_1109), .B1(n_1110), .B2(n_1171), .Y(n_1108) );
CKINVDCx16_ASAP7_75t_R g1109 ( .A(n_160), .Y(n_1109) );
INVx1_ASAP7_75t_L g1811 ( .A(n_161), .Y(n_1811) );
INVx1_ASAP7_75t_L g904 ( .A(n_162), .Y(n_904) );
OAI22xp33_ASAP7_75t_SL g921 ( .A1(n_162), .A2(n_173), .B1(n_390), .B2(n_463), .Y(n_921) );
INVxp33_ASAP7_75t_SL g1884 ( .A(n_163), .Y(n_1884) );
AOI22xp33_ASAP7_75t_L g1908 ( .A1(n_163), .A2(n_170), .B1(n_1130), .B2(n_1189), .Y(n_1908) );
INVx1_ASAP7_75t_L g1561 ( .A(n_164), .Y(n_1561) );
NAND2xp5_ASAP7_75t_L g1566 ( .A(n_164), .B(n_1559), .Y(n_1566) );
INVxp33_ASAP7_75t_SL g1347 ( .A(n_165), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g1369 ( .A1(n_165), .A2(n_341), .B1(n_1216), .B2(n_1370), .Y(n_1369) );
AOI22xp33_ASAP7_75t_SL g1816 ( .A1(n_167), .A2(n_192), .B1(n_1817), .B2(n_1818), .Y(n_1816) );
INVxp67_ASAP7_75t_SL g1856 ( .A(n_167), .Y(n_1856) );
OAI22xp5_ASAP7_75t_L g1421 ( .A1(n_168), .A2(n_179), .B1(n_448), .B2(n_630), .Y(n_1421) );
AOI221xp5_ASAP7_75t_L g1436 ( .A1(n_168), .A2(n_319), .B1(n_1135), .B2(n_1137), .C(n_1437), .Y(n_1436) );
INVx2_ASAP7_75t_L g393 ( .A(n_169), .Y(n_393) );
INVxp67_ASAP7_75t_SL g1887 ( .A(n_170), .Y(n_1887) );
AO221x2_ASAP7_75t_L g1614 ( .A1(n_171), .A2(n_218), .B1(n_1586), .B2(n_1615), .C(n_1616), .Y(n_1614) );
INVxp33_ASAP7_75t_L g1178 ( .A(n_172), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_172), .A2(n_344), .B1(n_1133), .B2(n_1213), .Y(n_1212) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_173), .A2(n_298), .B1(n_548), .B2(n_550), .Y(n_908) );
INVx1_ASAP7_75t_L g745 ( .A(n_174), .Y(n_745) );
OAI22xp33_ASAP7_75t_L g760 ( .A1(n_174), .A2(n_371), .B1(n_453), .B2(n_620), .Y(n_760) );
BUFx3_ASAP7_75t_L g414 ( .A(n_175), .Y(n_414) );
INVx1_ASAP7_75t_L g441 ( .A(n_175), .Y(n_441) );
INVx1_ASAP7_75t_L g1250 ( .A(n_176), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_176), .A2(n_265), .B1(n_995), .B2(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g994 ( .A(n_177), .Y(n_994) );
INVx1_ASAP7_75t_L g1242 ( .A(n_178), .Y(n_1242) );
INVx1_ASAP7_75t_L g1438 ( .A(n_179), .Y(n_1438) );
AOI22xp33_ASAP7_75t_SL g860 ( .A1(n_180), .A2(n_253), .B1(n_568), .B2(n_808), .Y(n_860) );
AOI22xp33_ASAP7_75t_SL g868 ( .A1(n_180), .A2(n_253), .B1(n_550), .B2(n_831), .Y(n_868) );
INVx1_ASAP7_75t_L g1793 ( .A(n_181), .Y(n_1793) );
AOI22xp33_ASAP7_75t_SL g1258 ( .A1(n_182), .A2(n_369), .B1(n_1130), .B2(n_1259), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1268 ( .A1(n_182), .A2(n_369), .B1(n_1101), .B2(n_1153), .Y(n_1268) );
INVx1_ASAP7_75t_L g838 ( .A(n_183), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_183), .A2(n_320), .B1(n_571), .B2(n_792), .Y(n_865) );
OAI211xp5_ASAP7_75t_SL g595 ( .A1(n_184), .A2(n_483), .B(n_596), .C(n_599), .Y(n_595) );
INVx1_ASAP7_75t_L g1292 ( .A(n_185), .Y(n_1292) );
INVxp33_ASAP7_75t_L g989 ( .A(n_186), .Y(n_989) );
AOI221xp5_ASAP7_75t_L g1025 ( .A1(n_186), .A2(n_309), .B1(n_507), .B2(n_529), .C(n_1026), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_187), .A2(n_249), .B1(n_1135), .B2(n_1137), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_187), .A2(n_249), .B1(n_1149), .B2(n_1150), .Y(n_1148) );
INVx1_ASAP7_75t_L g1236 ( .A(n_189), .Y(n_1236) );
INVx1_ASAP7_75t_L g752 ( .A(n_190), .Y(n_752) );
OAI211xp5_ASAP7_75t_L g756 ( .A1(n_190), .A2(n_443), .B(n_757), .C(n_759), .Y(n_756) );
INVx1_ASAP7_75t_L g1291 ( .A(n_191), .Y(n_1291) );
INVxp67_ASAP7_75t_SL g1861 ( .A(n_192), .Y(n_1861) );
AOI22xp33_ASAP7_75t_SL g1128 ( .A1(n_193), .A2(n_366), .B1(n_1129), .B2(n_1131), .Y(n_1128) );
AOI22xp33_ASAP7_75t_SL g1152 ( .A1(n_193), .A2(n_366), .B1(n_1101), .B2(n_1153), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_194), .A2(n_356), .B1(n_517), .B2(n_521), .Y(n_575) );
INVx1_ASAP7_75t_L g606 ( .A(n_194), .Y(n_606) );
INVx1_ASAP7_75t_L g1119 ( .A(n_195), .Y(n_1119) );
CKINVDCx5p33_ASAP7_75t_R g1833 ( .A(n_196), .Y(n_1833) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_197), .A2(n_702), .B1(n_761), .B2(n_762), .Y(n_701) );
INVx1_ASAP7_75t_L g762 ( .A(n_197), .Y(n_762) );
INVx1_ASAP7_75t_L g425 ( .A(n_198), .Y(n_425) );
INVx1_ASAP7_75t_L g442 ( .A(n_199), .Y(n_442) );
INVx1_ASAP7_75t_L g1384 ( .A(n_200), .Y(n_1384) );
XNOR2xp5_ASAP7_75t_L g1418 ( .A(n_201), .B(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g942 ( .A(n_204), .Y(n_942) );
OAI211xp5_ASAP7_75t_SL g972 ( .A1(n_204), .A2(n_478), .B(n_483), .C(n_973), .Y(n_972) );
AO22x2_ASAP7_75t_L g1376 ( .A1(n_205), .A2(n_1377), .B1(n_1411), .B2(n_1412), .Y(n_1376) );
INVx1_ASAP7_75t_L g1411 ( .A(n_205), .Y(n_1411) );
INVxp33_ASAP7_75t_SL g1064 ( .A(n_206), .Y(n_1064) );
INVx1_ASAP7_75t_L g855 ( .A(n_207), .Y(n_855) );
INVx1_ASAP7_75t_L g458 ( .A(n_208), .Y(n_458) );
INVx1_ASAP7_75t_L g1792 ( .A(n_208), .Y(n_1792) );
INVx1_ASAP7_75t_L g601 ( .A(n_209), .Y(n_601) );
INVx1_ASAP7_75t_L g715 ( .A(n_210), .Y(n_715) );
INVxp33_ASAP7_75t_SL g1247 ( .A(n_211), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_211), .A2(n_248), .B1(n_1149), .B2(n_1279), .Y(n_1278) );
INVxp67_ASAP7_75t_L g803 ( .A(n_212), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_212), .A2(n_303), .B1(n_831), .B2(n_832), .Y(n_830) );
INVxp67_ASAP7_75t_SL g885 ( .A(n_215), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_215), .A2(n_343), .B1(n_550), .B2(n_586), .Y(n_900) );
INVx1_ASAP7_75t_L g1492 ( .A(n_216), .Y(n_1492) );
OAI22xp5_ASAP7_75t_L g1507 ( .A1(n_216), .A2(n_223), .B1(n_448), .B2(n_630), .Y(n_1507) );
INVx1_ASAP7_75t_L g1298 ( .A(n_217), .Y(n_1298) );
AOI22xp33_ASAP7_75t_SL g1823 ( .A1(n_219), .A2(n_300), .B1(n_1818), .B2(n_1824), .Y(n_1823) );
OAI211xp5_ASAP7_75t_SL g1840 ( .A1(n_219), .A2(n_1841), .B(n_1842), .C(n_1847), .Y(n_1840) );
INVx1_ASAP7_75t_L g1481 ( .A(n_220), .Y(n_1481) );
AOI22xp5_ASAP7_75t_L g1555 ( .A1(n_221), .A2(n_286), .B1(n_1556), .B2(n_1564), .Y(n_1555) );
AOI22xp5_ASAP7_75t_L g1577 ( .A1(n_222), .A2(n_312), .B1(n_1568), .B2(n_1572), .Y(n_1577) );
INVx1_ASAP7_75t_L g1489 ( .A(n_223), .Y(n_1489) );
INVxp33_ASAP7_75t_SL g1516 ( .A(n_224), .Y(n_1516) );
INVxp33_ASAP7_75t_SL g1114 ( .A(n_225), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_226), .A2(n_311), .B1(n_586), .B2(n_587), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_226), .A2(n_311), .B1(n_463), .B2(n_471), .Y(n_594) );
INVxp33_ASAP7_75t_L g1080 ( .A(n_228), .Y(n_1080) );
INVxp67_ASAP7_75t_SL g1194 ( .A(n_229), .Y(n_1194) );
INVx1_ASAP7_75t_L g946 ( .A(n_230), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g1422 ( .A1(n_231), .A2(n_319), .B1(n_453), .B2(n_620), .Y(n_1422) );
INVx1_ASAP7_75t_L g1433 ( .A(n_231), .Y(n_1433) );
INVx1_ASAP7_75t_L g743 ( .A(n_232), .Y(n_743) );
INVxp67_ASAP7_75t_SL g1890 ( .A(n_233), .Y(n_1890) );
INVxp33_ASAP7_75t_L g1380 ( .A(n_234), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g1410 ( .A1(n_234), .A2(n_325), .B1(n_548), .B2(n_587), .Y(n_1410) );
INVxp33_ASAP7_75t_L g1395 ( .A(n_235), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_235), .A2(n_292), .B1(n_507), .B2(n_1007), .Y(n_1402) );
INVx1_ASAP7_75t_L g1116 ( .A(n_236), .Y(n_1116) );
INVx1_ASAP7_75t_L g881 ( .A(n_237), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g1400 ( .A1(n_238), .A2(n_359), .B1(n_521), .B2(n_810), .Y(n_1400) );
AOI22xp33_ASAP7_75t_L g1405 ( .A1(n_238), .A2(n_359), .B1(n_580), .B2(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1303 ( .A(n_239), .Y(n_1303) );
INVx1_ASAP7_75t_L g1892 ( .A(n_241), .Y(n_1892) );
INVxp33_ASAP7_75t_SL g1343 ( .A(n_242), .Y(n_1343) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_242), .A2(n_260), .B1(n_1189), .B2(n_1213), .Y(n_1360) );
INVx1_ASAP7_75t_L g416 ( .A(n_243), .Y(n_416) );
INVx1_ASAP7_75t_L g1602 ( .A(n_245), .Y(n_1602) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_246), .A2(n_316), .B1(n_448), .B2(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g653 ( .A(n_246), .Y(n_653) );
INVxp33_ASAP7_75t_SL g1248 ( .A(n_248), .Y(n_1248) );
CKINVDCx20_ASAP7_75t_R g1617 ( .A(n_250), .Y(n_1617) );
INVxp33_ASAP7_75t_SL g1234 ( .A(n_251), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_252), .A2(n_278), .B1(n_517), .B2(n_521), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_252), .A2(n_278), .B1(n_544), .B2(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g628 ( .A(n_255), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g1464 ( .A(n_256), .Y(n_1464) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_257), .A2(n_288), .B1(n_568), .B2(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g612 ( .A(n_257), .Y(n_612) );
INVx1_ASAP7_75t_L g1336 ( .A(n_260), .Y(n_1336) );
CKINVDCx5p33_ASAP7_75t_R g1023 ( .A(n_261), .Y(n_1023) );
INVxp67_ASAP7_75t_SL g687 ( .A(n_262), .Y(n_687) );
INVxp67_ASAP7_75t_SL g1919 ( .A(n_263), .Y(n_1919) );
INVx1_ASAP7_75t_L g948 ( .A(n_264), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_264), .A2(n_273), .B1(n_471), .B2(n_500), .Y(n_971) );
INVxp33_ASAP7_75t_SL g1252 ( .A(n_265), .Y(n_1252) );
INVxp33_ASAP7_75t_L g798 ( .A(n_266), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g1430 ( .A(n_267), .Y(n_1430) );
INVxp33_ASAP7_75t_L g1170 ( .A(n_268), .Y(n_1170) );
BUFx3_ASAP7_75t_L g415 ( .A(n_269), .Y(n_415) );
INVx1_ASAP7_75t_L g434 ( .A(n_269), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_270), .A2(n_340), .B1(n_390), .B2(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g1471 ( .A(n_272), .Y(n_1471) );
OAI22xp5_ASAP7_75t_L g1499 ( .A1(n_272), .A2(n_331), .B1(n_390), .B2(n_500), .Y(n_1499) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_273), .A2(n_282), .B1(n_453), .B2(n_620), .Y(n_964) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_275), .Y(n_389) );
INVx1_ASAP7_75t_L g541 ( .A(n_275), .Y(n_541) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_275), .B(n_467), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_275), .B(n_349), .Y(n_1017) );
INVx1_ASAP7_75t_L g997 ( .A(n_277), .Y(n_997) );
OAI221xp5_ASAP7_75t_L g1010 ( .A1(n_277), .A2(n_373), .B1(n_1011), .B2(n_1018), .C(n_1020), .Y(n_1010) );
AO22x2_ASAP7_75t_L g1229 ( .A1(n_279), .A2(n_1230), .B1(n_1280), .B2(n_1281), .Y(n_1229) );
INVx1_ASAP7_75t_L g1280 ( .A(n_279), .Y(n_1280) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_280), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_281), .A2(n_321), .B1(n_851), .B2(n_1213), .Y(n_1358) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_281), .A2(n_321), .B1(n_967), .B2(n_1312), .Y(n_1368) );
INVx1_ASAP7_75t_L g958 ( .A(n_282), .Y(n_958) );
INVx1_ASAP7_75t_L g627 ( .A(n_283), .Y(n_627) );
XNOR2xp5_ASAP7_75t_L g922 ( .A(n_284), .B(n_923), .Y(n_922) );
INVx2_ASAP7_75t_L g420 ( .A(n_285), .Y(n_420) );
OR2x2_ASAP7_75t_L g1791 ( .A(n_285), .B(n_1792), .Y(n_1791) );
INVx1_ASAP7_75t_L g770 ( .A(n_286), .Y(n_770) );
INVxp67_ASAP7_75t_SL g1003 ( .A(n_287), .Y(n_1003) );
INVxp67_ASAP7_75t_SL g611 ( .A(n_288), .Y(n_611) );
INVx1_ASAP7_75t_L g1307 ( .A(n_289), .Y(n_1307) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_289), .A2(n_295), .B1(n_1312), .B2(n_1314), .Y(n_1311) );
INVx1_ASAP7_75t_L g1181 ( .A(n_290), .Y(n_1181) );
INVx1_ASAP7_75t_L g1073 ( .A(n_291), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_291), .A2(n_327), .B1(n_794), .B2(n_795), .Y(n_1078) );
INVxp33_ASAP7_75t_L g1393 ( .A(n_292), .Y(n_1393) );
INVx1_ASAP7_75t_L g969 ( .A(n_294), .Y(n_969) );
INVx1_ASAP7_75t_L g1301 ( .A(n_295), .Y(n_1301) );
OAI211xp5_ASAP7_75t_L g621 ( .A1(n_296), .A2(n_443), .B(n_622), .C(n_625), .Y(n_621) );
INVx1_ASAP7_75t_L g655 ( .A(n_296), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_298), .A2(n_338), .B1(n_471), .B2(n_500), .Y(n_918) );
INVx1_ASAP7_75t_L g1186 ( .A(n_299), .Y(n_1186) );
OAI221xp5_ASAP7_75t_L g1852 ( .A1(n_300), .A2(n_1853), .B1(n_1854), .B2(n_1860), .C(n_1864), .Y(n_1852) );
INVxp67_ASAP7_75t_SL g1190 ( .A(n_301), .Y(n_1190) );
INVx1_ASAP7_75t_L g888 ( .A(n_302), .Y(n_888) );
INVx1_ASAP7_75t_L g800 ( .A(n_303), .Y(n_800) );
INVx1_ASAP7_75t_L g1239 ( .A(n_304), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_305), .A2(n_348), .B1(n_1200), .B2(n_1256), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_305), .A2(n_348), .B1(n_1270), .B2(n_1272), .Y(n_1269) );
INVx1_ASAP7_75t_L g907 ( .A(n_306), .Y(n_907) );
OAI211xp5_ASAP7_75t_SL g919 ( .A1(n_306), .A2(n_478), .B(n_483), .C(n_920), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_308), .A2(n_346), .B1(n_782), .B2(n_783), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_308), .A2(n_346), .B1(n_794), .B2(n_795), .Y(n_793) );
INVxp67_ASAP7_75t_SL g992 ( .A(n_309), .Y(n_992) );
INVxp67_ASAP7_75t_SL g1341 ( .A(n_310), .Y(n_1341) );
INVxp33_ASAP7_75t_L g1541 ( .A(n_314), .Y(n_1541) );
INVx1_ASAP7_75t_L g1123 ( .A(n_315), .Y(n_1123) );
INVx1_ASAP7_75t_L g646 ( .A(n_316), .Y(n_646) );
INVx1_ASAP7_75t_L g854 ( .A(n_317), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_317), .A2(n_351), .B1(n_557), .B2(n_829), .Y(n_870) );
INVxp67_ASAP7_75t_SL g1338 ( .A(n_318), .Y(n_1338) );
INVx1_ASAP7_75t_L g845 ( .A(n_320), .Y(n_845) );
OAI22xp33_ASAP7_75t_L g447 ( .A1(n_324), .A2(n_340), .B1(n_448), .B2(n_453), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_324), .A2(n_355), .B1(n_532), .B2(n_533), .Y(n_531) );
INVxp33_ASAP7_75t_L g1381 ( .A(n_325), .Y(n_1381) );
INVx1_ASAP7_75t_L g934 ( .A(n_326), .Y(n_934) );
INVx1_ASAP7_75t_L g1072 ( .A(n_327), .Y(n_1072) );
INVx1_ASAP7_75t_L g1385 ( .A(n_328), .Y(n_1385) );
INVxp33_ASAP7_75t_SL g1524 ( .A(n_329), .Y(n_1524) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_330), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g1563 ( .A(n_330), .B(n_381), .Y(n_1563) );
AND3x2_ASAP7_75t_L g1569 ( .A(n_330), .B(n_381), .C(n_1560), .Y(n_1569) );
OAI22xp5_ASAP7_75t_L g1508 ( .A1(n_331), .A2(n_361), .B1(n_453), .B2(n_620), .Y(n_1508) );
INVxp33_ASAP7_75t_SL g1885 ( .A(n_332), .Y(n_1885) );
INVx2_ASAP7_75t_L g394 ( .A(n_333), .Y(n_394) );
INVx1_ASAP7_75t_L g1391 ( .A(n_334), .Y(n_1391) );
INVx1_ASAP7_75t_L g709 ( .A(n_335), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g1021 ( .A1(n_337), .A2(n_535), .B(n_1022), .Y(n_1021) );
INVxp67_ASAP7_75t_SL g1046 ( .A(n_337), .Y(n_1046) );
INVx1_ASAP7_75t_L g1036 ( .A(n_339), .Y(n_1036) );
INVxp67_ASAP7_75t_SL g1349 ( .A(n_341), .Y(n_1349) );
AOI22xp5_ASAP7_75t_L g1877 ( .A1(n_342), .A2(n_1878), .B1(n_1879), .B2(n_1880), .Y(n_1877) );
CKINVDCx5p33_ASAP7_75t_R g1878 ( .A(n_342), .Y(n_1878) );
INVxp67_ASAP7_75t_SL g883 ( .A(n_343), .Y(n_883) );
INVxp67_ASAP7_75t_SL g1184 ( .A(n_344), .Y(n_1184) );
CKINVDCx5p33_ASAP7_75t_R g1425 ( .A(n_345), .Y(n_1425) );
INVx1_ASAP7_75t_L g878 ( .A(n_347), .Y(n_878) );
INVx1_ASAP7_75t_L g396 ( .A(n_349), .Y(n_396) );
INVx2_ASAP7_75t_L g467 ( .A(n_349), .Y(n_467) );
XNOR2xp5_ASAP7_75t_L g834 ( .A(n_350), .B(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g850 ( .A(n_351), .Y(n_850) );
INVx1_ASAP7_75t_L g1034 ( .A(n_352), .Y(n_1034) );
INVxp67_ASAP7_75t_SL g1863 ( .A(n_353), .Y(n_1863) );
INVxp33_ASAP7_75t_L g1182 ( .A(n_354), .Y(n_1182) );
INVx1_ASAP7_75t_L g409 ( .A(n_355), .Y(n_409) );
INVx1_ASAP7_75t_L g650 ( .A(n_357), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g1426 ( .A(n_358), .Y(n_1426) );
INVx1_ASAP7_75t_L g708 ( .A(n_360), .Y(n_708) );
INVx1_ASAP7_75t_L g1495 ( .A(n_361), .Y(n_1495) );
XOR2x2_ASAP7_75t_L g1059 ( .A(n_363), .B(n_1060), .Y(n_1059) );
INVxp67_ASAP7_75t_SL g1538 ( .A(n_364), .Y(n_1538) );
INVx1_ASAP7_75t_L g843 ( .A(n_365), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_367), .A2(n_372), .B1(n_1158), .B2(n_1159), .Y(n_1157) );
INVxp33_ASAP7_75t_L g1167 ( .A(n_367), .Y(n_1167) );
INVx1_ASAP7_75t_L g991 ( .A(n_370), .Y(n_991) );
INVxp67_ASAP7_75t_SL g1168 ( .A(n_372), .Y(n_1168) );
INVx1_ASAP7_75t_L g996 ( .A(n_373), .Y(n_996) );
AO22x1_ASAP7_75t_L g1173 ( .A1(n_374), .A2(n_1174), .B1(n_1175), .B2(n_1225), .Y(n_1173) );
INVxp67_ASAP7_75t_L g1174 ( .A(n_374), .Y(n_1174) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_397), .B(n_1549), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_384), .Y(n_378) );
AND2x4_ASAP7_75t_L g1874 ( .A(n_379), .B(n_385), .Y(n_1874) );
NOR2xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_SL g1926 ( .A(n_380), .Y(n_1926) );
NAND2xp5_ASAP7_75t_L g1932 ( .A(n_380), .B(n_382), .Y(n_1932) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g1925 ( .A(n_382), .B(n_1926), .Y(n_1925) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x6_ASAP7_75t_L g502 ( .A(n_387), .B(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g804 ( .A(n_387), .B(n_503), .Y(n_804) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g525 ( .A(n_388), .B(n_396), .Y(n_525) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g668 ( .A(n_389), .B(n_466), .Y(n_668) );
INVx8_ASAP7_75t_L g797 ( .A(n_390), .Y(n_797) );
OR2x6_ASAP7_75t_L g390 ( .A(n_391), .B(n_395), .Y(n_390) );
OR2x6_ASAP7_75t_L g500 ( .A(n_391), .B(n_465), .Y(n_500) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_391), .Y(n_654) );
INVx1_ASAP7_75t_L g749 ( .A(n_391), .Y(n_749) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_391), .Y(n_893) );
INVx2_ASAP7_75t_SL g953 ( .A(n_391), .Y(n_953) );
OAI21xp33_ASAP7_75t_L g1022 ( .A1(n_391), .A2(n_525), .B(n_1023), .Y(n_1022) );
INVx2_ASAP7_75t_SL g1440 ( .A(n_391), .Y(n_1440) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx2_ASAP7_75t_L g470 ( .A(n_393), .Y(n_470) );
AND2x4_ASAP7_75t_L g475 ( .A(n_393), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g482 ( .A(n_393), .Y(n_482) );
INVx1_ASAP7_75t_L g489 ( .A(n_393), .Y(n_489) );
AND2x2_ASAP7_75t_L g520 ( .A(n_393), .B(n_394), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_394), .B(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g476 ( .A(n_394), .Y(n_476) );
INVx1_ASAP7_75t_L g481 ( .A(n_394), .Y(n_481) );
INVx1_ASAP7_75t_L g494 ( .A(n_394), .Y(n_494) );
INVx1_ASAP7_75t_L g511 ( .A(n_394), .Y(n_511) );
AND2x4_ASAP7_75t_L g493 ( .A(n_395), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g795 ( .A(n_396), .B(n_497), .Y(n_795) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_396), .B(n_497), .Y(n_1165) );
XNOR2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_977), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
XNOR2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_766), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_615), .B1(n_764), .B2(n_765), .Y(n_402) );
INVx2_ASAP7_75t_L g764 ( .A(n_403), .Y(n_764) );
XOR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_563), .Y(n_403) );
NAND3x1_ASAP7_75t_L g405 ( .A(n_406), .B(n_461), .C(n_504), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_447), .B(n_456), .Y(n_406) );
NAND3xp33_ASAP7_75t_SL g407 ( .A(n_408), .B(n_430), .C(n_443), .Y(n_407) );
AOI222xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_416), .B2(n_417), .C1(n_425), .C2(n_426), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g607 ( .A(n_411), .Y(n_607) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g546 ( .A(n_412), .Y(n_546) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_412), .Y(n_829) );
BUFx3_ASAP7_75t_L g995 ( .A(n_412), .Y(n_995) );
BUFx4f_ASAP7_75t_L g1101 ( .A(n_412), .Y(n_1101) );
INVx1_ASAP7_75t_L g1371 ( .A(n_412), .Y(n_1371) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_413), .Y(n_446) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx2_ASAP7_75t_L g428 ( .A(n_414), .Y(n_428) );
AND2x4_ASAP7_75t_L g433 ( .A(n_414), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g424 ( .A(n_415), .Y(n_424) );
AND2x4_ASAP7_75t_L g440 ( .A(n_415), .B(n_441), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_416), .A2(n_425), .B1(n_491), .B2(n_495), .Y(n_490) );
AOI222xp33_ASAP7_75t_L g993 ( .A1(n_417), .A2(n_426), .B1(n_994), .B2(n_995), .C1(n_996), .C2(n_997), .Y(n_993) );
AOI222xp33_ASAP7_75t_L g1068 ( .A1(n_417), .A2(n_426), .B1(n_1069), .B2(n_1070), .C1(n_1072), .C2(n_1073), .Y(n_1068) );
AOI222xp33_ASAP7_75t_L g1183 ( .A1(n_417), .A2(n_426), .B1(n_829), .B2(n_1184), .C1(n_1185), .C2(n_1186), .Y(n_1183) );
AOI222xp33_ASAP7_75t_L g1390 ( .A1(n_417), .A2(n_426), .B1(n_1070), .B2(n_1384), .C1(n_1385), .C2(n_1391), .Y(n_1390) );
AOI222xp33_ASAP7_75t_L g1518 ( .A1(n_417), .A2(n_426), .B1(n_1370), .B2(n_1519), .C1(n_1520), .C2(n_1521), .Y(n_1518) );
AOI222xp33_ASAP7_75t_L g1886 ( .A1(n_417), .A2(n_426), .B1(n_1887), .B2(n_1888), .C1(n_1889), .C2(n_1890), .Y(n_1886) );
AND2x2_ASAP7_75t_SL g417 ( .A(n_418), .B(n_421), .Y(n_417) );
AND2x4_ASAP7_75t_L g454 ( .A(n_418), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g626 ( .A(n_418), .B(n_421), .Y(n_626) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g429 ( .A(n_420), .Y(n_429) );
INVx1_ASAP7_75t_L g438 ( .A(n_420), .Y(n_438) );
AND2x2_ASAP7_75t_L g554 ( .A(n_420), .B(n_458), .Y(n_554) );
INVx2_ASAP7_75t_L g562 ( .A(n_420), .Y(n_562) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g609 ( .A(n_422), .Y(n_609) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g691 ( .A(n_423), .Y(n_691) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g455 ( .A(n_424), .B(n_428), .Y(n_455) );
AOI222xp33_ASAP7_75t_L g605 ( .A1(n_426), .A2(n_600), .B1(n_601), .B2(n_606), .C1(n_607), .C2(n_608), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_426), .A2(n_626), .B1(n_627), .B2(n_628), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_426), .A2(n_626), .B1(n_708), .B2(n_709), .Y(n_759) );
INVx3_ASAP7_75t_L g783 ( .A(n_426), .Y(n_783) );
AOI222xp33_ASAP7_75t_L g912 ( .A1(n_426), .A2(n_608), .B1(n_895), .B2(n_913), .C1(n_914), .C2(n_915), .Y(n_912) );
AOI222xp33_ASAP7_75t_L g966 ( .A1(n_426), .A2(n_608), .B1(n_961), .B2(n_967), .C1(n_968), .C2(n_969), .Y(n_966) );
AOI222xp33_ASAP7_75t_L g1118 ( .A1(n_426), .A2(n_1119), .B1(n_1120), .B2(n_1121), .C1(n_1122), .C2(n_1123), .Y(n_1118) );
AOI222xp33_ASAP7_75t_L g1238 ( .A1(n_426), .A2(n_1122), .B1(n_1239), .B2(n_1240), .C1(n_1242), .C2(n_1243), .Y(n_1238) );
AOI222xp33_ASAP7_75t_L g1335 ( .A1(n_426), .A2(n_626), .B1(n_823), .B2(n_1336), .C1(n_1337), .C2(n_1338), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1424 ( .A1(n_426), .A2(n_626), .B1(n_1425), .B2(n_1426), .Y(n_1424) );
AOI22xp33_ASAP7_75t_L g1510 ( .A1(n_426), .A2(n_626), .B1(n_1503), .B2(n_1504), .Y(n_1510) );
AND2x6_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
BUFx3_ASAP7_75t_L g693 ( .A(n_427), .Y(n_693) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g432 ( .A(n_429), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_435), .B1(n_436), .B2(n_442), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_431), .A2(n_436), .B1(n_611), .B2(n_612), .Y(n_610) );
CKINVDCx6p67_ASAP7_75t_R g630 ( .A(n_431), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_431), .A2(n_436), .B1(n_785), .B2(n_786), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_431), .A2(n_436), .B1(n_842), .B2(n_843), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_431), .A2(n_839), .B1(n_988), .B2(n_989), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_431), .A2(n_775), .B1(n_1063), .B2(n_1064), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_431), .A2(n_775), .B1(n_1113), .B2(n_1114), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_431), .A2(n_839), .B1(n_1178), .B2(n_1179), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_431), .A2(n_775), .B1(n_1233), .B2(n_1234), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g1290 ( .A1(n_431), .A2(n_839), .B1(n_1291), .B2(n_1292), .Y(n_1290) );
AOI22xp33_ASAP7_75t_L g1342 ( .A1(n_431), .A2(n_775), .B1(n_1343), .B2(n_1344), .Y(n_1342) );
AOI22xp5_ASAP7_75t_L g1394 ( .A1(n_431), .A2(n_839), .B1(n_1395), .B2(n_1396), .Y(n_1394) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_431), .A2(n_775), .B1(n_1516), .B2(n_1517), .Y(n_1515) );
AOI221xp5_ASAP7_75t_L g1883 ( .A1(n_431), .A2(n_444), .B1(n_775), .B2(n_1884), .C(n_1885), .Y(n_1883) );
AND2x6_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g445 ( .A(n_432), .Y(n_445) );
INVx1_ASAP7_75t_L g449 ( .A(n_432), .Y(n_449) );
AND2x2_ASAP7_75t_L g779 ( .A(n_432), .B(n_580), .Y(n_779) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_433), .Y(n_548) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_433), .Y(n_586) );
BUFx2_ASAP7_75t_L g681 ( .A(n_433), .Y(n_681) );
INVx2_ASAP7_75t_SL g718 ( .A(n_433), .Y(n_718) );
BUFx3_ASAP7_75t_L g831 ( .A(n_433), .Y(n_831) );
BUFx6f_ASAP7_75t_L g930 ( .A(n_433), .Y(n_930) );
BUFx6f_ASAP7_75t_L g945 ( .A(n_433), .Y(n_945) );
HB1xp67_ASAP7_75t_L g1149 ( .A(n_433), .Y(n_1149) );
HB1xp67_ASAP7_75t_L g1223 ( .A(n_433), .Y(n_1223) );
INVx1_ASAP7_75t_L g452 ( .A(n_434), .Y(n_452) );
INVx4_ASAP7_75t_L g620 ( .A(n_436), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_436), .A2(n_454), .B1(n_991), .B2(n_992), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_436), .A2(n_454), .B1(n_1066), .B2(n_1067), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_436), .A2(n_454), .B1(n_1116), .B2(n_1117), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_436), .A2(n_454), .B1(n_1181), .B2(n_1182), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_436), .A2(n_454), .B1(n_1236), .B2(n_1237), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1293 ( .A1(n_436), .A2(n_454), .B1(n_1294), .B2(n_1295), .Y(n_1293) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_436), .A2(n_454), .B1(n_1340), .B2(n_1341), .Y(n_1339) );
AOI221xp5_ASAP7_75t_L g1392 ( .A1(n_436), .A2(n_444), .B1(n_454), .B2(n_1388), .C(n_1393), .Y(n_1392) );
AOI22xp33_ASAP7_75t_L g1522 ( .A1(n_436), .A2(n_454), .B1(n_1523), .B2(n_1524), .Y(n_1522) );
AOI22xp33_ASAP7_75t_L g1891 ( .A1(n_436), .A2(n_454), .B1(n_1892), .B2(n_1893), .Y(n_1891) );
AND2x6_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
AND2x4_ASAP7_75t_L g775 ( .A(n_437), .B(n_776), .Y(n_775) );
AND2x4_ASAP7_75t_L g839 ( .A(n_437), .B(n_776), .Y(n_839) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g608 ( .A(n_438), .B(n_609), .Y(n_608) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_439), .Y(n_587) );
INVx1_ASAP7_75t_L g683 ( .A(n_439), .Y(n_683) );
BUFx6f_ASAP7_75t_L g832 ( .A(n_439), .Y(n_832) );
INVx2_ASAP7_75t_L g947 ( .A(n_439), .Y(n_947) );
INVx1_ASAP7_75t_L g1367 ( .A(n_439), .Y(n_1367) );
INVx1_ASAP7_75t_L g1822 ( .A(n_439), .Y(n_1822) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_440), .Y(n_550) );
INVx1_ASAP7_75t_L g583 ( .A(n_440), .Y(n_583) );
INVx2_ASAP7_75t_L g722 ( .A(n_440), .Y(n_722) );
INVx1_ASAP7_75t_L g1151 ( .A(n_440), .Y(n_1151) );
INVx1_ASAP7_75t_L g451 ( .A(n_441), .Y(n_451) );
NAND3xp33_ASAP7_75t_SL g604 ( .A(n_443), .B(n_605), .C(n_610), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g911 ( .A(n_443), .B(n_912), .Y(n_911) );
NAND2xp5_ASAP7_75t_SL g965 ( .A(n_443), .B(n_966), .Y(n_965) );
NAND4xp25_ASAP7_75t_L g1061 ( .A(n_443), .B(n_1062), .C(n_1065), .D(n_1068), .Y(n_1061) );
NAND4xp25_ASAP7_75t_SL g1334 ( .A(n_443), .B(n_1335), .C(n_1339), .D(n_1342), .Y(n_1334) );
NAND4xp25_ASAP7_75t_L g1514 ( .A(n_443), .B(n_1515), .C(n_1518), .D(n_1522), .Y(n_1514) );
CKINVDCx8_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
INVx5_ASAP7_75t_L g787 ( .A(n_444), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g1286 ( .A(n_444), .B(n_1287), .Y(n_1286) );
AND2x4_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_446), .Y(n_580) );
INVx2_ASAP7_75t_L g592 ( .A(n_446), .Y(n_592) );
INVx1_ASAP7_75t_L g824 ( .A(n_446), .Y(n_824) );
BUFx6f_ASAP7_75t_L g1071 ( .A(n_446), .Y(n_1071) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx2_ASAP7_75t_L g674 ( .A(n_450), .Y(n_674) );
INVx1_ASAP7_75t_L g695 ( .A(n_450), .Y(n_695) );
BUFx2_ASAP7_75t_L g724 ( .A(n_450), .Y(n_724) );
INVx1_ASAP7_75t_L g936 ( .A(n_450), .Y(n_936) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
AND2x2_ASAP7_75t_L g624 ( .A(n_451), .B(n_452), .Y(n_624) );
INVx4_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI22xp5_ASAP7_75t_SL g773 ( .A1(n_454), .A2(n_774), .B1(n_775), .B2(n_777), .Y(n_773) );
AOI22xp5_ASAP7_75t_SL g837 ( .A1(n_454), .A2(n_838), .B1(n_839), .B2(n_840), .Y(n_837) );
BUFx2_ASAP7_75t_L g544 ( .A(n_455), .Y(n_544) );
INVx2_ASAP7_75t_L g558 ( .A(n_455), .Y(n_558) );
INVx6_ASAP7_75t_L g590 ( .A(n_455), .Y(n_590) );
AND2x2_ASAP7_75t_L g1836 ( .A(n_455), .B(n_1809), .Y(n_1836) );
OAI21xp5_ASAP7_75t_SL g603 ( .A1(n_456), .A2(n_604), .B(n_613), .Y(n_603) );
OAI31xp33_ASAP7_75t_SL g754 ( .A1(n_456), .A2(n_755), .A3(n_756), .B(n_760), .Y(n_754) );
AOI211xp5_ASAP7_75t_L g771 ( .A1(n_456), .A2(n_772), .B(n_788), .C(n_805), .Y(n_771) );
AOI211xp5_ASAP7_75t_L g835 ( .A1(n_456), .A2(n_836), .B(n_848), .C(n_858), .Y(n_835) );
OAI31xp33_ASAP7_75t_SL g909 ( .A1(n_456), .A2(n_910), .A3(n_911), .B(n_916), .Y(n_909) );
OAI31xp33_ASAP7_75t_L g962 ( .A1(n_456), .A2(n_963), .A3(n_964), .B(n_965), .Y(n_962) );
OAI31xp33_ASAP7_75t_SL g1420 ( .A1(n_456), .A2(n_1421), .A3(n_1422), .B(n_1423), .Y(n_1420) );
AOI211x1_ASAP7_75t_L g1513 ( .A1(n_456), .A2(n_1514), .B(n_1525), .C(n_1536), .Y(n_1513) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_459), .Y(n_456) );
AND2x4_ASAP7_75t_L g632 ( .A(n_457), .B(n_459), .Y(n_632) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g561 ( .A(n_458), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g1869 ( .A(n_459), .Y(n_1869) );
BUFx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g524 ( .A(n_460), .Y(n_524) );
OR2x6_ASAP7_75t_L g667 ( .A(n_460), .B(n_668), .Y(n_667) );
OAI31xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_477), .A3(n_499), .B(n_501), .Y(n_461) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_468), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g472 ( .A(n_465), .B(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g799 ( .A(n_465), .B(n_509), .Y(n_799) );
AND2x4_ASAP7_75t_L g1081 ( .A(n_465), .B(n_473), .Y(n_1081) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g487 ( .A(n_467), .Y(n_487) );
INVx2_ASAP7_75t_L g661 ( .A(n_468), .Y(n_661) );
BUFx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g649 ( .A(n_469), .Y(n_649) );
INVx1_ASAP7_75t_L g738 ( .A(n_469), .Y(n_738) );
AND2x4_ASAP7_75t_L g509 ( .A(n_470), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g1019 ( .A(n_470), .Y(n_1019) );
INVx5_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g801 ( .A1(n_472), .A2(n_777), .B1(n_802), .B2(n_803), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_472), .A2(n_802), .B1(n_840), .B2(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_472), .A2(n_799), .B1(n_1167), .B2(n_1168), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g1297 ( .A1(n_472), .A2(n_799), .B1(n_1298), .B2(n_1299), .Y(n_1297) );
AOI22xp5_ASAP7_75t_L g1351 ( .A1(n_472), .A2(n_799), .B1(n_1352), .B2(n_1353), .Y(n_1351) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_474), .Y(n_816) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g515 ( .A(n_475), .Y(n_515) );
BUFx6f_ASAP7_75t_L g808 ( .A(n_475), .Y(n_808) );
INVx1_ASAP7_75t_L g1008 ( .A(n_475), .Y(n_1008) );
AND2x4_ASAP7_75t_L g488 ( .A(n_476), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g656 ( .A(n_479), .Y(n_656) );
INVx1_ASAP7_75t_L g733 ( .A(n_479), .Y(n_733) );
BUFx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g598 ( .A(n_480), .Y(n_598) );
INVx3_ASAP7_75t_L g638 ( .A(n_480), .Y(n_638) );
INVx2_ASAP7_75t_L g751 ( .A(n_480), .Y(n_751) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_481), .B(n_482), .Y(n_880) );
INVx1_ASAP7_75t_L g497 ( .A(n_482), .Y(n_497) );
NAND4xp25_ASAP7_75t_SL g1245 ( .A(n_483), .B(n_1246), .C(n_1249), .D(n_1251), .Y(n_1245) );
NAND4xp25_ASAP7_75t_SL g1296 ( .A(n_483), .B(n_1297), .C(n_1300), .D(n_1306), .Y(n_1296) );
NAND4xp25_ASAP7_75t_L g1378 ( .A(n_483), .B(n_1379), .C(n_1382), .D(n_1386), .Y(n_1378) );
NAND3xp33_ASAP7_75t_SL g1428 ( .A(n_483), .B(n_1429), .C(n_1431), .Y(n_1428) );
CKINVDCx11_ASAP7_75t_R g483 ( .A(n_484), .Y(n_483) );
AOI211xp5_ASAP7_75t_L g789 ( .A1(n_484), .A2(n_790), .B(n_791), .C(n_793), .Y(n_789) );
AOI211xp5_ASAP7_75t_L g849 ( .A1(n_484), .A2(n_850), .B(n_851), .C(n_852), .Y(n_849) );
AOI211xp5_ASAP7_75t_L g1075 ( .A1(n_484), .A2(n_1076), .B(n_1077), .C(n_1078), .Y(n_1075) );
AOI211xp5_ASAP7_75t_L g1162 ( .A1(n_484), .A2(n_521), .B(n_1163), .C(n_1164), .Y(n_1162) );
AOI211xp5_ASAP7_75t_L g1188 ( .A1(n_484), .A2(n_1189), .B(n_1190), .C(n_1191), .Y(n_1188) );
AOI211xp5_ASAP7_75t_L g1348 ( .A1(n_484), .A2(n_811), .B(n_1349), .C(n_1350), .Y(n_1348) );
AOI211xp5_ASAP7_75t_L g1537 ( .A1(n_484), .A2(n_1189), .B(n_1538), .C(n_1539), .Y(n_1537) );
AOI211xp5_ASAP7_75t_L g1915 ( .A1(n_484), .A2(n_521), .B(n_1916), .C(n_1917), .Y(n_1915) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_488), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVxp67_ASAP7_75t_L g498 ( .A(n_486), .Y(n_498) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g540 ( .A(n_487), .B(n_541), .Y(n_540) );
BUFx3_ASAP7_75t_L g522 ( .A(n_488), .Y(n_522) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_488), .Y(n_535) );
BUFx3_ASAP7_75t_L g792 ( .A(n_488), .Y(n_792) );
INVx1_ASAP7_75t_L g812 ( .A(n_488), .Y(n_812) );
BUFx6f_ASAP7_75t_L g1133 ( .A(n_488), .Y(n_1133) );
BUFx2_ASAP7_75t_L g1145 ( .A(n_488), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_491), .A2(n_495), .B1(n_708), .B2(n_709), .Y(n_707) );
AOI222xp33_ASAP7_75t_L g1382 ( .A1(n_491), .A2(n_1145), .B1(n_1305), .B2(n_1383), .C1(n_1384), .C2(n_1385), .Y(n_1382) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_493), .A2(n_495), .B1(n_600), .B2(n_601), .Y(n_599) );
INVx2_ASAP7_75t_L g641 ( .A(n_493), .Y(n_641) );
INVx2_ASAP7_75t_L g794 ( .A(n_493), .Y(n_794) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_493), .A2(n_495), .B1(n_914), .B2(n_915), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_493), .A2(n_495), .B1(n_968), .B2(n_969), .Y(n_973) );
AOI222xp33_ASAP7_75t_SL g1429 ( .A1(n_493), .A2(n_1259), .B1(n_1305), .B2(n_1425), .C1(n_1426), .C2(n_1430), .Y(n_1429) );
AOI22xp33_ASAP7_75t_L g1502 ( .A1(n_493), .A2(n_495), .B1(n_1503), .B2(n_1504), .Y(n_1502) );
INVx1_ASAP7_75t_L g1013 ( .A(n_494), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1850 ( .A(n_494), .Y(n_1850) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_495), .A2(n_627), .B1(n_628), .B2(n_640), .Y(n_639) );
AOI222xp33_ASAP7_75t_L g1249 ( .A1(n_495), .A2(n_640), .B1(n_1143), .B2(n_1242), .C1(n_1243), .C2(n_1250), .Y(n_1249) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
AND2x4_ASAP7_75t_L g1305 ( .A(n_496), .B(n_498), .Y(n_1305) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx5_ASAP7_75t_L g802 ( .A(n_500), .Y(n_802) );
INVx4_ASAP7_75t_L g1308 ( .A(n_500), .Y(n_1308) );
OAI31xp33_ASAP7_75t_SL g593 ( .A1(n_501), .A2(n_594), .A3(n_595), .B(n_602), .Y(n_593) );
OAI31xp33_ASAP7_75t_L g633 ( .A1(n_501), .A2(n_634), .A3(n_635), .B(n_642), .Y(n_633) );
OAI31xp33_ASAP7_75t_L g703 ( .A1(n_501), .A2(n_704), .A3(n_705), .B(n_710), .Y(n_703) );
OAI31xp33_ASAP7_75t_SL g917 ( .A1(n_501), .A2(n_918), .A3(n_919), .B(n_921), .Y(n_917) );
OAI31xp33_ASAP7_75t_SL g970 ( .A1(n_501), .A2(n_971), .A3(n_972), .B(n_974), .Y(n_970) );
AOI221xp5_ASAP7_75t_L g1060 ( .A1(n_501), .A2(n_632), .B1(n_1061), .B2(n_1074), .C(n_1085), .Y(n_1060) );
AOI221x1_ASAP7_75t_L g1230 ( .A1(n_501), .A2(n_631), .B1(n_1231), .B2(n_1245), .C(n_1253), .Y(n_1230) );
AOI221x1_ASAP7_75t_L g1284 ( .A1(n_501), .A2(n_631), .B1(n_1285), .B2(n_1296), .C(n_1309), .Y(n_1284) );
AOI221x1_ASAP7_75t_L g1377 ( .A1(n_501), .A2(n_632), .B1(n_1378), .B2(n_1389), .C(n_1397), .Y(n_1377) );
OAI21xp5_ASAP7_75t_L g1427 ( .A1(n_501), .A2(n_1428), .B(n_1434), .Y(n_1427) );
OAI31xp33_ASAP7_75t_SL g1498 ( .A1(n_501), .A2(n_1499), .A3(n_1500), .B(n_1505), .Y(n_1498) );
CKINVDCx16_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
AOI31xp33_ASAP7_75t_L g1161 ( .A1(n_502), .A2(n_1162), .A3(n_1166), .B(n_1169), .Y(n_1161) );
AOI31xp33_ASAP7_75t_L g1187 ( .A1(n_502), .A2(n_1188), .A3(n_1192), .B(n_1195), .Y(n_1187) );
AOI31xp33_ASAP7_75t_SL g1914 ( .A1(n_502), .A2(n_1915), .A3(n_1918), .B(n_1920), .Y(n_1914) );
AND2x4_ASAP7_75t_L g560 ( .A(n_503), .B(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_L g671 ( .A(n_503), .B(n_561), .Y(n_671) );
AND2x4_ASAP7_75t_L g1835 ( .A(n_503), .B(n_1836), .Y(n_1835) );
AND4x1_ASAP7_75t_L g504 ( .A(n_505), .B(n_526), .C(n_542), .D(n_555), .Y(n_504) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_516), .C(n_523), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g1362 ( .A(n_508), .Y(n_1362) );
INVx1_ASAP7_75t_L g1906 ( .A(n_508), .Y(n_1906) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_509), .Y(n_528) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_509), .Y(n_568) );
BUFx6f_ASAP7_75t_L g864 ( .A(n_509), .Y(n_864) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_509), .B(n_1002), .Y(n_1001) );
BUFx2_ASAP7_75t_L g1140 ( .A(n_509), .Y(n_1140) );
BUFx2_ASAP7_75t_L g1200 ( .A(n_509), .Y(n_1200) );
INVx1_ASAP7_75t_L g1209 ( .A(n_509), .Y(n_1209) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g1494 ( .A(n_512), .Y(n_1494) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g886 ( .A(n_514), .Y(n_886) );
INVx2_ASAP7_75t_L g1202 ( .A(n_514), .Y(n_1202) );
INVx2_ASAP7_75t_L g1211 ( .A(n_514), .Y(n_1211) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_515), .Y(n_530) );
INVx3_ASAP7_75t_L g890 ( .A(n_515), .Y(n_890) );
INVx2_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g571 ( .A(n_518), .Y(n_571) );
INVx2_ASAP7_75t_L g810 ( .A(n_518), .Y(n_810) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx2_ASAP7_75t_L g532 ( .A(n_519), .Y(n_532) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_519), .B(n_1002), .Y(n_1037) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx3_ASAP7_75t_L g1029 ( .A(n_520), .Y(n_1029) );
HB1xp67_ASAP7_75t_L g1076 ( .A(n_521), .Y(n_1076) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x4_ASAP7_75t_L g1035 ( .A(n_522), .B(n_1005), .Y(n_1035) );
INVx1_ASAP7_75t_L g1328 ( .A(n_522), .Y(n_1328) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_523), .B(n_567), .C(n_570), .Y(n_566) );
NAND3xp33_ASAP7_75t_L g806 ( .A(n_523), .B(n_807), .C(n_809), .Y(n_806) );
NAND3xp33_ASAP7_75t_L g859 ( .A(n_523), .B(n_860), .C(n_861), .Y(n_859) );
NAND3xp33_ASAP7_75t_L g1089 ( .A(n_523), .B(n_1090), .C(n_1093), .Y(n_1089) );
INVx2_ASAP7_75t_L g1127 ( .A(n_523), .Y(n_1127) );
NAND3xp33_ASAP7_75t_L g1198 ( .A(n_523), .B(n_1199), .C(n_1203), .Y(n_1198) );
AOI33xp33_ASAP7_75t_L g1318 ( .A1(n_523), .A2(n_536), .A3(n_1319), .B1(n_1321), .B2(n_1322), .B3(n_1326), .Y(n_1318) );
NAND3xp33_ASAP7_75t_L g1398 ( .A(n_523), .B(n_1399), .C(n_1400), .Y(n_1398) );
BUFx3_ASAP7_75t_L g1449 ( .A(n_523), .Y(n_1449) );
AOI33xp33_ASAP7_75t_L g1531 ( .A1(n_523), .A2(n_560), .A3(n_1532), .B1(n_1533), .B2(n_1534), .B3(n_1535), .Y(n_1531) );
AND2x4_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
OR2x2_ASAP7_75t_L g552 ( .A(n_524), .B(n_553), .Y(n_552) );
OR2x6_ASAP7_75t_L g696 ( .A(n_524), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g818 ( .A(n_524), .B(n_819), .Y(n_818) );
OR2x2_ASAP7_75t_L g926 ( .A(n_524), .B(n_697), .Y(n_926) );
BUFx2_ASAP7_75t_L g1043 ( .A(n_524), .Y(n_1043) );
AND2x4_ASAP7_75t_L g1357 ( .A(n_524), .B(n_525), .Y(n_1357) );
INVx2_ASAP7_75t_L g1838 ( .A(n_524), .Y(n_1838) );
INVx1_ASAP7_75t_L g1859 ( .A(n_525), .Y(n_1859) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_531), .C(n_536), .Y(n_526) );
INVx1_ASAP7_75t_L g746 ( .A(n_529), .Y(n_746) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g569 ( .A(n_530), .Y(n_569) );
INVx2_ASAP7_75t_L g574 ( .A(n_530), .Y(n_574) );
INVx2_ASAP7_75t_L g664 ( .A(n_530), .Y(n_664) );
INVx3_ASAP7_75t_L g741 ( .A(n_530), .Y(n_741) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g851 ( .A(n_534), .Y(n_851) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g1205 ( .A(n_535), .Y(n_1205) );
NAND3xp33_ASAP7_75t_L g1086 ( .A(n_536), .B(n_1087), .C(n_1088), .Y(n_1086) );
NAND3xp33_ASAP7_75t_L g1206 ( .A(n_536), .B(n_1207), .C(n_1212), .Y(n_1206) );
NAND3xp33_ASAP7_75t_L g1260 ( .A(n_536), .B(n_1261), .C(n_1264), .Y(n_1260) );
AOI33xp33_ASAP7_75t_L g1355 ( .A1(n_536), .A2(n_1356), .A3(n_1358), .B1(n_1359), .B2(n_1360), .B3(n_1361), .Y(n_1355) );
CKINVDCx8_ASAP7_75t_R g1497 ( .A(n_536), .Y(n_1497) );
NAND3xp33_ASAP7_75t_L g1904 ( .A(n_536), .B(n_1905), .C(n_1908), .Y(n_1904) );
INVx5_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx6_ASAP7_75t_L g576 ( .A(n_537), .Y(n_576) );
OR2x6_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
NAND2x1p5_ASAP7_75t_L g1808 ( .A(n_538), .B(n_1809), .Y(n_1808) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g1790 ( .A(n_539), .B(n_1791), .Y(n_1790) );
INVx2_ASAP7_75t_L g819 ( .A(n_540), .Y(n_819) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .C(n_551), .Y(n_542) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_544), .Y(n_685) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g913 ( .A(n_546), .Y(n_913) );
INVx1_ASAP7_75t_L g1314 ( .A(n_546), .Y(n_1314) );
INVx2_ASAP7_75t_L g1271 ( .A(n_548), .Y(n_1271) );
BUFx3_ASAP7_75t_L g1899 ( .A(n_548), .Y(n_1899) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g932 ( .A(n_550), .Y(n_932) );
INVx1_ASAP7_75t_L g1827 ( .A(n_550), .Y(n_1827) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_551), .B(n_578), .C(n_581), .Y(n_577) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_551), .B(n_821), .C(n_825), .Y(n_820) );
NAND3xp33_ASAP7_75t_L g866 ( .A(n_551), .B(n_867), .C(n_868), .Y(n_866) );
NAND3xp33_ASAP7_75t_L g1097 ( .A(n_551), .B(n_1098), .C(n_1102), .Y(n_1097) );
NAND3xp33_ASAP7_75t_L g1214 ( .A(n_551), .B(n_1215), .C(n_1219), .Y(n_1214) );
AOI33xp33_ASAP7_75t_L g1310 ( .A1(n_551), .A2(n_670), .A3(n_1311), .B1(n_1315), .B2(n_1316), .B3(n_1317), .Y(n_1310) );
NAND3xp33_ASAP7_75t_L g1404 ( .A(n_551), .B(n_1405), .C(n_1407), .Y(n_1404) );
AOI33xp33_ASAP7_75t_L g1526 ( .A1(n_551), .A2(n_818), .A3(n_1527), .B1(n_1528), .B2(n_1529), .B3(n_1530), .Y(n_1526) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OAI22xp5_ASAP7_75t_SL g897 ( .A1(n_552), .A2(n_898), .B1(n_901), .B2(n_902), .Y(n_897) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g697 ( .A(n_554), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .C(n_560), .Y(n_555) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_SL g579 ( .A(n_558), .Y(n_579) );
NAND3xp33_ASAP7_75t_L g584 ( .A(n_560), .B(n_585), .C(n_588), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g827 ( .A(n_560), .B(n_828), .C(n_830), .Y(n_827) );
NAND3xp33_ASAP7_75t_L g869 ( .A(n_560), .B(n_870), .C(n_871), .Y(n_869) );
INVx1_ASAP7_75t_L g949 ( .A(n_560), .Y(n_949) );
NAND3xp33_ASAP7_75t_L g1103 ( .A(n_560), .B(n_1104), .C(n_1105), .Y(n_1103) );
NAND3xp33_ASAP7_75t_L g1220 ( .A(n_560), .B(n_1221), .C(n_1222), .Y(n_1220) );
AOI33xp33_ASAP7_75t_L g1364 ( .A1(n_560), .A2(n_1050), .A3(n_1365), .B1(n_1368), .B2(n_1369), .B3(n_1372), .Y(n_1364) );
NAND3xp33_ASAP7_75t_L g1408 ( .A(n_560), .B(n_1409), .C(n_1410), .Y(n_1408) );
AND2x4_ASAP7_75t_L g1809 ( .A(n_562), .B(n_1810), .Y(n_1809) );
XOR2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_614), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_593), .C(n_603), .Y(n_564) );
AND4x1_ASAP7_75t_L g565 ( .A(n_566), .B(n_572), .C(n_577), .D(n_584), .Y(n_565) );
INVx1_ASAP7_75t_L g651 ( .A(n_569), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .C(n_576), .Y(n_572) );
INVx2_ASAP7_75t_L g657 ( .A(n_576), .Y(n_657) );
INVx1_ASAP7_75t_L g753 ( .A(n_576), .Y(n_753) );
AOI33xp33_ASAP7_75t_L g1125 ( .A1(n_576), .A2(n_1126), .A3(n_1128), .B1(n_1134), .B2(n_1139), .B3(n_1142), .Y(n_1125) );
AOI221xp5_ASAP7_75t_L g1435 ( .A1(n_576), .A2(n_1436), .B1(n_1444), .B2(n_1449), .C(n_1450), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1798 ( .A(n_579), .B(n_1789), .Y(n_1798) );
HB1xp67_ASAP7_75t_L g1120 ( .A(n_580), .Y(n_1120) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x6_ASAP7_75t_L g1795 ( .A(n_583), .B(n_1790), .Y(n_1795) );
BUFx3_ASAP7_75t_L g1158 ( .A(n_586), .Y(n_1158) );
INVx1_ASAP7_75t_L g1476 ( .A(n_586), .Y(n_1476) );
INVx1_ASAP7_75t_L g1472 ( .A(n_587), .Y(n_1472) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g776 ( .A(n_590), .Y(n_776) );
INVx1_ASAP7_75t_L g822 ( .A(n_590), .Y(n_822) );
BUFx6f_ASAP7_75t_L g1100 ( .A(n_590), .Y(n_1100) );
INVx2_ASAP7_75t_L g1156 ( .A(n_590), .Y(n_1156) );
INVx2_ASAP7_75t_SL g1218 ( .A(n_590), .Y(n_1218) );
HB1xp67_ASAP7_75t_L g1277 ( .A(n_590), .Y(n_1277) );
INVx2_ASAP7_75t_L g1313 ( .A(n_590), .Y(n_1313) );
INVx1_ASAP7_75t_L g1241 ( .A(n_591), .Y(n_1241) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx3_ASAP7_75t_L g967 ( .A(n_592), .Y(n_967) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x6_ASAP7_75t_L g1032 ( .A(n_598), .B(n_1015), .Y(n_1032) );
OR2x2_ASAP7_75t_L g1864 ( .A(n_598), .B(n_1015), .Y(n_1864) );
INVx2_ASAP7_75t_L g782 ( .A(n_608), .Y(n_782) );
INVx1_ASAP7_75t_L g847 ( .A(n_608), .Y(n_847) );
INVx1_ASAP7_75t_L g765 ( .A(n_615), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_700), .B1(n_701), .B2(n_763), .Y(n_615) );
INVx1_ASAP7_75t_L g763 ( .A(n_616), .Y(n_763) );
INVx1_ASAP7_75t_L g698 ( .A(n_617), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_633), .C(n_643), .Y(n_617) );
OAI31xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .A3(n_629), .B(n_631), .Y(n_618) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g1289 ( .A(n_623), .Y(n_1289) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g678 ( .A(n_624), .Y(n_678) );
INVx1_ASAP7_75t_L g727 ( .A(n_624), .Y(n_727) );
BUFx2_ASAP7_75t_L g906 ( .A(n_624), .Y(n_906) );
BUFx4f_ASAP7_75t_L g939 ( .A(n_624), .Y(n_939) );
BUFx4f_ASAP7_75t_L g1122 ( .A(n_626), .Y(n_1122) );
AOI221x1_ASAP7_75t_L g985 ( .A1(n_631), .A2(n_986), .B1(n_998), .B2(n_1041), .C(n_1044), .Y(n_985) );
AOI211x1_ASAP7_75t_SL g1110 ( .A1(n_631), .A2(n_1111), .B(n_1124), .C(n_1161), .Y(n_1110) );
AOI211xp5_ASAP7_75t_L g1175 ( .A1(n_631), .A2(n_1176), .B(n_1187), .C(n_1197), .Y(n_1175) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI211x1_ASAP7_75t_SL g1333 ( .A1(n_632), .A2(n_1334), .B(n_1345), .C(n_1354), .Y(n_1333) );
OAI31xp33_ASAP7_75t_SL g1506 ( .A1(n_632), .A2(n_1507), .A3(n_1508), .B(n_1509), .Y(n_1506) );
INVx1_ASAP7_75t_L g1894 ( .A(n_632), .Y(n_1894) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g1487 ( .A(n_637), .Y(n_1487) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx2_ASAP7_75t_L g706 ( .A(n_638), .Y(n_706) );
OAI22xp33_ASAP7_75t_L g959 ( .A1(n_638), .A2(n_952), .B1(n_960), .B2(n_961), .Y(n_959) );
OAI21xp5_ASAP7_75t_SL g1026 ( .A1(n_638), .A2(n_994), .B(n_1027), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1446 ( .A1(n_638), .A2(n_654), .B1(n_1447), .B2(n_1448), .Y(n_1446) );
AOI222xp33_ASAP7_75t_L g1300 ( .A1(n_640), .A2(n_1301), .B1(n_1302), .B2(n_1303), .C1(n_1304), .C2(n_1305), .Y(n_1300) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NOR3xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_658), .C(n_684), .Y(n_643) );
NOR3xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_652), .C(n_657), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B1(n_650), .B2(n_651), .Y(n_645) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g884 ( .A(n_649), .Y(n_884) );
INVx1_ASAP7_75t_L g956 ( .A(n_649), .Y(n_956) );
HB1xp67_ASAP7_75t_L g1491 ( .A(n_649), .Y(n_1491) );
OAI22xp33_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_652) );
OAI22xp33_ASAP7_75t_L g732 ( .A1(n_654), .A2(n_714), .B1(n_715), .B2(n_733), .Y(n_732) );
OAI22xp33_ASAP7_75t_L g877 ( .A1(n_654), .A2(n_878), .B1(n_879), .B2(n_881), .Y(n_877) );
OAI22xp33_ASAP7_75t_L g1493 ( .A1(n_656), .A2(n_1494), .B1(n_1495), .B2(n_1496), .Y(n_1493) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_667), .B1(n_669), .B2(n_672), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_662), .B1(n_663), .B2(n_665), .C(n_666), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI33xp33_ASAP7_75t_L g731 ( .A1(n_667), .A2(n_732), .A3(n_734), .B1(n_742), .B2(n_747), .B3(n_753), .Y(n_731) );
OAI33xp33_ASAP7_75t_L g876 ( .A1(n_667), .A2(n_877), .A3(n_882), .B1(n_887), .B2(n_892), .B3(n_896), .Y(n_876) );
OAI33xp33_ASAP7_75t_L g950 ( .A1(n_667), .A2(n_896), .A3(n_951), .B1(n_954), .B2(n_955), .B3(n_959), .Y(n_950) );
INVx1_ASAP7_75t_L g1479 ( .A(n_667), .Y(n_1479) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_669), .A2(n_696), .B1(n_713), .B2(n_723), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_669), .A2(n_1045), .B1(n_1049), .B2(n_1051), .Y(n_1044) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_670), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g1896 ( .A(n_670), .B(n_1897), .C(n_1898), .Y(n_1896) );
BUFx4f_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx4_ASAP7_75t_L g901 ( .A(n_671), .Y(n_901) );
BUFx4f_ASAP7_75t_L g1160 ( .A(n_671), .Y(n_1160) );
AOI33xp33_ASAP7_75t_L g1815 ( .A1(n_671), .A2(n_1273), .A3(n_1816), .B1(n_1819), .B2(n_1823), .B3(n_1825), .Y(n_1815) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .B1(n_676), .B2(n_679), .C(n_680), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_673), .A2(n_676), .B1(n_714), .B2(n_715), .C(n_716), .Y(n_713) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g899 ( .A(n_674), .Y(n_899) );
INVx2_ASAP7_75t_L g903 ( .A(n_674), .Y(n_903) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_674), .Y(n_1053) );
OAI21xp33_ASAP7_75t_SL g686 ( .A1(n_676), .A2(n_687), .B(n_688), .Y(n_686) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI221xp5_ASAP7_75t_SL g1045 ( .A1(n_678), .A2(n_694), .B1(n_1023), .B2(n_1046), .C(n_1047), .Y(n_1045) );
BUFx3_ASAP7_75t_L g1452 ( .A(n_678), .Y(n_1452) );
OR2x6_ASAP7_75t_L g1801 ( .A(n_678), .B(n_1790), .Y(n_1801) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g1056 ( .A(n_683), .Y(n_1056) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2x1p5_ASAP7_75t_L g1806 ( .A(n_690), .B(n_1807), .Y(n_1806) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g1814 ( .A(n_693), .Y(n_1814) );
BUFx2_ASAP7_75t_L g1470 ( .A(n_694), .Y(n_1470) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g1050 ( .A(n_696), .Y(n_1050) );
CKINVDCx5p33_ASAP7_75t_R g1147 ( .A(n_696), .Y(n_1147) );
CKINVDCx5p33_ASAP7_75t_R g1273 ( .A(n_696), .Y(n_1273) );
OAI22xp5_ASAP7_75t_L g1462 ( .A1(n_696), .A2(n_901), .B1(n_1463), .B2(n_1469), .Y(n_1462) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g761 ( .A(n_702), .Y(n_761) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_711), .C(n_754), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_731), .Y(n_711) );
AND2x2_ASAP7_75t_L g1788 ( .A(n_717), .B(n_1789), .Y(n_1788) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_SL g826 ( .A(n_718), .Y(n_826) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g1224 ( .A(n_720), .Y(n_1224) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
BUFx2_ASAP7_75t_L g730 ( .A(n_721), .Y(n_730) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g1159 ( .A(n_722), .Y(n_1159) );
OAI221xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B1(n_726), .B2(n_728), .C(n_729), .Y(n_723) );
OAI221xp5_ASAP7_75t_L g1463 ( .A1(n_724), .A2(n_757), .B1(n_1464), .B2(n_1465), .C(n_1466), .Y(n_1463) );
BUFx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g758 ( .A(n_727), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B1(n_739), .B2(n_740), .Y(n_734) );
INVx2_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g744 ( .A(n_737), .Y(n_744) );
INVx2_ASAP7_75t_L g1482 ( .A(n_737), .Y(n_1482) );
INVx2_ASAP7_75t_L g1843 ( .A(n_737), .Y(n_1843) );
BUFx3_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_743), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_742) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_750), .B1(n_751), .B2(n_752), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OAI22xp33_ASAP7_75t_L g892 ( .A1(n_751), .A2(n_893), .B1(n_894), .B2(n_895), .Y(n_892) );
OAI221xp5_ASAP7_75t_L g898 ( .A1(n_757), .A2(n_878), .B1(n_881), .B2(n_899), .C(n_900), .Y(n_898) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
XOR2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_872), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_769), .B1(n_833), .B2(n_834), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
XNOR2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
NAND4xp25_ASAP7_75t_L g772 ( .A(n_773), .B(n_778), .C(n_784), .D(n_787), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_780), .B(n_781), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g844 ( .A1(n_779), .A2(n_845), .B(n_846), .Y(n_844) );
NAND4xp25_ASAP7_75t_L g836 ( .A(n_787), .B(n_837), .C(n_841), .D(n_844), .Y(n_836) );
NAND4xp25_ASAP7_75t_L g986 ( .A(n_787), .B(n_987), .C(n_990), .D(n_993), .Y(n_986) );
NAND4xp25_ASAP7_75t_SL g1111 ( .A(n_787), .B(n_1112), .C(n_1115), .D(n_1118), .Y(n_1111) );
NAND4xp25_ASAP7_75t_SL g1176 ( .A(n_787), .B(n_1177), .C(n_1180), .D(n_1183), .Y(n_1176) );
BUFx2_ASAP7_75t_L g1244 ( .A(n_787), .Y(n_1244) );
AOI31xp33_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_796), .A3(n_801), .B(n_804), .Y(n_788) );
BUFx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_SL g796 ( .A1(n_797), .A2(n_798), .B1(n_799), .B2(n_800), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_797), .A2(n_799), .B1(n_854), .B2(n_855), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_797), .A2(n_802), .B1(n_1066), .B2(n_1084), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_797), .A2(n_802), .B1(n_1116), .B2(n_1170), .Y(n_1169) );
AOI22xp33_ASAP7_75t_SL g1195 ( .A1(n_797), .A2(n_802), .B1(n_1181), .B2(n_1196), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1251 ( .A1(n_797), .A2(n_802), .B1(n_1236), .B2(n_1252), .Y(n_1251) );
AOI22xp33_ASAP7_75t_L g1306 ( .A1(n_797), .A2(n_1294), .B1(n_1307), .B2(n_1308), .Y(n_1306) );
AOI22xp5_ASAP7_75t_L g1346 ( .A1(n_797), .A2(n_802), .B1(n_1340), .B2(n_1347), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_797), .A2(n_802), .B1(n_1387), .B2(n_1388), .Y(n_1386) );
AOI22xp33_ASAP7_75t_L g1431 ( .A1(n_797), .A2(n_1308), .B1(n_1432), .B2(n_1433), .Y(n_1431) );
AOI22xp33_ASAP7_75t_SL g1543 ( .A1(n_797), .A2(n_802), .B1(n_1523), .B2(n_1544), .Y(n_1543) );
AOI22xp5_ASAP7_75t_L g1918 ( .A1(n_797), .A2(n_1308), .B1(n_1892), .B2(n_1919), .Y(n_1918) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_799), .A2(n_1080), .B1(n_1081), .B2(n_1082), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_799), .A2(n_1081), .B1(n_1193), .B2(n_1194), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_799), .A2(n_1081), .B1(n_1247), .B2(n_1248), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_799), .A2(n_1081), .B1(n_1380), .B2(n_1381), .Y(n_1379) );
AOI22xp33_ASAP7_75t_SL g1540 ( .A1(n_799), .A2(n_1081), .B1(n_1541), .B2(n_1542), .Y(n_1540) );
AOI22xp5_ASAP7_75t_SL g1920 ( .A1(n_799), .A2(n_1081), .B1(n_1921), .B2(n_1922), .Y(n_1920) );
AOI31xp33_ASAP7_75t_L g848 ( .A1(n_804), .A2(n_849), .A3(n_853), .B(n_856), .Y(n_848) );
AOI31xp33_ASAP7_75t_L g1345 ( .A1(n_804), .A2(n_1346), .A3(n_1348), .B(n_1351), .Y(n_1345) );
AOI31xp33_ASAP7_75t_L g1536 ( .A1(n_804), .A2(n_1537), .A3(n_1540), .B(n_1543), .Y(n_1536) );
NAND4xp25_ASAP7_75t_L g805 ( .A(n_806), .B(n_813), .C(n_820), .D(n_827), .Y(n_805) );
INVx2_ASAP7_75t_SL g1138 ( .A(n_808), .Y(n_1138) );
BUFx3_ASAP7_75t_L g1141 ( .A(n_808), .Y(n_1141) );
INVx2_ASAP7_75t_SL g1257 ( .A(n_808), .Y(n_1257) );
INVx4_ASAP7_75t_L g1263 ( .A(n_808), .Y(n_1263) );
INVx2_ASAP7_75t_SL g1844 ( .A(n_808), .Y(n_1844) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NAND3xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_817), .C(n_818), .Y(n_813) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND3xp33_ASAP7_75t_L g862 ( .A(n_818), .B(n_863), .C(n_865), .Y(n_862) );
INVx1_ASAP7_75t_L g896 ( .A(n_818), .Y(n_896) );
NAND3xp33_ASAP7_75t_L g1401 ( .A(n_818), .B(n_1402), .C(n_1403), .Y(n_1401) );
INVx1_ASAP7_75t_L g1030 ( .A(n_819), .Y(n_1030) );
INVx2_ASAP7_75t_SL g1846 ( .A(n_819), .Y(n_1846) );
BUFx2_ASAP7_75t_L g1820 ( .A(n_822), .Y(n_1820) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
HB1xp67_ASAP7_75t_L g1818 ( .A(n_829), .Y(n_1818) );
NAND2xp5_ASAP7_75t_L g1830 ( .A(n_829), .B(n_1831), .Y(n_1830) );
BUFx2_ASAP7_75t_SL g1888 ( .A(n_829), .Y(n_1888) );
BUFx3_ASAP7_75t_L g1817 ( .A(n_831), .Y(n_1817) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NAND4xp25_ASAP7_75t_L g858 ( .A(n_859), .B(n_862), .C(n_866), .D(n_869), .Y(n_858) );
INVx2_ASAP7_75t_SL g1136 ( .A(n_864), .Y(n_1136) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_922), .B1(n_975), .B2(n_976), .Y(n_872) );
INVx1_ASAP7_75t_L g975 ( .A(n_873), .Y(n_975) );
NAND3xp33_ASAP7_75t_L g874 ( .A(n_875), .B(n_909), .C(n_917), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_897), .Y(n_875) );
OAI22xp33_ASAP7_75t_L g951 ( .A1(n_879), .A2(n_934), .B1(n_937), .B2(n_952), .Y(n_951) );
INVx2_ASAP7_75t_L g1443 ( .A(n_879), .Y(n_1443) );
BUFx3_ASAP7_75t_L g1501 ( .A(n_879), .Y(n_1501) );
BUFx6f_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
OAI22xp33_ASAP7_75t_SL g882 ( .A1(n_883), .A2(n_884), .B1(n_885), .B2(n_886), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_884), .A2(n_888), .B1(n_889), .B2(n_891), .Y(n_887) );
OAI22xp33_ASAP7_75t_L g954 ( .A1(n_884), .A2(n_889), .B1(n_928), .B2(n_931), .Y(n_954) );
INVx1_ASAP7_75t_L g1445 ( .A(n_886), .Y(n_1445) );
INVx1_ASAP7_75t_L g1484 ( .A(n_886), .Y(n_1484) );
OAI22xp33_ASAP7_75t_L g955 ( .A1(n_889), .A2(n_956), .B1(n_957), .B2(n_958), .Y(n_955) );
INVx2_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
BUFx3_ASAP7_75t_L g1907 ( .A(n_890), .Y(n_1907) );
OAI22xp5_ASAP7_75t_SL g1450 ( .A1(n_901), .A2(n_926), .B1(n_1451), .B2(n_1454), .Y(n_1450) );
OAI221xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_904), .B1(n_905), .B2(n_907), .C(n_908), .Y(n_902) );
OAI221xp5_ASAP7_75t_L g1451 ( .A1(n_903), .A2(n_1447), .B1(n_1448), .B2(n_1452), .C(n_1453), .Y(n_1451) );
OAI221xp5_ASAP7_75t_L g1454 ( .A1(n_903), .A2(n_1430), .B1(n_1432), .B2(n_1455), .C(n_1456), .Y(n_1454) );
HB1xp67_ASAP7_75t_L g1054 ( .A(n_905), .Y(n_1054) );
INVx2_ASAP7_75t_SL g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g976 ( .A(n_922), .Y(n_976) );
NAND3xp33_ASAP7_75t_L g923 ( .A(n_924), .B(n_962), .C(n_970), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g924 ( .A(n_925), .B(n_950), .Y(n_924) );
OAI33xp33_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_927), .A3(n_933), .B1(n_940), .B2(n_943), .B3(n_949), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_928), .A2(n_929), .B1(n_931), .B2(n_932), .Y(n_927) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
BUFx4f_ASAP7_75t_L g1048 ( .A(n_930), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_935), .B1(n_937), .B2(n_938), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_935), .A2(n_938), .B1(n_941), .B2(n_942), .Y(n_940) );
INVx2_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx2_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g1455 ( .A(n_939), .Y(n_1455) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_944), .A2(n_946), .B1(n_947), .B2(n_948), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx2_ASAP7_75t_SL g1468 ( .A(n_945), .Y(n_1468) );
INVx1_ASAP7_75t_L g1272 ( .A(n_947), .Y(n_1272) );
INVx1_ASAP7_75t_L g1279 ( .A(n_947), .Y(n_1279) );
OAI22xp33_ASAP7_75t_L g1486 ( .A1(n_952), .A2(n_1464), .B1(n_1465), .B2(n_1487), .Y(n_1486) );
OAI22xp33_ASAP7_75t_L g1488 ( .A1(n_952), .A2(n_1489), .B1(n_1490), .B2(n_1492), .Y(n_1488) );
OAI221xp5_ASAP7_75t_L g1854 ( .A1(n_952), .A2(n_1855), .B1(n_1856), .B2(n_1857), .C(n_1858), .Y(n_1854) );
INVx2_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_978), .A2(n_979), .B1(n_1415), .B2(n_1548), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
XNOR2xp5_ASAP7_75t_L g979 ( .A(n_980), .B(n_1227), .Y(n_979) );
XNOR2xp5_ASAP7_75t_L g980 ( .A(n_981), .B(n_1107), .Y(n_980) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_982), .A2(n_983), .B1(n_1057), .B2(n_1106), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
AOI222xp33_ASAP7_75t_L g1033 ( .A1(n_991), .A2(n_1034), .B1(n_1035), .B2(n_1036), .C1(n_1037), .C2(n_1038), .Y(n_1033) );
NAND3xp33_ASAP7_75t_L g998 ( .A(n_999), .B(n_1009), .C(n_1033), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g999 ( .A1(n_1000), .A2(n_1001), .B1(n_1003), .B2(n_1004), .Y(n_999) );
INVx3_ASAP7_75t_L g1866 ( .A(n_1001), .Y(n_1866) );
INVx2_ASAP7_75t_L g1006 ( .A(n_1002), .Y(n_1006) );
INVx3_ASAP7_75t_L g1867 ( .A(n_1004), .Y(n_1867) );
AND2x4_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1007), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1007), .Y(n_1092) );
INVx2_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1008), .Y(n_1325) );
NOR3xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1025), .C(n_1031), .Y(n_1009) );
NAND2x1p5_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1014), .Y(n_1011) );
INVx2_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
OR2x6_ASAP7_75t_L g1018 ( .A(n_1015), .B(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1015), .Y(n_1040) );
INVx2_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
CKINVDCx11_ASAP7_75t_R g1851 ( .A(n_1018), .Y(n_1851) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1024), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_1028), .B(n_1040), .Y(n_1039) );
BUFx2_ASAP7_75t_L g1204 ( .A(n_1028), .Y(n_1204) );
INVx2_ASAP7_75t_SL g1028 ( .A(n_1029), .Y(n_1028) );
INVx2_ASAP7_75t_SL g1096 ( .A(n_1029), .Y(n_1096) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1029), .Y(n_1130) );
INVx2_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
OAI221xp5_ASAP7_75t_SL g1051 ( .A1(n_1034), .A2(n_1036), .B1(n_1052), .B2(n_1054), .C(n_1055), .Y(n_1051) );
INVx8_ASAP7_75t_L g1841 ( .A(n_1035), .Y(n_1841) );
CKINVDCx6p67_ASAP7_75t_R g1853 ( .A(n_1037), .Y(n_1853) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
NOR2xp67_ASAP7_75t_L g1837 ( .A(n_1039), .B(n_1838), .Y(n_1837) );
AND2x2_ASAP7_75t_L g1849 ( .A(n_1040), .B(n_1850), .Y(n_1849) );
INVx2_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
CKINVDCx8_ASAP7_75t_R g1042 ( .A(n_1043), .Y(n_1042) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1059), .Y(n_1106) );
BUFx6f_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
NAND3xp33_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1079), .C(n_1083), .Y(n_1074) );
NAND4xp25_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1089), .C(n_1097), .D(n_1103), .Y(n_1085) );
INVx1_ASAP7_75t_L g1862 ( .A(n_1091), .Y(n_1862) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1092), .Y(n_1320) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
BUFx2_ASAP7_75t_L g1213 ( .A(n_1096), .Y(n_1213) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1096), .Y(n_1266) );
HB1xp67_ASAP7_75t_L g1824 ( .A(n_1099), .Y(n_1824) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx4_ASAP7_75t_L g1153 ( .A(n_1100), .Y(n_1153) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1100), .Y(n_1406) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_1108), .A2(n_1172), .B1(n_1173), .B2(n_1226), .Y(n_1107) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1108), .Y(n_1226) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1110), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1146), .Y(n_1124) );
NAND3xp33_ASAP7_75t_L g1254 ( .A(n_1126), .B(n_1255), .C(n_1258), .Y(n_1254) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
BUFx3_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
INVx2_ASAP7_75t_SL g1131 ( .A(n_1132), .Y(n_1131) );
INVx2_ASAP7_75t_SL g1132 ( .A(n_1133), .Y(n_1132) );
BUFx6f_ASAP7_75t_L g1189 ( .A(n_1133), .Y(n_1189) );
INVx3_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1144), .Y(n_1259) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1144), .Y(n_1302) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
AOI33xp33_ASAP7_75t_L g1146 ( .A1(n_1147), .A2(n_1148), .A3(n_1152), .B1(n_1154), .B2(n_1157), .B3(n_1160), .Y(n_1146) );
NAND3xp33_ASAP7_75t_L g1900 ( .A(n_1147), .B(n_1901), .C(n_1902), .Y(n_1900) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
BUFx3_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
NAND3xp33_ASAP7_75t_L g1274 ( .A(n_1160), .B(n_1275), .C(n_1278), .Y(n_1274) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1175), .Y(n_1225) );
NAND4xp25_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1206), .C(n_1214), .D(n_1220), .Y(n_1197) );
INVx2_ASAP7_75t_SL g1201 ( .A(n_1202), .Y(n_1201) );
INVx2_ASAP7_75t_L g1363 ( .A(n_1202), .Y(n_1363) );
INVx2_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx2_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AO22x2_ASAP7_75t_L g1227 ( .A1(n_1228), .A2(n_1330), .B1(n_1331), .B2(n_1414), .Y(n_1227) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1228), .Y(n_1414) );
XNOR2xp5_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1282), .Y(n_1228) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1230), .Y(n_1281) );
NAND4xp25_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1235), .C(n_1238), .D(n_1244), .Y(n_1231) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
NAND4xp25_ASAP7_75t_L g1253 ( .A(n_1254), .B(n_1260), .C(n_1267), .D(n_1274), .Y(n_1253) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
INVx2_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
NAND3xp33_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1269), .C(n_1273), .Y(n_1267) );
INVx2_ASAP7_75t_SL g1270 ( .A(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
NAND3xp33_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1290), .C(n_1293), .Y(n_1285) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1318), .Y(n_1309) );
BUFx6f_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1912 ( .A(n_1325), .Y(n_1912) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
OAI22xp33_ASAP7_75t_L g1589 ( .A1(n_1329), .A2(n_1590), .B1(n_1591), .B2(n_1594), .Y(n_1589) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
AOI22xp5_ASAP7_75t_L g1331 ( .A1(n_1332), .A2(n_1375), .B1(n_1376), .B2(n_1413), .Y(n_1331) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1332), .Y(n_1413) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1333), .Y(n_1374) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1364), .Y(n_1354) );
BUFx2_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
NAND3xp33_ASAP7_75t_L g1909 ( .A(n_1357), .B(n_1910), .C(n_1913), .Y(n_1909) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1903 ( .A(n_1367), .Y(n_1903) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1377), .Y(n_1412) );
NAND3xp33_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1392), .C(n_1394), .Y(n_1389) );
NAND4xp25_ASAP7_75t_L g1397 ( .A(n_1398), .B(n_1401), .C(n_1404), .D(n_1408), .Y(n_1397) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1415), .Y(n_1548) );
XOR2x2_ASAP7_75t_SL g1415 ( .A(n_1416), .B(n_1457), .Y(n_1415) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
NAND3x1_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1427), .C(n_1435), .Y(n_1419) );
OAI22xp5_ASAP7_75t_L g1437 ( .A1(n_1438), .A2(n_1439), .B1(n_1441), .B2(n_1442), .Y(n_1437) );
INVx3_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
INVx2_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
AOI22xp5_ASAP7_75t_L g1458 ( .A1(n_1459), .A2(n_1511), .B1(n_1512), .B2(n_1547), .Y(n_1458) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1459), .Y(n_1547) );
NAND3xp33_ASAP7_75t_L g1460 ( .A(n_1461), .B(n_1498), .C(n_1506), .Y(n_1460) );
NOR2xp33_ASAP7_75t_L g1461 ( .A(n_1462), .B(n_1477), .Y(n_1461) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
OAI221xp5_ASAP7_75t_L g1469 ( .A1(n_1470), .A2(n_1471), .B1(n_1472), .B2(n_1473), .C(n_1474), .Y(n_1469) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
OAI33xp33_ASAP7_75t_L g1477 ( .A1(n_1478), .A2(n_1480), .A3(n_1486), .B1(n_1488), .B2(n_1493), .B3(n_1497), .Y(n_1477) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
OAI22xp5_ASAP7_75t_L g1480 ( .A1(n_1481), .A2(n_1482), .B1(n_1483), .B2(n_1485), .Y(n_1480) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
OAI22xp5_ASAP7_75t_L g1860 ( .A1(n_1490), .A2(n_1861), .B1(n_1862), .B2(n_1863), .Y(n_1860) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
BUFx3_ASAP7_75t_L g1855 ( .A(n_1501), .Y(n_1855) );
INVx2_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1513), .Y(n_1546) );
NAND2xp5_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1531), .Y(n_1525) );
OAI221xp5_ASAP7_75t_L g1549 ( .A1(n_1550), .A2(n_1781), .B1(n_1782), .B2(n_1870), .C(n_1875), .Y(n_1549) );
NOR4xp25_ASAP7_75t_L g1550 ( .A(n_1551), .B(n_1645), .C(n_1731), .D(n_1758), .Y(n_1550) );
O2A1O1Ixp33_ASAP7_75t_L g1551 ( .A1(n_1552), .A2(n_1582), .B(n_1603), .C(n_1637), .Y(n_1551) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
OAI211xp5_ASAP7_75t_L g1729 ( .A1(n_1553), .A2(n_1624), .B(n_1661), .C(n_1730), .Y(n_1729) );
AOI21xp5_ASAP7_75t_L g1756 ( .A1(n_1553), .A2(n_1609), .B(n_1676), .Y(n_1756) );
NAND2xp5_ASAP7_75t_L g1761 ( .A(n_1553), .B(n_1762), .Y(n_1761) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1573), .Y(n_1553) );
CKINVDCx5p33_ASAP7_75t_R g1610 ( .A(n_1554), .Y(n_1610) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_1554), .B(n_1579), .Y(n_1669) );
AND2x2_ASAP7_75t_L g1690 ( .A(n_1554), .B(n_1613), .Y(n_1690) );
NOR2xp33_ASAP7_75t_L g1700 ( .A(n_1554), .B(n_1701), .Y(n_1700) );
OR2x2_ASAP7_75t_L g1704 ( .A(n_1554), .B(n_1705), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1717 ( .A(n_1554), .B(n_1701), .Y(n_1717) );
NOR2xp33_ASAP7_75t_L g1727 ( .A(n_1554), .B(n_1663), .Y(n_1727) );
AND2x2_ASAP7_75t_L g1733 ( .A(n_1554), .B(n_1641), .Y(n_1733) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1554), .B(n_1673), .Y(n_1739) );
AND2x2_ASAP7_75t_L g1769 ( .A(n_1554), .B(n_1664), .Y(n_1769) );
AND2x4_ASAP7_75t_SL g1554 ( .A(n_1555), .B(n_1567), .Y(n_1554) );
AND2x4_ASAP7_75t_L g1556 ( .A(n_1557), .B(n_1562), .Y(n_1556) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
OR2x2_ASAP7_75t_L g1593 ( .A(n_1558), .B(n_1563), .Y(n_1593) );
NAND2xp5_ASAP7_75t_L g1558 ( .A(n_1559), .B(n_1561), .Y(n_1558) );
HB1xp67_ASAP7_75t_L g1931 ( .A(n_1559), .Y(n_1931) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1561), .Y(n_1571) );
AND2x4_ASAP7_75t_L g1564 ( .A(n_1562), .B(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
OR2x2_ASAP7_75t_L g1596 ( .A(n_1563), .B(n_1566), .Y(n_1596) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1566), .Y(n_1565) );
AND2x2_ASAP7_75t_L g1568 ( .A(n_1569), .B(n_1570), .Y(n_1568) );
AND2x4_ASAP7_75t_L g1572 ( .A(n_1569), .B(n_1571), .Y(n_1572) );
AND2x4_ASAP7_75t_L g1586 ( .A(n_1569), .B(n_1570), .Y(n_1586) );
HB1xp67_ASAP7_75t_L g1929 ( .A(n_1570), .Y(n_1929) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx2_ASAP7_75t_L g1588 ( .A(n_1572), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1634 ( .A(n_1573), .B(n_1610), .Y(n_1634) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1573), .Y(n_1689) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_1573), .B(n_1690), .Y(n_1714) );
AOI22xp33_ASAP7_75t_L g1779 ( .A1(n_1573), .A2(n_1638), .B1(n_1697), .B2(n_1780), .Y(n_1779) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_1574), .B(n_1578), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1641 ( .A(n_1574), .B(n_1579), .Y(n_1641) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1574), .Y(n_1701) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1621 ( .A(n_1575), .B(n_1622), .Y(n_1621) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_1575), .B(n_1579), .Y(n_1673) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_1576), .B(n_1577), .Y(n_1575) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
INVxp67_ASAP7_75t_SL g1622 ( .A(n_1579), .Y(n_1622) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1579), .Y(n_1664) );
AND2x2_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1581), .Y(n_1579) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1582), .Y(n_1707) );
NAND2xp5_ASAP7_75t_L g1582 ( .A(n_1583), .B(n_1597), .Y(n_1582) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1583), .Y(n_1648) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1584), .Y(n_1583) );
BUFx3_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1586), .Y(n_1600) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1587), .Y(n_1781) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
OAI22xp5_ASAP7_75t_SL g1599 ( .A1(n_1588), .A2(n_1600), .B1(n_1601), .B2(n_1602), .Y(n_1599) );
INVx2_ASAP7_75t_L g1615 ( .A(n_1588), .Y(n_1615) );
BUFx3_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
OAI22xp33_ASAP7_75t_L g1616 ( .A1(n_1592), .A2(n_1617), .B1(n_1618), .B2(n_1619), .Y(n_1616) );
BUFx6f_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
HB1xp67_ASAP7_75t_L g1619 ( .A(n_1596), .Y(n_1619) );
CKINVDCx6p67_ASAP7_75t_R g1657 ( .A(n_1597), .Y(n_1657) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_1597), .B(n_1667), .Y(n_1671) );
OR2x2_ASAP7_75t_L g1698 ( .A(n_1597), .B(n_1667), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1597), .B(n_1627), .Y(n_1721) );
OR2x2_ASAP7_75t_L g1728 ( .A(n_1597), .B(n_1642), .Y(n_1728) );
OR2x6_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1599), .Y(n_1597) );
OR2x2_ASAP7_75t_L g1661 ( .A(n_1598), .B(n_1599), .Y(n_1661) );
OAI22xp5_ASAP7_75t_L g1603 ( .A1(n_1604), .A2(n_1623), .B1(n_1630), .B2(n_1635), .Y(n_1603) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1605), .B(n_1609), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1706 ( .A(n_1605), .B(n_1613), .Y(n_1706) );
A2O1A1Ixp33_ASAP7_75t_L g1753 ( .A1(n_1605), .A2(n_1667), .B(n_1754), .C(n_1756), .Y(n_1753) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1606), .Y(n_1625) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1606), .Y(n_1631) );
NAND2xp5_ASAP7_75t_L g1642 ( .A(n_1606), .B(n_1626), .Y(n_1642) );
AND2x2_ASAP7_75t_L g1644 ( .A(n_1606), .B(n_1627), .Y(n_1644) );
AND2x2_ASAP7_75t_L g1656 ( .A(n_1606), .B(n_1657), .Y(n_1656) );
OAI321xp33_ASAP7_75t_L g1692 ( .A1(n_1606), .A2(n_1646), .A3(n_1693), .B1(n_1695), .B2(n_1696), .C(n_1702), .Y(n_1692) );
NAND3xp33_ASAP7_75t_L g1713 ( .A(n_1606), .B(n_1697), .C(n_1714), .Y(n_1713) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1607), .B(n_1608), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1610), .B(n_1611), .Y(n_1609) );
OR2x2_ASAP7_75t_L g1639 ( .A(n_1610), .B(n_1640), .Y(n_1639) );
OR2x2_ASAP7_75t_L g1651 ( .A(n_1610), .B(n_1652), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1682 ( .A(n_1610), .B(n_1614), .Y(n_1682) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_1610), .B(n_1621), .Y(n_1694) );
AND2x2_ASAP7_75t_L g1724 ( .A(n_1610), .B(n_1641), .Y(n_1724) );
AND2x2_ASAP7_75t_L g1747 ( .A(n_1610), .B(n_1673), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1755 ( .A(n_1610), .B(n_1654), .Y(n_1755) );
NOR2xp33_ASAP7_75t_L g1611 ( .A(n_1612), .B(n_1620), .Y(n_1611) );
NAND2xp5_ASAP7_75t_L g1640 ( .A(n_1612), .B(n_1641), .Y(n_1640) );
NOR2x1p5_ASAP7_75t_L g1654 ( .A(n_1612), .B(n_1655), .Y(n_1654) );
AND2x2_ASAP7_75t_L g1699 ( .A(n_1612), .B(n_1700), .Y(n_1699) );
AND2x2_ASAP7_75t_L g1718 ( .A(n_1612), .B(n_1624), .Y(n_1718) );
HB1xp67_ASAP7_75t_L g1762 ( .A(n_1612), .Y(n_1762) );
INVx2_ASAP7_75t_SL g1612 ( .A(n_1613), .Y(n_1612) );
BUFx3_ASAP7_75t_L g1633 ( .A(n_1613), .Y(n_1633) );
BUFx2_ASAP7_75t_L g1653 ( .A(n_1613), .Y(n_1653) );
NOR2xp33_ASAP7_75t_L g1776 ( .A(n_1613), .B(n_1625), .Y(n_1776) );
INVx2_ASAP7_75t_SL g1613 ( .A(n_1614), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1614), .B(n_1625), .Y(n_1676) );
OR2x2_ASAP7_75t_L g1652 ( .A(n_1620), .B(n_1653), .Y(n_1652) );
NOR2xp33_ASAP7_75t_L g1763 ( .A(n_1620), .B(n_1764), .Y(n_1763) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1621), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1681 ( .A(n_1621), .B(n_1682), .Y(n_1681) );
AND2x2_ASAP7_75t_L g1712 ( .A(n_1621), .B(n_1690), .Y(n_1712) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
NAND2xp5_ASAP7_75t_SL g1772 ( .A(n_1624), .B(n_1657), .Y(n_1772) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1625), .B(n_1626), .Y(n_1624) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_1625), .B(n_1657), .Y(n_1683) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1625), .B(n_1627), .Y(n_1691) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
BUFx6f_ASAP7_75t_L g1636 ( .A(n_1627), .Y(n_1636) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1627), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1628), .B(n_1629), .Y(n_1627) );
INVxp67_ASAP7_75t_L g1735 ( .A(n_1630), .Y(n_1735) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1631), .B(n_1632), .Y(n_1630) );
INVx3_ASAP7_75t_L g1711 ( .A(n_1631), .Y(n_1711) );
AOI221xp5_ASAP7_75t_L g1744 ( .A1(n_1631), .A2(n_1646), .B1(n_1691), .B2(n_1745), .C(n_1748), .Y(n_1744) );
O2A1O1Ixp33_ASAP7_75t_L g1719 ( .A1(n_1632), .A2(n_1720), .B(n_1721), .C(n_1722), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1633), .B(n_1634), .Y(n_1632) );
NAND2xp5_ASAP7_75t_L g1749 ( .A(n_1633), .B(n_1747), .Y(n_1749) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1633), .Y(n_1771) );
A2O1A1Ixp33_ASAP7_75t_L g1750 ( .A1(n_1635), .A2(n_1699), .B(n_1751), .C(n_1753), .Y(n_1750) );
CKINVDCx14_ASAP7_75t_R g1635 ( .A(n_1636), .Y(n_1635) );
AOI32xp33_ASAP7_75t_L g1740 ( .A1(n_1636), .A2(n_1640), .A3(n_1646), .B1(n_1741), .B2(n_1742), .Y(n_1740) );
OAI21xp5_ASAP7_75t_L g1637 ( .A1(n_1638), .A2(n_1642), .B(n_1643), .Y(n_1637) );
INVx2_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
INVx2_ASAP7_75t_L g1655 ( .A(n_1641), .Y(n_1655) );
INVx2_ASAP7_75t_L g1734 ( .A(n_1642), .Y(n_1734) );
AOI21xp33_ASAP7_75t_L g1777 ( .A1(n_1643), .A2(n_1680), .B(n_1778), .Y(n_1777) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1644), .B(n_1653), .Y(n_1660) );
AOI21xp33_ASAP7_75t_L g1736 ( .A1(n_1644), .A2(n_1737), .B(n_1740), .Y(n_1736) );
OAI211xp5_ASAP7_75t_L g1645 ( .A1(n_1646), .A2(n_1649), .B(n_1678), .C(n_1719), .Y(n_1645) );
INVx3_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
AOI31xp33_ASAP7_75t_L g1758 ( .A1(n_1647), .A2(n_1759), .A3(n_1765), .B(n_1779), .Y(n_1758) );
INVx2_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
NAND2xp5_ASAP7_75t_L g1695 ( .A(n_1648), .B(n_1657), .Y(n_1695) );
NAND2xp5_ASAP7_75t_L g1743 ( .A(n_1648), .B(n_1667), .Y(n_1743) );
O2A1O1Ixp33_ASAP7_75t_L g1649 ( .A1(n_1650), .A2(n_1654), .B(n_1656), .C(n_1658), .Y(n_1649) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1651), .Y(n_1650) );
NAND2xp5_ASAP7_75t_L g1745 ( .A(n_1652), .B(n_1746), .Y(n_1745) );
OR2x2_ASAP7_75t_L g1668 ( .A(n_1653), .B(n_1669), .Y(n_1668) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_1653), .B(n_1673), .Y(n_1672) );
NAND2xp5_ASAP7_75t_L g1726 ( .A(n_1653), .B(n_1727), .Y(n_1726) );
INVx2_ASAP7_75t_L g1730 ( .A(n_1653), .Y(n_1730) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1654), .Y(n_1773) );
AOI221xp5_ASAP7_75t_L g1679 ( .A1(n_1656), .A2(n_1680), .B1(n_1683), .B2(n_1684), .C(n_1686), .Y(n_1679) );
CKINVDCx5p33_ASAP7_75t_R g1770 ( .A(n_1656), .Y(n_1770) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1657), .B(n_1667), .Y(n_1666) );
AOI31xp33_ASAP7_75t_L g1686 ( .A1(n_1657), .A2(n_1687), .A3(n_1690), .B(n_1691), .Y(n_1686) );
AND2x2_ASAP7_75t_L g1766 ( .A(n_1657), .B(n_1691), .Y(n_1766) );
OAI321xp33_ASAP7_75t_L g1658 ( .A1(n_1659), .A2(n_1661), .A3(n_1662), .B1(n_1665), .B2(n_1668), .C(n_1670), .Y(n_1658) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
NOR3xp33_ASAP7_75t_L g1674 ( .A(n_1661), .B(n_1675), .C(n_1677), .Y(n_1674) );
OAI211xp5_ASAP7_75t_L g1715 ( .A1(n_1661), .A2(n_1716), .B(n_1717), .C(n_1718), .Y(n_1715) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
OAI221xp5_ASAP7_75t_SL g1722 ( .A1(n_1665), .A2(n_1684), .B1(n_1723), .B2(n_1728), .C(n_1729), .Y(n_1722) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
INVx1_ASAP7_75t_L g1775 ( .A(n_1669), .Y(n_1775) );
AOI21xp5_ASAP7_75t_L g1670 ( .A1(n_1671), .A2(n_1672), .B(n_1674), .Y(n_1670) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1671), .Y(n_1709) );
AOI211xp5_ASAP7_75t_L g1765 ( .A1(n_1672), .A2(n_1766), .B(n_1767), .C(n_1777), .Y(n_1765) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1673), .Y(n_1677) );
OAI211xp5_ASAP7_75t_L g1702 ( .A1(n_1673), .A2(n_1703), .B(n_1706), .C(n_1707), .Y(n_1702) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1676), .Y(n_1675) );
OR2x2_ASAP7_75t_L g1684 ( .A(n_1677), .B(n_1685), .Y(n_1684) );
NAND2xp5_ASAP7_75t_L g1688 ( .A(n_1677), .B(n_1689), .Y(n_1688) );
NOR3xp33_ASAP7_75t_SL g1678 ( .A(n_1679), .B(n_1692), .C(n_1708), .Y(n_1678) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
AND2x2_ASAP7_75t_L g1720 ( .A(n_1681), .B(n_1711), .Y(n_1720) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1682), .Y(n_1685) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
AOI21xp5_ASAP7_75t_L g1759 ( .A1(n_1691), .A2(n_1760), .B(n_1763), .Y(n_1759) );
NAND2xp5_ASAP7_75t_L g1737 ( .A(n_1693), .B(n_1738), .Y(n_1737) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1695), .Y(n_1757) );
NAND2xp5_ASAP7_75t_L g1696 ( .A(n_1697), .B(n_1699), .Y(n_1696) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1698), .Y(n_1697) );
HB1xp67_ASAP7_75t_L g1716 ( .A(n_1700), .Y(n_1716) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1701), .Y(n_1705) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
OAI211xp5_ASAP7_75t_L g1708 ( .A1(n_1709), .A2(n_1710), .B(n_1713), .C(n_1715), .Y(n_1708) );
NAND2xp5_ASAP7_75t_L g1710 ( .A(n_1711), .B(n_1712), .Y(n_1710) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1711), .Y(n_1752) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1714), .Y(n_1778) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1718), .Y(n_1764) );
AOI21xp5_ASAP7_75t_L g1732 ( .A1(n_1720), .A2(n_1733), .B(n_1734), .Y(n_1732) );
NOR2xp33_ASAP7_75t_L g1723 ( .A(n_1724), .B(n_1725), .Y(n_1723) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1724), .Y(n_1741) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1726), .Y(n_1725) );
INVx1_ASAP7_75t_L g1780 ( .A(n_1728), .Y(n_1780) );
AOI321xp33_ASAP7_75t_L g1731 ( .A1(n_1732), .A2(n_1735), .A3(n_1736), .B1(n_1744), .B2(n_1750), .C(n_1757), .Y(n_1731) );
INVx1_ASAP7_75t_L g1738 ( .A(n_1739), .Y(n_1738) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1747), .Y(n_1746) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1752), .Y(n_1751) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
OAI321xp33_ASAP7_75t_L g1767 ( .A1(n_1768), .A2(n_1770), .A3(n_1771), .B1(n_1772), .B2(n_1773), .C(n_1774), .Y(n_1767) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
NAND2xp5_ASAP7_75t_L g1774 ( .A(n_1775), .B(n_1776), .Y(n_1774) );
NAND3xp33_ASAP7_75t_L g1783 ( .A(n_1784), .B(n_1832), .C(n_1839), .Y(n_1783) );
NOR2xp33_ASAP7_75t_L g1784 ( .A(n_1785), .B(n_1802), .Y(n_1784) );
NAND2xp5_ASAP7_75t_L g1785 ( .A(n_1786), .B(n_1796), .Y(n_1785) );
AOI22xp33_ASAP7_75t_L g1786 ( .A1(n_1787), .A2(n_1788), .B1(n_1793), .B2(n_1794), .Y(n_1786) );
OAI221xp5_ASAP7_75t_L g1842 ( .A1(n_1787), .A2(n_1793), .B1(n_1843), .B2(n_1844), .C(n_1845), .Y(n_1842) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1790), .Y(n_1789) );
INVx1_ASAP7_75t_L g1810 ( .A(n_1792), .Y(n_1810) );
CKINVDCx6p67_ASAP7_75t_R g1794 ( .A(n_1795), .Y(n_1794) );
AOI22xp33_ASAP7_75t_L g1796 ( .A1(n_1797), .A2(n_1798), .B1(n_1799), .B2(n_1800), .Y(n_1796) );
CKINVDCx6p67_ASAP7_75t_R g1800 ( .A(n_1801), .Y(n_1800) );
NAND3xp33_ASAP7_75t_SL g1802 ( .A(n_1803), .B(n_1815), .C(n_1828), .Y(n_1802) );
AOI22xp33_ASAP7_75t_L g1803 ( .A1(n_1804), .A2(n_1805), .B1(n_1811), .B2(n_1812), .Y(n_1803) );
AOI22xp33_ASAP7_75t_L g1847 ( .A1(n_1804), .A2(n_1811), .B1(n_1848), .B2(n_1851), .Y(n_1847) );
INVx2_ASAP7_75t_L g1805 ( .A(n_1806), .Y(n_1805) );
INVx2_ASAP7_75t_SL g1807 ( .A(n_1808), .Y(n_1807) );
OR2x6_ASAP7_75t_L g1813 ( .A(n_1808), .B(n_1814), .Y(n_1813) );
INVx1_ASAP7_75t_L g1831 ( .A(n_1808), .Y(n_1831) );
INVx2_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1822), .Y(n_1821) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
INVx1_ASAP7_75t_L g1828 ( .A(n_1829), .Y(n_1828) );
INVx1_ASAP7_75t_L g1829 ( .A(n_1830), .Y(n_1829) );
NAND2xp5_ASAP7_75t_L g1832 ( .A(n_1833), .B(n_1834), .Y(n_1832) );
OR2x6_ASAP7_75t_L g1834 ( .A(n_1835), .B(n_1837), .Y(n_1834) );
OAI31xp33_ASAP7_75t_L g1839 ( .A1(n_1840), .A2(n_1852), .A3(n_1865), .B(n_1868), .Y(n_1839) );
HB1xp67_ASAP7_75t_L g1848 ( .A(n_1849), .Y(n_1848) );
INVx2_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
BUFx8_ASAP7_75t_SL g1868 ( .A(n_1869), .Y(n_1868) );
CKINVDCx14_ASAP7_75t_R g1870 ( .A(n_1871), .Y(n_1870) );
BUFx2_ASAP7_75t_L g1871 ( .A(n_1872), .Y(n_1871) );
INVx1_ASAP7_75t_L g1872 ( .A(n_1873), .Y(n_1872) );
INVx1_ASAP7_75t_L g1873 ( .A(n_1874), .Y(n_1873) );
INVxp33_ASAP7_75t_SL g1876 ( .A(n_1877), .Y(n_1876) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1880), .Y(n_1879) );
INVx1_ASAP7_75t_L g1880 ( .A(n_1881), .Y(n_1880) );
NOR3xp33_ASAP7_75t_L g1881 ( .A(n_1882), .B(n_1895), .C(n_1914), .Y(n_1881) );
AOI31xp33_ASAP7_75t_L g1882 ( .A1(n_1883), .A2(n_1886), .A3(n_1891), .B(n_1894), .Y(n_1882) );
NAND4xp25_ASAP7_75t_L g1895 ( .A(n_1896), .B(n_1900), .C(n_1904), .D(n_1909), .Y(n_1895) );
INVx1_ASAP7_75t_L g1911 ( .A(n_1912), .Y(n_1911) );
INVx1_ASAP7_75t_L g1923 ( .A(n_1924), .Y(n_1923) );
CKINVDCx5p33_ASAP7_75t_R g1924 ( .A(n_1925), .Y(n_1924) );
A2O1A1Ixp33_ASAP7_75t_L g1927 ( .A1(n_1926), .A2(n_1928), .B(n_1930), .C(n_1932), .Y(n_1927) );
INVx1_ASAP7_75t_L g1928 ( .A(n_1929), .Y(n_1928) );
INVx1_ASAP7_75t_L g1930 ( .A(n_1931), .Y(n_1930) );
endmodule