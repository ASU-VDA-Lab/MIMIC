module real_aes_863_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_815;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_0), .B(n_142), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_1), .A2(n_151), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_2), .B(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_3), .B(n_158), .Y(n_221) );
INVx1_ASAP7_75t_L g149 ( .A(n_4), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_5), .B(n_158), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_6), .B(n_162), .Y(n_486) );
INVx1_ASAP7_75t_L g520 ( .A(n_7), .Y(n_520) );
OAI22xp5_ASAP7_75t_SL g806 ( .A1(n_8), .A2(n_807), .B1(n_810), .B2(n_811), .Y(n_806) );
INVx1_ASAP7_75t_L g810 ( .A(n_8), .Y(n_810) );
CKINVDCx16_ASAP7_75t_R g821 ( .A(n_9), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_10), .Y(n_558) );
NAND2xp33_ASAP7_75t_L g159 ( .A(n_11), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g139 ( .A(n_12), .Y(n_139) );
AOI221x1_ASAP7_75t_L g237 ( .A1(n_13), .A2(n_25), .B1(n_142), .B2(n_151), .C(n_238), .Y(n_237) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_14), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_15), .B(n_142), .Y(n_141) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_16), .A2(n_137), .B(n_140), .Y(n_136) );
INVx1_ASAP7_75t_L g495 ( .A(n_17), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_18), .B(n_176), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_19), .B(n_158), .Y(n_185) );
AO21x1_ASAP7_75t_L g216 ( .A1(n_20), .A2(n_142), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g120 ( .A(n_21), .Y(n_120) );
INVx1_ASAP7_75t_L g493 ( .A(n_22), .Y(n_493) );
INVx1_ASAP7_75t_SL g503 ( .A(n_23), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_24), .B(n_143), .Y(n_586) );
NAND2x1_ASAP7_75t_L g207 ( .A(n_26), .B(n_158), .Y(n_207) );
AOI33xp33_ASAP7_75t_L g532 ( .A1(n_27), .A2(n_53), .A3(n_470), .B1(n_475), .B2(n_533), .B3(n_534), .Y(n_532) );
NAND2x1_ASAP7_75t_L g195 ( .A(n_28), .B(n_160), .Y(n_195) );
INVx1_ASAP7_75t_L g552 ( .A(n_29), .Y(n_552) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_30), .A2(n_88), .B(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g163 ( .A(n_30), .B(n_88), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_31), .B(n_478), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_32), .B(n_160), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_33), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_34), .B(n_160), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_35), .A2(n_151), .B(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g148 ( .A(n_36), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g152 ( .A(n_36), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g469 ( .A(n_36), .Y(n_469) );
OR2x6_ASAP7_75t_L g118 ( .A(n_37), .B(n_119), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g819 ( .A(n_37), .B(n_820), .C(n_822), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_38), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_39), .B(n_142), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_40), .B(n_478), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_41), .A2(n_162), .B1(n_169), .B2(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_42), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_43), .B(n_143), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_44), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_45), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_46), .B(n_160), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_47), .B(n_137), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_48), .B(n_143), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_49), .A2(n_151), .B(n_194), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_50), .Y(n_583) );
XOR2xp5_ASAP7_75t_L g124 ( .A(n_51), .B(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_52), .B(n_160), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_54), .B(n_143), .Y(n_544) );
INVx1_ASAP7_75t_L g145 ( .A(n_55), .Y(n_145) );
INVx1_ASAP7_75t_L g155 ( .A(n_55), .Y(n_155) );
AND2x2_ASAP7_75t_L g545 ( .A(n_56), .B(n_176), .Y(n_545) );
AOI221xp5_ASAP7_75t_L g518 ( .A1(n_57), .A2(n_73), .B1(n_467), .B2(n_478), .C(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_58), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_59), .B(n_158), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_60), .B(n_169), .Y(n_560) );
AOI21xp5_ASAP7_75t_SL g466 ( .A1(n_61), .A2(n_467), .B(n_472), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_62), .A2(n_151), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g489 ( .A(n_63), .Y(n_489) );
AO21x1_ASAP7_75t_L g218 ( .A1(n_64), .A2(n_151), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_65), .B(n_142), .Y(n_171) );
INVx1_ASAP7_75t_L g543 ( .A(n_66), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_67), .B(n_142), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_68), .A2(n_467), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g231 ( .A(n_69), .B(n_177), .Y(n_231) );
INVx1_ASAP7_75t_L g147 ( .A(n_70), .Y(n_147) );
INVx1_ASAP7_75t_L g153 ( .A(n_70), .Y(n_153) );
AND2x2_ASAP7_75t_L g199 ( .A(n_71), .B(n_168), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_72), .B(n_478), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g807 ( .A1(n_74), .A2(n_84), .B1(n_808), .B2(n_809), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_74), .Y(n_808) );
AND2x2_ASAP7_75t_L g505 ( .A(n_75), .B(n_168), .Y(n_505) );
INVx1_ASAP7_75t_L g490 ( .A(n_76), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_77), .A2(n_467), .B(n_502), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g584 ( .A1(n_78), .A2(n_467), .B(n_527), .C(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g121 ( .A(n_79), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_79), .B(n_120), .Y(n_823) );
AND2x2_ASAP7_75t_L g167 ( .A(n_80), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_81), .B(n_142), .Y(n_187) );
AND2x2_ASAP7_75t_SL g464 ( .A(n_82), .B(n_168), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_83), .A2(n_467), .B1(n_530), .B2(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g809 ( .A(n_84), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_85), .Y(n_798) );
AND2x2_ASAP7_75t_L g217 ( .A(n_86), .B(n_162), .Y(n_217) );
INVxp33_ASAP7_75t_L g825 ( .A(n_87), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_89), .B(n_160), .Y(n_186) );
AND2x2_ASAP7_75t_L g211 ( .A(n_90), .B(n_168), .Y(n_211) );
INVx1_ASAP7_75t_L g473 ( .A(n_91), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_92), .B(n_158), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_93), .A2(n_151), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_94), .B(n_160), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_95), .A2(n_96), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_95), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_96), .Y(n_127) );
AND2x2_ASAP7_75t_L g536 ( .A(n_97), .B(n_168), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_98), .B(n_158), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_99), .A2(n_550), .B(n_551), .C(n_553), .Y(n_549) );
BUFx2_ASAP7_75t_L g108 ( .A(n_100), .Y(n_108) );
BUFx2_ASAP7_75t_SL g801 ( .A(n_100), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_101), .A2(n_151), .B(n_156), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_102), .B(n_143), .Y(n_476) );
AOI21xp33_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_815), .B(n_824), .Y(n_103) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_123), .B(n_799), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_110), .A2(n_803), .B(n_812), .Y(n_802) );
NOR2xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_122), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g814 ( .A(n_115), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
AND2x6_ASAP7_75t_SL g455 ( .A(n_116), .B(n_118), .Y(n_455) );
OR2x6_ASAP7_75t_SL g790 ( .A(n_116), .B(n_117), .Y(n_790) );
OR2x2_ASAP7_75t_L g797 ( .A(n_116), .B(n_118), .Y(n_797) );
CKINVDCx16_ASAP7_75t_R g822 ( .A(n_116), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
OAI222xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_128), .B1(n_791), .B2(n_792), .C1(n_795), .C2(n_798), .Y(n_123) );
INVx1_ASAP7_75t_L g791 ( .A(n_124), .Y(n_791) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_452), .B1(n_456), .B2(n_790), .Y(n_129) );
INVx2_ASAP7_75t_L g794 ( .A(n_130), .Y(n_794) );
OAI22x1_ASAP7_75t_SL g803 ( .A1(n_130), .A2(n_804), .B1(n_805), .B2(n_806), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_130), .Y(n_804) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_373), .Y(n_130) );
NOR3xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_285), .C(n_325), .Y(n_131) );
OAI221xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_200), .B1(n_249), .B2(n_264), .C(n_267), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_164), .Y(n_134) );
INVx2_ASAP7_75t_L g282 ( .A(n_135), .Y(n_282) );
AND2x2_ASAP7_75t_L g312 ( .A(n_135), .B(n_313), .Y(n_312) );
BUFx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g250 ( .A(n_136), .B(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g257 ( .A(n_136), .B(n_190), .Y(n_257) );
INVx2_ASAP7_75t_L g263 ( .A(n_136), .Y(n_263) );
AND2x2_ASAP7_75t_L g272 ( .A(n_136), .B(n_166), .Y(n_272) );
INVx1_ASAP7_75t_L g288 ( .A(n_136), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_136), .B(n_334), .Y(n_333) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_137), .A2(n_518), .B(n_522), .Y(n_517) );
INVx2_ASAP7_75t_SL g527 ( .A(n_137), .Y(n_527) );
BUFx4f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
AND2x4_ASAP7_75t_L g162 ( .A(n_139), .B(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_139), .B(n_163), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_150), .B(n_162), .Y(n_140) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_148), .Y(n_142) );
INVx1_ASAP7_75t_L g491 ( .A(n_143), .Y(n_491) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
AND2x6_ASAP7_75t_L g160 ( .A(n_144), .B(n_153), .Y(n_160) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g158 ( .A(n_146), .B(n_155), .Y(n_158) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx5_ASAP7_75t_L g161 ( .A(n_148), .Y(n_161) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_148), .Y(n_553) );
AND2x2_ASAP7_75t_L g154 ( .A(n_149), .B(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_149), .Y(n_480) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_154), .Y(n_151) );
BUFx3_ASAP7_75t_L g481 ( .A(n_152), .Y(n_481) );
INVx2_ASAP7_75t_L g471 ( .A(n_153), .Y(n_471) );
AND2x4_ASAP7_75t_L g467 ( .A(n_154), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g475 ( .A(n_155), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_161), .Y(n_156) );
INVxp67_ASAP7_75t_L g496 ( .A(n_158), .Y(n_496) );
INVxp67_ASAP7_75t_L g494 ( .A(n_160), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_161), .A2(n_174), .B(n_175), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_161), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_161), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_161), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_161), .A2(n_220), .B(n_221), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_161), .A2(n_228), .B(n_229), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_161), .A2(n_239), .B(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_161), .A2(n_473), .B(n_474), .C(n_476), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_161), .B(n_162), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_SL g502 ( .A1(n_161), .A2(n_474), .B(n_503), .C(n_504), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_SL g519 ( .A1(n_161), .A2(n_474), .B(n_520), .C(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g530 ( .A(n_161), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_161), .A2(n_474), .B(n_543), .C(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_161), .A2(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_SL g181 ( .A(n_162), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_162), .B(n_223), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_162), .A2(n_466), .B(n_477), .Y(n_465) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_165), .B(n_178), .Y(n_164) );
INVx4_ASAP7_75t_L g253 ( .A(n_165), .Y(n_253) );
AND2x2_ASAP7_75t_L g284 ( .A(n_165), .B(n_191), .Y(n_284) );
AND2x2_ASAP7_75t_L g360 ( .A(n_165), .B(n_334), .Y(n_360) );
NAND2x1p5_ASAP7_75t_L g402 ( .A(n_165), .B(n_190), .Y(n_402) );
INVx5_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_166), .B(n_190), .Y(n_289) );
AND2x2_ASAP7_75t_L g313 ( .A(n_166), .B(n_191), .Y(n_313) );
BUFx2_ASAP7_75t_L g329 ( .A(n_166), .Y(n_329) );
NOR2x1_ASAP7_75t_SL g432 ( .A(n_166), .B(n_334), .Y(n_432) );
OR2x6_ASAP7_75t_L g166 ( .A(n_167), .B(n_170), .Y(n_166) );
INVx3_ASAP7_75t_L g210 ( .A(n_168), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_168), .A2(n_210), .B1(n_549), .B2(n_554), .Y(n_548) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_169), .B(n_557), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_176), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_176), .Y(n_198) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_176), .A2(n_237), .B(n_241), .Y(n_236) );
OA21x2_ASAP7_75t_L g299 ( .A1(n_176), .A2(n_237), .B(n_241), .Y(n_299) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g309 ( .A(n_178), .Y(n_309) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_178), .A2(n_376), .B1(n_378), .B2(n_380), .C(n_385), .Y(n_375) );
AND2x2_ASAP7_75t_L g395 ( .A(n_178), .B(n_288), .Y(n_395) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_190), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g251 ( .A(n_180), .Y(n_251) );
INVx1_ASAP7_75t_L g304 ( .A(n_180), .Y(n_304) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_188), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_181), .B(n_189), .Y(n_188) );
AO21x2_ASAP7_75t_L g334 ( .A1(n_181), .A2(n_182), .B(n_188), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_187), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_190), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g273 ( .A(n_190), .B(n_261), .Y(n_273) );
INVx2_ASAP7_75t_L g315 ( .A(n_190), .Y(n_315) );
AND2x2_ASAP7_75t_L g448 ( .A(n_190), .B(n_263), .Y(n_448) );
INVx4_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_191), .Y(n_305) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_198), .B(n_199), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_197), .Y(n_192) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_198), .A2(n_499), .B(n_505), .Y(n_498) );
NOR3xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_232), .C(n_247), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_212), .Y(n_201) );
INVx2_ASAP7_75t_L g362 ( .A(n_202), .Y(n_362) );
AND2x2_ASAP7_75t_L g407 ( .A(n_202), .B(n_284), .Y(n_407) );
BUFx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g352 ( .A(n_203), .Y(n_352) );
AND2x4_ASAP7_75t_SL g367 ( .A(n_203), .B(n_279), .Y(n_367) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_210), .B(n_211), .Y(n_203) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_204), .A2(n_210), .B(n_211), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_209), .Y(n_204) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_210), .A2(n_225), .B(n_231), .Y(n_224) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_210), .A2(n_225), .B(n_231), .Y(n_244) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_210), .A2(n_539), .B(n_545), .Y(n_538) );
AO21x2_ASAP7_75t_L g568 ( .A1(n_210), .A2(n_539), .B(n_545), .Y(n_568) );
INVx2_ASAP7_75t_L g321 ( .A(n_212), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_212), .B(n_351), .Y(n_377) );
AND2x4_ASAP7_75t_L g410 ( .A(n_212), .B(n_357), .Y(n_410) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_224), .Y(n_212) );
AND2x2_ASAP7_75t_L g248 ( .A(n_213), .B(n_243), .Y(n_248) );
OR2x2_ASAP7_75t_L g278 ( .A(n_213), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_SL g347 ( .A(n_213), .B(n_299), .Y(n_347) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
BUFx2_ASAP7_75t_L g292 ( .A(n_214), .Y(n_292) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g266 ( .A(n_215), .Y(n_266) );
OAI21x1_ASAP7_75t_SL g215 ( .A1(n_216), .A2(n_218), .B(n_222), .Y(n_215) );
INVx1_ASAP7_75t_L g223 ( .A(n_217), .Y(n_223) );
INVx2_ASAP7_75t_L g279 ( .A(n_224), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_226), .B(n_230), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_232), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_242), .Y(n_233) );
AND2x2_ASAP7_75t_L g247 ( .A(n_234), .B(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g320 ( .A(n_234), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g405 ( .A(n_234), .Y(n_405) );
BUFx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x4_ASAP7_75t_L g265 ( .A(n_235), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g384 ( .A(n_235), .B(n_244), .Y(n_384) );
AND2x2_ASAP7_75t_L g388 ( .A(n_235), .B(n_254), .Y(n_388) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g357 ( .A(n_236), .Y(n_357) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_236), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_242), .B(n_265), .Y(n_341) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_245), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_243), .B(n_266), .Y(n_451) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g255 ( .A(n_244), .B(n_246), .Y(n_255) );
AND2x2_ASAP7_75t_L g337 ( .A(n_244), .B(n_299), .Y(n_337) );
AND2x2_ASAP7_75t_L g356 ( .A(n_244), .B(n_245), .Y(n_356) );
BUFx2_ASAP7_75t_L g277 ( .A(n_245), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_245), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
BUFx3_ASAP7_75t_L g254 ( .A(n_246), .Y(n_254) );
INVxp67_ASAP7_75t_L g297 ( .A(n_246), .Y(n_297) );
INVx1_ASAP7_75t_L g270 ( .A(n_248), .Y(n_270) );
AND2x2_ASAP7_75t_L g306 ( .A(n_248), .B(n_277), .Y(n_306) );
NAND2xp33_ASAP7_75t_L g387 ( .A(n_248), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g424 ( .A(n_248), .B(n_425), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_252), .B1(n_255), .B2(n_256), .C(n_258), .Y(n_249) );
AND2x2_ASAP7_75t_L g353 ( .A(n_250), .B(n_253), .Y(n_353) );
AND2x2_ASAP7_75t_SL g372 ( .A(n_250), .B(n_313), .Y(n_372) );
AND2x2_ASAP7_75t_L g390 ( .A(n_250), .B(n_315), .Y(n_390) );
AND2x2_ASAP7_75t_L g445 ( .A(n_250), .B(n_284), .Y(n_445) );
INVx1_ASAP7_75t_L g261 ( .A(n_251), .Y(n_261) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_251), .Y(n_317) );
CKINVDCx16_ASAP7_75t_R g397 ( .A(n_252), .Y(n_397) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_253), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_253), .B(n_304), .Y(n_379) );
AND2x2_ASAP7_75t_L g346 ( .A(n_254), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g382 ( .A(n_254), .Y(n_382) );
AND2x2_ASAP7_75t_L g291 ( .A(n_255), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_255), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g433 ( .A(n_255), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_255), .B(n_357), .Y(n_443) );
AND2x4_ASAP7_75t_L g359 ( .A(n_256), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g430 ( .A(n_257), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
OR2x2_ASAP7_75t_L g301 ( .A(n_262), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g308 ( .A(n_263), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g339 ( .A(n_263), .B(n_313), .Y(n_339) );
AND2x2_ASAP7_75t_L g413 ( .A(n_263), .B(n_334), .Y(n_413) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g361 ( .A(n_265), .B(n_362), .Y(n_361) );
OAI32xp33_ASAP7_75t_L g426 ( .A1(n_265), .A2(n_427), .A3(n_429), .B1(n_430), .B2(n_433), .Y(n_426) );
AND2x4_ASAP7_75t_L g298 ( .A(n_266), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g396 ( .A(n_266), .B(n_299), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .B1(n_274), .B2(n_280), .Y(n_267) );
INVxp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_SL g385 ( .A1(n_269), .A2(n_283), .B(n_386), .C(n_387), .Y(n_385) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g369 ( .A(n_270), .B(n_297), .Y(n_369) );
INVx1_ASAP7_75t_SL g440 ( .A(n_271), .Y(n_440) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
AND2x4_ASAP7_75t_L g343 ( .A(n_273), .B(n_282), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_273), .A2(n_422), .B1(n_423), .B2(n_424), .C(n_426), .Y(n_421) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_278), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OAI22xp33_ASAP7_75t_L g363 ( .A1(n_281), .A2(n_311), .B1(n_364), .B2(n_365), .Y(n_363) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
OAI211xp5_ASAP7_75t_SL g399 ( .A1(n_282), .A2(n_400), .B(n_408), .C(n_421), .Y(n_399) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g319 ( .A(n_284), .B(n_288), .Y(n_319) );
OAI211xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_290), .B(n_293), .C(n_322), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g316 ( .A(n_288), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g436 ( .A(n_288), .B(n_432), .Y(n_436) );
OAI32xp33_ASAP7_75t_L g393 ( .A1(n_289), .A2(n_394), .A3(n_396), .B1(n_397), .B2(n_398), .Y(n_393) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_SL g383 ( .A(n_292), .B(n_384), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_300), .B1(n_306), .B2(n_307), .C(n_310), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g450 ( .A(n_297), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_298), .B(n_362), .Y(n_364) );
A2O1A1O1Ixp25_ASAP7_75t_L g435 ( .A1(n_298), .A2(n_367), .B(n_383), .C(n_429), .D(n_436), .Y(n_435) );
AOI31xp33_ASAP7_75t_L g437 ( .A1(n_298), .A2(n_319), .A3(n_429), .B(n_436), .Y(n_437) );
AND2x2_ASAP7_75t_L g351 ( .A(n_299), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_301), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx2_ASAP7_75t_L g428 ( .A(n_303), .Y(n_428) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g423 ( .A(n_304), .B(n_315), .Y(n_423) );
INVx1_ASAP7_75t_L g338 ( .A(n_306), .Y(n_338) );
AND2x2_ASAP7_75t_L g323 ( .A(n_307), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AOI31xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_314), .A3(n_318), .B(n_320), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_313), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g446 ( .A(n_313), .B(n_392), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x2_ASAP7_75t_L g391 ( .A(n_315), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g417 ( .A(n_315), .Y(n_417) );
INVxp67_ASAP7_75t_L g386 ( .A(n_316), .Y(n_386) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g324 ( .A(n_320), .Y(n_324) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND3xp33_ASAP7_75t_SL g325 ( .A(n_326), .B(n_342), .C(n_358), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_335), .B1(n_339), .B2(n_340), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx2_ASAP7_75t_L g412 ( .A(n_329), .Y(n_412) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_333), .Y(n_392) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_333), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_333), .B(n_402), .Y(n_419) );
NAND2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g370 ( .A(n_337), .Y(n_370) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B1(n_353), .B2(n_354), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_345), .B(n_348), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_351), .A2(n_356), .B1(n_390), .B2(n_391), .C(n_393), .Y(n_389) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2x1_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g429 ( .A(n_356), .Y(n_429) );
AND2x2_ASAP7_75t_L g366 ( .A(n_357), .B(n_367), .Y(n_366) );
O2A1O1Ixp33_ASAP7_75t_SL g414 ( .A1(n_357), .A2(n_415), .B(n_419), .C(n_420), .Y(n_414) );
AOI211xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B(n_363), .C(n_368), .Y(n_358) );
AND2x2_ASAP7_75t_L g409 ( .A(n_362), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g420 ( .A(n_367), .Y(n_420) );
AOI21xp33_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_370), .B(n_371), .Y(n_368) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
NOR3xp33_ASAP7_75t_L g373 ( .A(n_374), .B(n_399), .C(n_434), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_375), .B(n_389), .Y(n_374) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g398 ( .A(n_383), .Y(n_398) );
INVxp67_ASAP7_75t_L g422 ( .A(n_387), .Y(n_422) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g406 ( .A(n_396), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B1(n_406), .B2(n_407), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B(n_414), .Y(n_408) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g447 ( .A(n_432), .B(n_448), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_438), .B2(n_441), .C(n_444), .Y(n_434) );
INVxp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI31xp33_ASAP7_75t_SL g444 ( .A1(n_445), .A2(n_446), .A3(n_447), .B(n_449), .Y(n_444) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx4_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx3_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_454), .A2(n_457), .B1(n_790), .B2(n_794), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND3x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_677), .C(n_754), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_629), .Y(n_458) );
NOR2xp67_ASAP7_75t_L g459 ( .A(n_460), .B(n_569), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_506), .B1(n_513), .B2(n_562), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_482), .Y(n_461) );
NOR2xp67_ASAP7_75t_SL g612 ( .A(n_462), .B(n_613), .Y(n_612) );
AND2x4_ASAP7_75t_L g627 ( .A(n_462), .B(n_628), .Y(n_627) );
NOR2x1_ASAP7_75t_L g644 ( .A(n_462), .B(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_SL g684 ( .A(n_462), .B(n_685), .Y(n_684) );
INVx4_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_463), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_463), .B(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g619 ( .A(n_463), .Y(n_619) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_463), .Y(n_624) );
AND2x2_ASAP7_75t_L g653 ( .A(n_463), .B(n_593), .Y(n_653) );
OR2x2_ASAP7_75t_L g657 ( .A(n_463), .B(n_498), .Y(n_657) );
AND2x4_ASAP7_75t_L g670 ( .A(n_463), .B(n_628), .Y(n_670) );
NOR2x1_ASAP7_75t_SL g672 ( .A(n_463), .B(n_485), .Y(n_672) );
AND2x2_ASAP7_75t_L g700 ( .A(n_463), .B(n_578), .Y(n_700) );
OR2x6_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVxp67_ASAP7_75t_L g559 ( .A(n_467), .Y(n_559) );
NOR2x1p5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g534 ( .A(n_470), .Y(n_534) );
INVx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OR2x6_ASAP7_75t_L g474 ( .A(n_471), .B(n_475), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_474), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_488) );
INVxp67_ASAP7_75t_L g550 ( .A(n_474), .Y(n_550) );
INVx2_ASAP7_75t_L g588 ( .A(n_474), .Y(n_588) );
AND2x2_ASAP7_75t_L g479 ( .A(n_475), .B(n_480), .Y(n_479) );
INVxp33_ASAP7_75t_L g533 ( .A(n_475), .Y(n_533) );
INVx1_ASAP7_75t_L g561 ( .A(n_478), .Y(n_561) );
AND2x4_ASAP7_75t_L g478 ( .A(n_479), .B(n_481), .Y(n_478) );
INVx1_ASAP7_75t_L g581 ( .A(n_479), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_481), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_482), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_483), .A2(n_758), .B1(n_760), .B2(n_763), .Y(n_757) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_498), .Y(n_483) );
INVx1_ASAP7_75t_L g512 ( .A(n_484), .Y(n_512) );
AND2x2_ASAP7_75t_L g615 ( .A(n_484), .B(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g620 ( .A(n_484), .B(n_578), .Y(n_620) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g577 ( .A(n_485), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g593 ( .A(n_485), .Y(n_593) );
AND2x2_ASAP7_75t_L g626 ( .A(n_485), .B(n_498), .Y(n_626) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_492), .B(n_497), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_491), .B(n_552), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_492) );
INVx2_ASAP7_75t_L g510 ( .A(n_498), .Y(n_510) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_498), .Y(n_595) );
INVx1_ASAP7_75t_L g614 ( .A(n_498), .Y(n_614) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_498), .Y(n_683) );
INVx1_ASAP7_75t_L g695 ( .A(n_498), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OAI31xp33_ASAP7_75t_SL g749 ( .A1(n_507), .A2(n_750), .A3(n_751), .B(n_752), .Y(n_749) );
NOR2x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_511), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g674 ( .A(n_509), .B(n_576), .Y(n_674) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g590 ( .A(n_510), .Y(n_590) );
AND2x4_ASAP7_75t_SL g710 ( .A(n_512), .B(n_614), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_513), .A2(n_631), .B(n_634), .Y(n_630) );
OR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_523), .Y(n_513) );
INVx2_ASAP7_75t_L g603 ( .A(n_514), .Y(n_603) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2x1p5_ASAP7_75t_L g730 ( .A(n_515), .B(n_638), .Y(n_730) );
BUFx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g640 ( .A(n_516), .B(n_546), .Y(n_640) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVxp67_ASAP7_75t_L g565 ( .A(n_517), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_517), .B(n_526), .Y(n_600) );
AND2x4_ASAP7_75t_L g610 ( .A(n_517), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g655 ( .A(n_517), .B(n_547), .Y(n_655) );
INVx2_ASAP7_75t_L g663 ( .A(n_517), .Y(n_663) );
INVx1_ASAP7_75t_L g762 ( .A(n_517), .Y(n_762) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_517), .Y(n_771) );
INVx1_ASAP7_75t_L g708 ( .A(n_523), .Y(n_708) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_524), .B(n_537), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g564 ( .A(n_525), .B(n_565), .Y(n_564) );
AND2x4_ASAP7_75t_L g703 ( .A(n_525), .B(n_638), .Y(n_703) );
AND2x2_ASAP7_75t_L g720 ( .A(n_525), .B(n_538), .Y(n_720) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_526), .B(n_568), .Y(n_743) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_536), .Y(n_526) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_527), .A2(n_528), .B(n_536), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_529), .B(n_535), .Y(n_528) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g666 ( .A(n_537), .B(n_564), .Y(n_666) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_546), .Y(n_537) );
INVx2_ASAP7_75t_L g572 ( .A(n_538), .Y(n_572) );
NOR2xp67_ASAP7_75t_L g753 ( .A(n_538), .B(n_546), .Y(n_753) );
NOR2x1_ASAP7_75t_L g761 ( .A(n_538), .B(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
AND2x2_ASAP7_75t_L g669 ( .A(n_546), .B(n_573), .Y(n_669) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_547), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g598 ( .A(n_547), .Y(n_598) );
AND2x4_ASAP7_75t_L g662 ( .A(n_547), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g692 ( .A(n_547), .Y(n_692) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_555), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_559), .B1(n_560), .B2(n_561), .Y(n_555) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_563), .A2(n_576), .B1(n_714), .B2(n_715), .C(n_716), .Y(n_713) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
AND2x2_ASAP7_75t_L g690 ( .A(n_564), .B(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_L g733 ( .A(n_564), .Y(n_733) );
INVx2_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g676 ( .A(n_567), .B(n_600), .Y(n_676) );
INVx3_ASAP7_75t_L g638 ( .A(n_568), .Y(n_638) );
AND2x2_ASAP7_75t_L g770 ( .A(n_568), .B(n_771), .Y(n_770) );
NAND3xp33_ASAP7_75t_SL g569 ( .A(n_570), .B(n_601), .C(n_617), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_574), .B1(n_591), .B2(n_596), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_571), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g701 ( .A(n_571), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g712 ( .A(n_571), .B(n_607), .Y(n_712) );
AND2x2_ASAP7_75t_L g782 ( .A(n_571), .B(n_655), .Y(n_782) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx2_ASAP7_75t_L g611 ( .A(n_573), .Y(n_611) );
INVx1_ASAP7_75t_L g660 ( .A(n_573), .Y(n_660) );
INVxp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI222xp33_ASAP7_75t_L g727 ( .A1(n_575), .A2(n_728), .B1(n_729), .B2(n_731), .C1(n_732), .C2(n_734), .Y(n_727) );
OR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_589), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_576), .B(n_603), .Y(n_602) );
NOR2x1_ASAP7_75t_L g735 ( .A(n_576), .B(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g694 ( .A(n_577), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g750 ( .A(n_577), .B(n_624), .Y(n_750) );
INVx2_ASAP7_75t_L g616 ( .A(n_578), .Y(n_616) );
INVx1_ASAP7_75t_L g628 ( .A(n_578), .Y(n_628) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_578), .Y(n_685) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_584), .Y(n_578) );
NOR3xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .C(n_583), .Y(n_580) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_590), .Y(n_633) );
INVx3_ASAP7_75t_L g652 ( .A(n_590), .Y(n_652) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g718 ( .A(n_592), .Y(n_718) );
NAND2x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g705 ( .A(n_594), .Y(n_705) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_L g706 ( .A(n_597), .Y(n_706) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g607 ( .A(n_598), .Y(n_607) );
AND2x2_ASAP7_75t_L g725 ( .A(n_598), .B(n_610), .Y(n_725) );
AND2x2_ASAP7_75t_L g788 ( .A(n_598), .B(n_720), .Y(n_788) );
AND2x2_ASAP7_75t_L g717 ( .A(n_599), .B(n_637), .Y(n_717) );
INVx1_ASAP7_75t_L g728 ( .A(n_599), .Y(n_728) );
AND2x2_ASAP7_75t_L g745 ( .A(n_599), .B(n_692), .Y(n_745) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_604), .B1(n_608), .B2(n_612), .Y(n_601) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_604), .A2(n_618), .B(n_621), .Y(n_617) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g649 ( .A(n_607), .B(n_610), .Y(n_649) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g752 ( .A(n_610), .B(n_753), .Y(n_752) );
BUFx2_ASAP7_75t_L g715 ( .A(n_613), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_614), .Y(n_643) );
AND2x2_ASAP7_75t_SL g623 ( .A(n_615), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g688 ( .A(n_615), .Y(n_688) );
AND2x2_ASAP7_75t_L g786 ( .A(n_615), .B(n_683), .Y(n_786) );
INVx1_ASAP7_75t_L g741 ( .A(n_616), .Y(n_741) );
INVx1_ASAP7_75t_L g647 ( .A(n_618), .Y(n_647) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx1_ASAP7_75t_L g736 ( .A(n_619), .Y(n_736) );
INVx4_ASAP7_75t_L g645 ( .A(n_620), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_625), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI32xp33_ASAP7_75t_L g716 ( .A1(n_623), .A2(n_717), .A3(n_718), .B1(n_719), .B2(n_720), .Y(n_716) );
AND2x2_ASAP7_75t_L g711 ( .A(n_624), .B(n_626), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_SL g774 ( .A1(n_624), .A2(n_775), .B(n_776), .C(n_778), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AND2x2_ASAP7_75t_SL g739 ( .A(n_626), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g778 ( .A(n_626), .Y(n_778) );
AND2x2_ASAP7_75t_L g632 ( .A(n_627), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g759 ( .A(n_627), .Y(n_759) );
AND2x2_ASAP7_75t_L g765 ( .A(n_627), .B(n_652), .Y(n_765) );
NOR3x1_ASAP7_75t_L g629 ( .A(n_630), .B(n_646), .C(n_664), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_641), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
AND2x2_ASAP7_75t_L g654 ( .A(n_637), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g697 ( .A(n_637), .B(n_662), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_637), .B(n_683), .Y(n_724) );
INVx3_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_645), .B(n_652), .Y(n_751) );
INVx2_ASAP7_75t_L g773 ( .A(n_645), .Y(n_773) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B(n_650), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_647), .A2(n_738), .B1(n_742), .B2(n_744), .C(n_749), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_648), .A2(n_768), .B1(n_769), .B2(n_772), .Y(n_767) );
INVx3_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B1(n_656), .B2(n_658), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
AND2x2_ASAP7_75t_L g696 ( .A(n_652), .B(n_672), .Y(n_696) );
INVx1_ASAP7_75t_L g702 ( .A(n_652), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_652), .B(n_670), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_655), .B(n_723), .Y(n_789) );
NAND2x1_ASAP7_75t_L g772 ( .A(n_656), .B(n_773), .Y(n_772) );
INVx2_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_657), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2x1_ASAP7_75t_SL g775 ( .A(n_660), .B(n_662), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_660), .B(n_760), .Y(n_781) );
OR2x2_ASAP7_75t_L g742 ( .A(n_661), .B(n_743), .Y(n_742) );
INVx3_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g777 ( .A(n_662), .B(n_703), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_665), .B(n_671), .Y(n_664) );
OAI21xp33_ASAP7_75t_SL g665 ( .A1(n_666), .A2(n_667), .B(n_670), .Y(n_665) );
OR2x2_ASAP7_75t_L g729 ( .A(n_668), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g763 ( .A(n_669), .B(n_761), .Y(n_763) );
AND2x2_ASAP7_75t_SL g709 ( .A(n_670), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g719 ( .A(n_670), .Y(n_719) );
OAI21xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B(n_675), .Y(n_671) );
AND2x2_ASAP7_75t_L g704 ( .A(n_672), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_721), .Y(n_678) );
NOR3xp33_ASAP7_75t_SL g679 ( .A(n_680), .B(n_698), .C(n_713), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_686), .B(n_689), .C(n_693), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
BUFx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g747 ( .A(n_692), .Y(n_747) );
AND2x2_ASAP7_75t_L g760 ( .A(n_692), .B(n_761), .Y(n_760) );
OAI21xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B(n_697), .Y(n_693) );
INVx1_ASAP7_75t_L g768 ( .A(n_694), .Y(n_768) );
OAI21xp5_ASAP7_75t_SL g698 ( .A1(n_699), .A2(n_706), .B(n_707), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_703), .B2(n_704), .Y(n_699) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_700), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_709), .B1(n_711), .B2(n_712), .Y(n_707) );
INVx1_ASAP7_75t_SL g714 ( .A(n_712), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_718), .B(n_759), .Y(n_758) );
OAI22xp33_ASAP7_75t_SL g784 ( .A1(n_719), .A2(n_785), .B1(n_787), .B2(n_789), .Y(n_784) );
AOI211x1_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_726), .B(n_727), .C(n_737), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
OAI21xp5_ASAP7_75t_L g779 ( .A1(n_739), .A2(n_780), .B(n_782), .Y(n_779) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g748 ( .A(n_743), .Y(n_748) );
NOR2xp67_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_746), .B(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NAND4xp25_ASAP7_75t_L g755 ( .A(n_756), .B(n_766), .C(n_779), .D(n_783), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_764), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_774), .Y(n_766) );
INVxp67_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx2_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
INVx3_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_802), .Y(n_799) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g811 ( .A(n_807), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_SL g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
BUFx4f_ASAP7_75t_SL g827 ( .A(n_818), .Y(n_827) );
NAND2xp5_ASAP7_75t_SL g818 ( .A(n_819), .B(n_823), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
endmodule