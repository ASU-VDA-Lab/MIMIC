module fake_jpeg_16308_n_113 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_113);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_113;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx8_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_19),
.B1(n_24),
.B2(n_23),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_14),
.B1(n_22),
.B2(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_50),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_33),
.Y(n_49)
);

NAND2x1_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_12),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_59),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_34),
.B1(n_31),
.B2(n_26),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_57),
.B1(n_33),
.B2(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_14),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_32),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_72),
.B1(n_3),
.B2(n_7),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_57),
.C(n_48),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_25),
.C(n_20),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_68),
.B(n_3),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_32),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_25),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_56),
.B1(n_54),
.B2(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_55),
.B(n_6),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_78),
.B(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_83),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_81),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_60),
.B1(n_17),
.B2(n_8),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_80),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_9),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_10),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_10),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_68),
.B(n_67),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_92),
.B(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_76),
.C(n_81),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_96),
.C(n_97),
.Y(n_100)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_62),
.B(n_77),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_64),
.C(n_71),
.Y(n_98)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_99),
.A2(n_85),
.B1(n_102),
.B2(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_88),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_104),
.B(n_106),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_89),
.C(n_87),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_100),
.C(n_101),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_109),
.B(n_107),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_110),
.Y(n_113)
);


endmodule