module real_aes_7282_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_532;
wire n_316;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_182;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
INVx1_ASAP7_75t_L g536 ( .A(n_1), .Y(n_536) );
INVx1_ASAP7_75t_L g198 ( .A(n_2), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_3), .A2(n_39), .B1(n_160), .B2(n_478), .Y(n_495) );
AOI21xp33_ASAP7_75t_L g139 ( .A1(n_4), .A2(n_140), .B(n_147), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_5), .B(n_133), .Y(n_527) );
AND2x6_ASAP7_75t_L g145 ( .A(n_6), .B(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_7), .A2(n_239), .B(n_240), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_8), .B(n_41), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_8), .B(n_41), .Y(n_446) );
INVx1_ASAP7_75t_L g157 ( .A(n_9), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_10), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g138 ( .A(n_11), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_12), .B(n_170), .Y(n_473) );
INVx1_ASAP7_75t_L g245 ( .A(n_13), .Y(n_245) );
INVx1_ASAP7_75t_L g531 ( .A(n_14), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_15), .B(n_134), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_16), .A2(n_747), .B1(n_748), .B2(n_751), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_16), .Y(n_751) );
AO32x2_ASAP7_75t_L g493 ( .A1(n_17), .A2(n_133), .A3(n_167), .B1(n_494), .B2(n_498), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_18), .B(n_160), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_19), .B(n_186), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_20), .B(n_134), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_21), .A2(n_52), .B1(n_160), .B2(n_478), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_22), .B(n_140), .Y(n_210) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_23), .A2(n_79), .B1(n_160), .B2(n_170), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_24), .B(n_160), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_25), .B(n_131), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_26), .A2(n_243), .B(n_244), .C(n_246), .Y(n_242) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_27), .A2(n_77), .B1(n_749), .B2(n_750), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_27), .Y(n_750) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_28), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_29), .B(n_163), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_30), .B(n_155), .Y(n_200) );
INVx1_ASAP7_75t_L g176 ( .A(n_31), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_32), .B(n_163), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_33), .B(n_442), .Y(n_450) );
INVx2_ASAP7_75t_L g143 ( .A(n_34), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_35), .B(n_160), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_36), .B(n_163), .Y(n_479) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_37), .A2(n_64), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_37), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_38), .A2(n_145), .B(n_150), .C(n_212), .Y(n_211) );
AOI222xp33_ASAP7_75t_L g452 ( .A1(n_40), .A2(n_453), .B1(n_745), .B2(n_746), .C1(n_752), .C2(n_756), .Y(n_452) );
INVx1_ASAP7_75t_L g174 ( .A(n_42), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_43), .B(n_155), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_44), .B(n_160), .Y(n_521) );
OAI321xp33_ASAP7_75t_L g118 ( .A1(n_45), .A2(n_119), .A3(n_442), .B1(n_447), .B2(n_448), .C(n_450), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_45), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_46), .A2(n_89), .B1(n_217), .B2(n_478), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_47), .B(n_160), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_48), .B(n_160), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_49), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_50), .B(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_51), .B(n_140), .Y(n_233) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_53), .A2(n_62), .B1(n_160), .B2(n_170), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_54), .A2(n_150), .B1(n_170), .B2(n_172), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_55), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_56), .B(n_160), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_57), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_58), .B(n_160), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_59), .A2(n_154), .B(n_156), .C(n_159), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_60), .Y(n_263) );
INVx1_ASAP7_75t_L g148 ( .A(n_61), .Y(n_148) );
INVx1_ASAP7_75t_L g146 ( .A(n_63), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_64), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_65), .B(n_160), .Y(n_537) );
INVx1_ASAP7_75t_L g137 ( .A(n_66), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_67), .Y(n_117) );
AO32x2_ASAP7_75t_L g503 ( .A1(n_68), .A2(n_133), .A3(n_225), .B1(n_498), .B2(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_69), .A2(n_104), .B1(n_112), .B2(n_760), .Y(n_103) );
INVx1_ASAP7_75t_L g548 ( .A(n_70), .Y(n_548) );
INVx1_ASAP7_75t_L g486 ( .A(n_71), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_SL g185 ( .A1(n_72), .A2(n_159), .B(n_186), .C(n_187), .Y(n_185) );
INVxp67_ASAP7_75t_L g188 ( .A(n_73), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_74), .B(n_170), .Y(n_487) );
INVx1_ASAP7_75t_L g111 ( .A(n_75), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_76), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_77), .Y(n_749) );
INVx1_ASAP7_75t_L g256 ( .A(n_78), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_80), .A2(n_145), .B(n_150), .C(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_81), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_82), .B(n_170), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_83), .B(n_199), .Y(n_213) );
INVx2_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_85), .B(n_186), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_86), .B(n_170), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_87), .A2(n_145), .B(n_150), .C(n_197), .Y(n_196) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_88), .B(n_108), .C(n_109), .Y(n_107) );
OR2x2_ASAP7_75t_L g443 ( .A(n_88), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g458 ( .A(n_88), .B(n_445), .Y(n_458) );
INVx2_ASAP7_75t_L g461 ( .A(n_88), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_90), .A2(n_102), .B1(n_170), .B2(n_171), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_91), .B(n_163), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_92), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_93), .A2(n_145), .B(n_150), .C(n_228), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_94), .Y(n_235) );
INVx1_ASAP7_75t_L g184 ( .A(n_95), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g241 ( .A(n_96), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_97), .B(n_199), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_98), .B(n_170), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_99), .B(n_133), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_100), .B(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_101), .A2(n_140), .B(n_183), .Y(n_182) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
CKINVDCx12_ASAP7_75t_R g761 ( .A(n_105), .Y(n_761) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
AND2x2_ASAP7_75t_L g445 ( .A(n_108), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AO21x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_118), .B(n_451), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_SL g759 ( .A(n_116), .Y(n_759) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_119), .B(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_121), .B1(n_124), .B2(n_441), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_124), .A2(n_463), .B1(n_754), .B2(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx2_ASAP7_75t_L g441 ( .A(n_125), .Y(n_441) );
AND3x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_363), .C(n_408), .Y(n_125) );
NOR4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_286), .C(n_327), .D(n_344), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_190), .B(n_206), .C(n_248), .Y(n_127) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_164), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_129), .B(n_191), .Y(n_190) );
NOR4xp25_ASAP7_75t_L g310 ( .A(n_129), .B(n_304), .C(n_311), .D(n_317), .Y(n_310) );
AND2x2_ASAP7_75t_L g383 ( .A(n_129), .B(n_272), .Y(n_383) );
AND2x2_ASAP7_75t_L g402 ( .A(n_129), .B(n_348), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_129), .B(n_397), .Y(n_411) );
AND2x2_ASAP7_75t_L g424 ( .A(n_129), .B(n_205), .Y(n_424) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_SL g269 ( .A(n_130), .Y(n_269) );
AND2x2_ASAP7_75t_L g276 ( .A(n_130), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g326 ( .A(n_130), .B(n_165), .Y(n_326) );
AND2x2_ASAP7_75t_SL g337 ( .A(n_130), .B(n_272), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_130), .B(n_165), .Y(n_341) );
AND2x2_ASAP7_75t_L g350 ( .A(n_130), .B(n_275), .Y(n_350) );
BUFx2_ASAP7_75t_L g373 ( .A(n_130), .Y(n_373) );
AND2x2_ASAP7_75t_L g377 ( .A(n_130), .B(n_181), .Y(n_377) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_139), .B(n_162), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2xp33_ASAP7_75t_SL g219 ( .A(n_132), .B(n_220), .Y(n_219) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_132), .B(n_498), .C(n_514), .Y(n_513) );
AO21x1_ASAP7_75t_L g551 ( .A1(n_132), .A2(n_514), .B(n_552), .Y(n_551) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_133), .A2(n_182), .B(n_189), .Y(n_181) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_133), .A2(n_519), .B(n_527), .Y(n_518) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g167 ( .A(n_134), .Y(n_167) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_135), .B(n_136), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx2_ASAP7_75t_L g239 ( .A(n_140), .Y(n_239) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_141), .B(n_145), .Y(n_178) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g526 ( .A(n_142), .Y(n_526) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
INVx1_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
INVx1_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
INVx3_ASAP7_75t_L g158 ( .A(n_144), .Y(n_158) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_144), .Y(n_173) );
INVx1_ASAP7_75t_L g186 ( .A(n_144), .Y(n_186) );
INVx4_ASAP7_75t_SL g161 ( .A(n_145), .Y(n_161) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_145), .A2(n_471), .B(n_475), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_145), .A2(n_485), .B(n_488), .Y(n_484) );
BUFx3_ASAP7_75t_L g498 ( .A(n_145), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_145), .A2(n_520), .B(n_523), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_145), .A2(n_530), .B(n_534), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_153), .C(n_161), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_149), .A2(n_161), .B(n_184), .C(n_185), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_149), .A2(n_161), .B(n_241), .C(n_242), .Y(n_240) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_151), .Y(n_160) );
BUFx3_ASAP7_75t_L g217 ( .A(n_151), .Y(n_217) );
INVx1_ASAP7_75t_L g478 ( .A(n_151), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_154), .A2(n_476), .B(n_477), .Y(n_475) );
O2A1O1Ixp5_ASAP7_75t_L g547 ( .A1(n_154), .A2(n_535), .B(n_548), .C(n_549), .Y(n_547) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx4_ASAP7_75t_L g231 ( .A(n_155), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_155), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_494) );
OAI22xp5_ASAP7_75t_SL g504 ( .A1(n_155), .A2(n_158), .B1(n_505), .B2(n_506), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_155), .A2(n_496), .B1(n_515), .B2(n_516), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_158), .B(n_188), .Y(n_187) );
INVx5_ASAP7_75t_L g199 ( .A(n_158), .Y(n_199) );
O2A1O1Ixp5_ASAP7_75t_SL g485 ( .A1(n_159), .A2(n_199), .B(n_486), .C(n_487), .Y(n_485) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_160), .Y(n_232) );
OAI22xp33_ASAP7_75t_L g168 ( .A1(n_161), .A2(n_169), .B1(n_177), .B2(n_178), .Y(n_168) );
INVx1_ASAP7_75t_L g204 ( .A(n_163), .Y(n_204) );
INVx2_ASAP7_75t_L g225 ( .A(n_163), .Y(n_225) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_163), .A2(n_238), .B(n_247), .Y(n_237) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_163), .A2(n_470), .B(n_479), .Y(n_469) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_163), .A2(n_484), .B(n_491), .Y(n_483) );
OR2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_181), .Y(n_164) );
AND2x2_ASAP7_75t_L g205 ( .A(n_165), .B(n_181), .Y(n_205) );
BUFx2_ASAP7_75t_L g279 ( .A(n_165), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_165), .A2(n_312), .B1(n_314), .B2(n_315), .Y(n_311) );
OR2x2_ASAP7_75t_L g333 ( .A(n_165), .B(n_193), .Y(n_333) );
AND2x2_ASAP7_75t_L g397 ( .A(n_165), .B(n_275), .Y(n_397) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g265 ( .A(n_166), .B(n_193), .Y(n_265) );
AND2x2_ASAP7_75t_L g272 ( .A(n_166), .B(n_181), .Y(n_272) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_166), .Y(n_314) );
OR2x2_ASAP7_75t_L g349 ( .A(n_166), .B(n_192), .Y(n_349) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_179), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_167), .B(n_180), .Y(n_179) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_167), .A2(n_194), .B(n_202), .Y(n_193) );
INVx2_ASAP7_75t_L g218 ( .A(n_167), .Y(n_218) );
INVx2_ASAP7_75t_L g201 ( .A(n_170), .Y(n_201) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI22xp5_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B1(n_175), .B2(n_176), .Y(n_172) );
INVx2_ASAP7_75t_L g175 ( .A(n_173), .Y(n_175) );
INVx4_ASAP7_75t_L g243 ( .A(n_173), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_178), .A2(n_195), .B(n_196), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_178), .A2(n_256), .B(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g268 ( .A(n_181), .Y(n_268) );
INVx3_ASAP7_75t_L g277 ( .A(n_181), .Y(n_277) );
BUFx2_ASAP7_75t_L g301 ( .A(n_181), .Y(n_301) );
AND2x2_ASAP7_75t_L g334 ( .A(n_181), .B(n_269), .Y(n_334) );
INVx1_ASAP7_75t_L g474 ( .A(n_186), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_190), .A2(n_420), .B1(n_421), .B2(n_422), .Y(n_419) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_205), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_192), .B(n_277), .Y(n_281) );
INVx1_ASAP7_75t_L g309 ( .A(n_192), .Y(n_309) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx3_ASAP7_75t_L g275 ( .A(n_193), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .C(n_201), .Y(n_197) );
INVx2_ASAP7_75t_L g496 ( .A(n_199), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_199), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_199), .A2(n_545), .B(n_546), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_201), .A2(n_531), .B(n_532), .C(n_533), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_204), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_204), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g287 ( .A(n_205), .Y(n_287) );
NAND2x1_ASAP7_75t_SL g206 ( .A(n_207), .B(n_221), .Y(n_206) );
AND2x2_ASAP7_75t_L g285 ( .A(n_207), .B(n_236), .Y(n_285) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_207), .Y(n_359) );
AND2x2_ASAP7_75t_L g386 ( .A(n_207), .B(n_306), .Y(n_386) );
AND2x2_ASAP7_75t_L g394 ( .A(n_207), .B(n_356), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_207), .B(n_251), .Y(n_421) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g252 ( .A(n_208), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g270 ( .A(n_208), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g291 ( .A(n_208), .Y(n_291) );
INVx1_ASAP7_75t_L g297 ( .A(n_208), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_208), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g330 ( .A(n_208), .B(n_254), .Y(n_330) );
OR2x2_ASAP7_75t_L g368 ( .A(n_208), .B(n_323), .Y(n_368) );
AOI32xp33_ASAP7_75t_L g380 ( .A1(n_208), .A2(n_381), .A3(n_384), .B1(n_385), .B2(n_386), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_208), .B(n_356), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_208), .B(n_316), .Y(n_431) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_219), .Y(n_208) );
AOI21xp5_ASAP7_75t_SL g209 ( .A1(n_210), .A2(n_211), .B(n_218), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_215), .A2(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g246 ( .A(n_217), .Y(n_246) );
INVx1_ASAP7_75t_L g261 ( .A(n_218), .Y(n_261) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_218), .A2(n_529), .B(n_538), .Y(n_528) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_218), .A2(n_543), .B(n_550), .Y(n_542) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g342 ( .A(n_222), .B(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_236), .Y(n_222) );
INVx1_ASAP7_75t_L g304 ( .A(n_223), .Y(n_304) );
AND2x2_ASAP7_75t_L g306 ( .A(n_223), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_223), .B(n_253), .Y(n_323) );
AND2x2_ASAP7_75t_L g356 ( .A(n_223), .B(n_332), .Y(n_356) );
AND2x2_ASAP7_75t_L g393 ( .A(n_223), .B(n_254), .Y(n_393) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g251 ( .A(n_224), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_224), .B(n_253), .Y(n_283) );
AND2x2_ASAP7_75t_L g290 ( .A(n_224), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g331 ( .A(n_224), .B(n_332), .Y(n_331) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_234), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_233), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_232), .Y(n_228) );
INVx2_ASAP7_75t_L g307 ( .A(n_236), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_236), .B(n_253), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_236), .B(n_298), .Y(n_379) );
INVx1_ASAP7_75t_L g401 ( .A(n_236), .Y(n_401) );
INVx1_ASAP7_75t_L g418 ( .A(n_236), .Y(n_418) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g271 ( .A(n_237), .B(n_253), .Y(n_271) );
AND2x2_ASAP7_75t_L g293 ( .A(n_237), .B(n_254), .Y(n_293) );
INVx1_ASAP7_75t_L g332 ( .A(n_237), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_243), .B(n_245), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_243), .A2(n_489), .B(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g533 ( .A(n_243), .Y(n_533) );
AOI221x1_ASAP7_75t_SL g248 ( .A1(n_249), .A2(n_264), .B1(n_270), .B2(n_272), .C(n_273), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_249), .A2(n_337), .B1(n_404), .B2(n_405), .Y(n_403) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_252), .Y(n_249) );
AND2x2_ASAP7_75t_L g295 ( .A(n_250), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g390 ( .A(n_250), .B(n_270), .Y(n_390) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g346 ( .A(n_251), .B(n_271), .Y(n_346) );
INVx1_ASAP7_75t_L g358 ( .A(n_252), .Y(n_358) );
AND2x2_ASAP7_75t_L g369 ( .A(n_252), .B(n_356), .Y(n_369) );
AND2x2_ASAP7_75t_L g436 ( .A(n_252), .B(n_331), .Y(n_436) );
INVx2_ASAP7_75t_L g298 ( .A(n_253), .Y(n_298) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_261), .B(n_262), .Y(n_254) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_265), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g388 ( .A(n_265), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_266), .B(n_349), .Y(n_352) );
INVx3_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_267), .A2(n_388), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NOR2xp33_ASAP7_75t_SL g410 ( .A(n_270), .B(n_296), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_271), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g362 ( .A(n_271), .B(n_290), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_271), .B(n_297), .Y(n_439) );
AND2x2_ASAP7_75t_L g308 ( .A(n_272), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g375 ( .A(n_272), .Y(n_375) );
AOI21xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_278), .B(n_282), .Y(n_273) );
NAND2x1_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_275), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g324 ( .A(n_275), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g336 ( .A(n_275), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_275), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g360 ( .A(n_276), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_276), .B(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_276), .B(n_279), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AOI211xp5_ASAP7_75t_L g347 ( .A1(n_279), .A2(n_318), .B(n_348), .C(n_350), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_279), .A2(n_366), .B1(n_369), .B2(n_370), .C(n_374), .Y(n_365) );
AND2x2_ASAP7_75t_L g361 ( .A(n_280), .B(n_314), .Y(n_361) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g321 ( .A(n_285), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g392 ( .A(n_285), .B(n_393), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B(n_294), .C(n_319), .Y(n_286) );
NAND3xp33_ASAP7_75t_SL g405 ( .A(n_287), .B(n_406), .C(n_407), .Y(n_405) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
OR2x2_ASAP7_75t_L g378 ( .A(n_289), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_299), .B1(n_302), .B2(n_308), .C(n_310), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_296), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_296), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g318 ( .A(n_301), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_301), .A2(n_358), .B1(n_359), .B2(n_360), .Y(n_357) );
OR2x2_ASAP7_75t_L g438 ( .A(n_301), .B(n_349), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVxp67_ASAP7_75t_L g412 ( .A(n_304), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_306), .B(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g313 ( .A(n_307), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_309), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_309), .B(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_309), .B(n_376), .Y(n_415) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_313), .Y(n_339) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g429 ( .A(n_318), .B(n_349), .Y(n_429) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_324), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g407 ( .A(n_324), .Y(n_407) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI322xp33_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_333), .A3(n_334), .B1(n_335), .B2(n_338), .C1(n_340), .C2(n_342), .Y(n_327) );
OAI322xp33_ASAP7_75t_L g409 ( .A1(n_328), .A2(n_410), .A3(n_411), .B1(n_412), .B2(n_413), .C1(n_414), .C2(n_416), .Y(n_409) );
CKINVDCx16_ASAP7_75t_R g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx4_ASAP7_75t_L g343 ( .A(n_330), .Y(n_343) );
AND2x2_ASAP7_75t_L g404 ( .A(n_330), .B(n_356), .Y(n_404) );
AND2x2_ASAP7_75t_L g417 ( .A(n_330), .B(n_418), .Y(n_417) );
CKINVDCx16_ASAP7_75t_R g428 ( .A(n_333), .Y(n_428) );
INVx1_ASAP7_75t_L g406 ( .A(n_334), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
OR2x2_ASAP7_75t_L g340 ( .A(n_336), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g423 ( .A(n_336), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_336), .B(n_377), .Y(n_434) );
OR2x2_ASAP7_75t_L g367 ( .A(n_339), .B(n_368), .Y(n_367) );
INVxp33_ASAP7_75t_L g384 ( .A(n_339), .Y(n_384) );
OAI221xp5_ASAP7_75t_SL g344 ( .A1(n_343), .A2(n_345), .B1(n_347), .B2(n_351), .C(n_353), .Y(n_344) );
NOR2xp67_ASAP7_75t_L g400 ( .A(n_343), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g427 ( .A(n_343), .Y(n_427) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx3_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AOI322xp5_ASAP7_75t_L g391 ( .A1(n_350), .A2(n_375), .A3(n_392), .B1(n_394), .B2(n_395), .C1(n_398), .C2(n_402), .Y(n_391) );
INVxp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .B1(n_361), .B2(n_362), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_387), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_365), .B(n_380), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_368), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NAND2xp33_ASAP7_75t_SL g385 ( .A(n_371), .B(n_382), .Y(n_385) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
OAI322xp33_ASAP7_75t_L g425 ( .A1(n_373), .A2(n_426), .A3(n_428), .B1(n_429), .B2(n_430), .C1(n_432), .C2(n_435), .Y(n_425) );
AOI21xp33_ASAP7_75t_SL g374 ( .A1(n_375), .A2(n_376), .B(n_378), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_383), .B(n_431), .Y(n_440) );
OAI211xp5_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_389), .B(n_391), .C(n_403), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NOR4xp25_ASAP7_75t_L g408 ( .A(n_409), .B(n_419), .C(n_425), .D(n_437), .Y(n_408) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
CKINVDCx14_ASAP7_75t_R g435 ( .A(n_436), .Y(n_435) );
OAI21xp5_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_439), .B(n_440), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_441), .A2(n_455), .B1(n_459), .B2(n_462), .Y(n_454) );
INVx1_ASAP7_75t_L g449 ( .A(n_442), .Y(n_449) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NOR2x2_ASAP7_75t_L g758 ( .A(n_444), .B(n_461), .Y(n_758) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g460 ( .A(n_445), .B(n_461), .Y(n_460) );
AOI21xp33_ASAP7_75t_L g451 ( .A1(n_450), .A2(n_452), .B(n_759), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g754 ( .A(n_458), .Y(n_754) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx6_ASAP7_75t_L g755 ( .A(n_460), .Y(n_755) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_667), .Y(n_463) );
NAND5xp2_ASAP7_75t_L g464 ( .A(n_465), .B(n_586), .C(n_601), .D(n_627), .E(n_649), .Y(n_464) );
NOR2xp33_ASAP7_75t_SL g465 ( .A(n_466), .B(n_566), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_507), .B1(n_539), .B2(n_555), .C(n_556), .Y(n_466) );
NOR2xp33_ASAP7_75t_SL g467 ( .A(n_468), .B(n_499), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_468), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g743 ( .A(n_468), .Y(n_743) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_480), .Y(n_468) );
INVx1_ASAP7_75t_L g583 ( .A(n_469), .Y(n_583) );
AND2x2_ASAP7_75t_L g585 ( .A(n_469), .B(n_493), .Y(n_585) );
AND2x2_ASAP7_75t_L g595 ( .A(n_469), .B(n_492), .Y(n_595) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_469), .Y(n_613) );
INVx1_ASAP7_75t_L g623 ( .A(n_469), .Y(n_623) );
OR2x2_ASAP7_75t_L g661 ( .A(n_469), .B(n_560), .Y(n_661) );
INVx2_ASAP7_75t_L g711 ( .A(n_469), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_469), .B(n_559), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_474), .Y(n_471) );
NOR2xp67_ASAP7_75t_L g480 ( .A(n_481), .B(n_492), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_482), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_482), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_SL g643 ( .A(n_482), .B(n_583), .Y(n_643) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_483), .Y(n_501) );
INVx2_ASAP7_75t_L g560 ( .A(n_483), .Y(n_560) );
OR2x2_ASAP7_75t_L g622 ( .A(n_483), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g561 ( .A(n_492), .B(n_503), .Y(n_561) );
AND2x2_ASAP7_75t_L g578 ( .A(n_492), .B(n_558), .Y(n_578) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g502 ( .A(n_493), .B(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g581 ( .A(n_493), .Y(n_581) );
AND2x2_ASAP7_75t_L g710 ( .A(n_493), .B(n_711), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_496), .A2(n_524), .B(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_496), .A2(n_535), .B(n_536), .C(n_537), .Y(n_534) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_498), .A2(n_544), .B(n_547), .Y(n_543) );
INVx1_ASAP7_75t_L g555 ( .A(n_499), .Y(n_555) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
AND2x2_ASAP7_75t_L g673 ( .A(n_500), .B(n_561), .Y(n_673) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g674 ( .A(n_501), .B(n_585), .Y(n_674) );
O2A1O1Ixp33_ASAP7_75t_L g641 ( .A1(n_502), .A2(n_642), .B(n_644), .C(n_646), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_502), .B(n_642), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_502), .A2(n_572), .B1(n_715), .B2(n_716), .C(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g558 ( .A(n_503), .Y(n_558) );
INVx1_ASAP7_75t_L g594 ( .A(n_503), .Y(n_594) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_503), .Y(n_603) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_517), .Y(n_508) );
AND2x2_ASAP7_75t_L g620 ( .A(n_509), .B(n_565), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_509), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_510), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g712 ( .A(n_510), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g744 ( .A(n_510), .Y(n_744) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g574 ( .A(n_511), .Y(n_574) );
AND2x2_ASAP7_75t_L g600 ( .A(n_511), .B(n_554), .Y(n_600) );
NOR2x1_ASAP7_75t_L g609 ( .A(n_511), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g616 ( .A(n_511), .B(n_617), .Y(n_616) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g552 ( .A(n_512), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_517), .B(n_656), .Y(n_691) );
INVx1_ASAP7_75t_SL g695 ( .A(n_517), .Y(n_695) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_528), .Y(n_517) );
INVx3_ASAP7_75t_L g554 ( .A(n_518), .Y(n_554) );
AND2x2_ASAP7_75t_L g565 ( .A(n_518), .B(n_542), .Y(n_565) );
AND2x2_ASAP7_75t_L g587 ( .A(n_518), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g632 ( .A(n_518), .B(n_626), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_518), .B(n_564), .Y(n_713) );
INVx2_ASAP7_75t_L g535 ( .A(n_526), .Y(n_535) );
AND2x2_ASAP7_75t_L g553 ( .A(n_528), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g564 ( .A(n_528), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_528), .B(n_542), .Y(n_589) );
AND2x2_ASAP7_75t_L g625 ( .A(n_528), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_553), .Y(n_540) );
INVx1_ASAP7_75t_L g605 ( .A(n_541), .Y(n_605) );
AND2x2_ASAP7_75t_L g647 ( .A(n_541), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_541), .B(n_568), .Y(n_653) );
AOI21xp5_ASAP7_75t_SL g727 ( .A1(n_541), .A2(n_559), .B(n_582), .Y(n_727) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_551), .Y(n_541) );
OR2x2_ASAP7_75t_L g570 ( .A(n_542), .B(n_551), .Y(n_570) );
AND2x2_ASAP7_75t_L g617 ( .A(n_542), .B(n_554), .Y(n_617) );
INVx2_ASAP7_75t_L g626 ( .A(n_542), .Y(n_626) );
INVx1_ASAP7_75t_L g732 ( .A(n_542), .Y(n_732) );
AND2x2_ASAP7_75t_L g656 ( .A(n_551), .B(n_626), .Y(n_656) );
INVx1_ASAP7_75t_L g681 ( .A(n_551), .Y(n_681) );
AND2x2_ASAP7_75t_L g590 ( .A(n_553), .B(n_574), .Y(n_590) );
AND2x2_ASAP7_75t_L g602 ( .A(n_553), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_SL g720 ( .A(n_553), .Y(n_720) );
INVx2_ASAP7_75t_L g610 ( .A(n_554), .Y(n_610) );
AND2x2_ASAP7_75t_L g648 ( .A(n_554), .B(n_564), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_554), .B(n_732), .Y(n_731) );
OAI21xp33_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_561), .B(n_562), .Y(n_556) );
AND2x2_ASAP7_75t_L g663 ( .A(n_557), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g717 ( .A(n_557), .Y(n_717) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g637 ( .A(n_558), .Y(n_637) );
BUFx2_ASAP7_75t_L g736 ( .A(n_558), .Y(n_736) );
BUFx2_ASAP7_75t_L g607 ( .A(n_559), .Y(n_607) );
AND2x2_ASAP7_75t_L g709 ( .A(n_559), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g692 ( .A(n_560), .Y(n_692) );
AND2x4_ASAP7_75t_L g619 ( .A(n_561), .B(n_582), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_561), .B(n_643), .Y(n_655) );
AOI32xp33_ASAP7_75t_L g579 ( .A1(n_562), .A2(n_580), .A3(n_582), .B1(n_584), .B2(n_585), .Y(n_579) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx3_ASAP7_75t_L g568 ( .A(n_563), .Y(n_568) );
OR2x2_ASAP7_75t_L g704 ( .A(n_563), .B(n_660), .Y(n_704) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g573 ( .A(n_564), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g680 ( .A(n_564), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g572 ( .A(n_565), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g584 ( .A(n_565), .B(n_574), .Y(n_584) );
INVx1_ASAP7_75t_L g705 ( .A(n_565), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_565), .B(n_680), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_571), .B(n_575), .C(n_579), .Y(n_566) );
OAI322xp33_ASAP7_75t_L g675 ( .A1(n_567), .A2(n_612), .A3(n_676), .B1(n_678), .B2(n_682), .C1(n_683), .C2(n_687), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVxp67_ASAP7_75t_L g640 ( .A(n_568), .Y(n_640) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g694 ( .A(n_570), .B(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_570), .B(n_610), .Y(n_741) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g633 ( .A(n_573), .Y(n_633) );
OR2x2_ASAP7_75t_L g719 ( .A(n_574), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_577), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g628 ( .A(n_578), .B(n_607), .Y(n_628) );
AND2x2_ASAP7_75t_L g699 ( .A(n_578), .B(n_612), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_578), .B(n_686), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_580), .A2(n_587), .B1(n_590), .B2(n_591), .C(n_596), .Y(n_586) );
OR2x2_ASAP7_75t_L g597 ( .A(n_580), .B(n_593), .Y(n_597) );
AND2x2_ASAP7_75t_L g685 ( .A(n_580), .B(n_686), .Y(n_685) );
AOI32xp33_ASAP7_75t_L g724 ( .A1(n_580), .A2(n_610), .A3(n_725), .B1(n_726), .B2(n_729), .Y(n_724) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_581), .B(n_617), .C(n_640), .Y(n_658) );
AND2x2_ASAP7_75t_L g684 ( .A(n_581), .B(n_677), .Y(n_684) );
INVxp67_ASAP7_75t_L g664 ( .A(n_582), .Y(n_664) );
BUFx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_585), .B(n_637), .Y(n_693) );
INVx2_ASAP7_75t_L g703 ( .A(n_585), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_585), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g672 ( .A(n_588), .Y(n_672) );
OR2x2_ASAP7_75t_L g598 ( .A(n_589), .B(n_599), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_591), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_594), .Y(n_677) );
AND2x2_ASAP7_75t_L g636 ( .A(n_595), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g682 ( .A(n_595), .Y(n_682) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_595), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AOI21xp33_ASAP7_75t_SL g621 ( .A1(n_597), .A2(n_622), .B(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g715 ( .A(n_600), .B(n_625), .Y(n_715) );
AOI211xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_604), .B(n_614), .C(n_621), .Y(n_601) );
AND2x2_ASAP7_75t_L g645 ( .A(n_603), .B(n_613), .Y(n_645) );
INVx2_ASAP7_75t_L g660 ( .A(n_603), .Y(n_660) );
OR2x2_ASAP7_75t_L g698 ( .A(n_603), .B(n_661), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_603), .B(n_741), .Y(n_740) );
AOI211xp5_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_606), .B(n_608), .C(n_611), .Y(n_604) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_607), .B(n_645), .Y(n_644) );
OAI211xp5_ASAP7_75t_L g726 ( .A1(n_608), .A2(n_703), .B(n_727), .C(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_609), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g666 ( .A(n_610), .B(n_656), .Y(n_666) );
INVx1_ASAP7_75t_L g671 ( .A(n_610), .Y(n_671) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_615), .B(n_618), .Y(n_614) );
INVxp33_ASAP7_75t_L g722 ( .A(n_616), .Y(n_722) );
AND2x2_ASAP7_75t_L g701 ( .A(n_617), .B(n_680), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_622), .A2(n_684), .B(n_685), .Y(n_683) );
OAI322xp33_ASAP7_75t_L g702 ( .A1(n_624), .A2(n_703), .A3(n_704), .B1(n_705), .B2(n_706), .C1(n_708), .C2(n_712), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B1(n_634), .B2(n_638), .C(n_641), .Y(n_627) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g679 ( .A(n_632), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g723 ( .A(n_636), .Y(n_723) );
INVxp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_639), .B(n_659), .Y(n_725) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g688 ( .A(n_648), .B(n_656), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B1(n_654), .B2(n_656), .C(n_657), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_652), .A2(n_669), .B1(n_673), .B2(n_674), .C(n_675), .Y(n_668) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_656), .B(n_671), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B1(n_662), .B2(n_665), .Y(n_657) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx2_ASAP7_75t_SL g686 ( .A(n_661), .Y(n_686) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND5xp2_ASAP7_75t_L g667 ( .A(n_668), .B(n_689), .C(n_714), .D(n_724), .E(n_734), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_670), .B(n_672), .Y(n_669) );
NOR4xp25_ASAP7_75t_L g742 ( .A(n_671), .B(n_677), .C(n_743), .D(n_744), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g734 ( .A1(n_674), .A2(n_735), .B1(n_737), .B2(n_739), .C(n_742), .Y(n_734) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g733 ( .A(n_680), .Y(n_733) );
OAI322xp33_ASAP7_75t_L g690 ( .A1(n_684), .A2(n_691), .A3(n_692), .B1(n_693), .B2(n_694), .C1(n_696), .C2(n_700), .Y(n_690) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_702), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g735 ( .A(n_710), .B(n_736), .Y(n_735) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_721), .B1(n_722), .B2(n_723), .Y(n_718) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
endmodule