module fake_jpeg_1865_n_675 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_675);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_675;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_483;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_650;
wire n_328;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

CKINVDCx6p67_ASAP7_75t_R g154 ( 
.A(n_60),
.Y(n_154)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_61),
.Y(n_170)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_36),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g195 ( 
.A(n_63),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_64),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_65),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_22),
.B(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_66),
.B(n_77),
.Y(n_142)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_69),
.B(n_72),
.Y(n_134)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_19),
.B(n_16),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_73),
.Y(n_178)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_79),
.B(n_86),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_82),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_31),
.B(n_16),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_84),
.B(n_3),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_38),
.B(n_49),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_90),
.Y(n_206)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

CKINVDCx9p33_ASAP7_75t_R g92 ( 
.A(n_54),
.Y(n_92)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_92),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_96),
.Y(n_147)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_53),
.B(n_1),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_40),
.B(n_2),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_32),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_25),
.B(n_2),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_109),
.Y(n_156)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_37),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_110),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_40),
.B(n_3),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_117),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_37),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_114),
.Y(n_210)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_50),
.Y(n_117)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_24),
.Y(n_119)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_24),
.Y(n_120)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_26),
.Y(n_121)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_121),
.Y(n_221)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx5_ASAP7_75t_SL g215 ( 
.A(n_124),
.Y(n_215)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_26),
.Y(n_125)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_54),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_129),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_28),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_28),
.Y(n_128)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_45),
.B(n_3),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_130),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_133),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_63),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_139),
.B(n_149),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_140),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_145),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_146),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_65),
.B(n_44),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_107),
.B(n_44),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_153),
.B(n_163),
.Y(n_286)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_157),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_88),
.B(n_34),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_82),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_175),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_62),
.A2(n_34),
.B1(n_57),
.B2(n_56),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_179),
.A2(n_216),
.B1(n_41),
.B2(n_52),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_70),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_214),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_96),
.B(n_27),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_186),
.A2(n_189),
.B(n_191),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_96),
.B(n_27),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_92),
.B(n_48),
.Y(n_191)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_192),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_194),
.B(n_48),
.Y(n_243)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_61),
.Y(n_197)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_197),
.Y(n_250)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_94),
.B(n_47),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_220),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_67),
.Y(n_209)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_90),
.Y(n_211)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_124),
.A2(n_47),
.B(n_33),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_212),
.B(n_110),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_116),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_114),
.A2(n_33),
.B1(n_51),
.B2(n_56),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_73),
.Y(n_217)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_64),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g303 ( 
.A(n_219),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_122),
.B(n_25),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_64),
.B(n_35),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_4),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_89),
.Y(n_223)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_225),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_195),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_228),
.B(n_244),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_128),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_231),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g232 ( 
.A(n_142),
.B(n_128),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_232),
.B(n_235),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_168),
.B(n_43),
.Y(n_235)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_136),
.Y(n_238)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_238),
.Y(n_314)
);

AND2x2_ASAP7_75t_SL g240 ( 
.A(n_165),
.B(n_105),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_240),
.Y(n_336)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_241),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_191),
.A2(n_43),
.B1(n_35),
.B2(n_41),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_242),
.A2(n_258),
.B1(n_280),
.B2(n_216),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_243),
.B(n_268),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_210),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_198),
.A2(n_144),
.B1(n_173),
.B2(n_51),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_245),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_246),
.A2(n_248),
.B1(n_249),
.B2(n_252),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_144),
.A2(n_51),
.B1(n_33),
.B2(n_57),
.Y(n_248)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_154),
.Y(n_249)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_143),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_251),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_186),
.A2(n_52),
.B1(n_91),
.B2(n_100),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_147),
.B(n_3),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_256),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_154),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_265),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_171),
.A2(n_58),
.B1(n_54),
.B2(n_30),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_148),
.A2(n_30),
.B1(n_54),
.B2(n_58),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_259),
.A2(n_141),
.B1(n_196),
.B2(n_182),
.Y(n_315)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_174),
.Y(n_260)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_260),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_261),
.B(n_151),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_189),
.B(n_4),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_262),
.B(n_266),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_210),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_263),
.B(n_285),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_154),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_148),
.B(n_4),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_168),
.B(n_142),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_147),
.A2(n_205),
.B1(n_213),
.B2(n_221),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g331 ( 
.A1(n_269),
.A2(n_287),
.B1(n_293),
.B2(n_169),
.Y(n_331)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_131),
.Y(n_270)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

HAxp5_ASAP7_75t_SL g271 ( 
.A(n_156),
.B(n_123),
.CON(n_271),
.SN(n_271)
);

NOR2x1_ASAP7_75t_L g322 ( 
.A(n_271),
.B(n_232),
.Y(n_322)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_135),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_272),
.B(n_288),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_274),
.B(n_282),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_177),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_275),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_161),
.A2(n_123),
.B1(n_111),
.B2(n_58),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_276),
.A2(n_299),
.B1(n_193),
.B2(n_141),
.Y(n_310)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_138),
.Y(n_278)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_155),
.Y(n_279)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_161),
.A2(n_58),
.B1(n_54),
.B2(n_111),
.Y(n_280)
);

CKINVDCx12_ASAP7_75t_R g281 ( 
.A(n_215),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_281),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_156),
.B(n_4),
.Y(n_282)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_176),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_283),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_170),
.Y(n_284)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_284),
.Y(n_305)
);

AOI21xp33_ASAP7_75t_L g285 ( 
.A1(n_134),
.A2(n_85),
.B(n_83),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_132),
.A2(n_54),
.B1(n_28),
.B2(n_8),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_172),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_289),
.B(n_296),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_190),
.B(n_5),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_290),
.B(n_291),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_203),
.B(n_5),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_150),
.Y(n_292)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_167),
.A2(n_28),
.B1(n_10),
.B2(n_11),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_207),
.B(n_6),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_301),
.Y(n_325)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_183),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_187),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_297),
.B(n_300),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_206),
.Y(n_298)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_212),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_133),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_222),
.B(n_6),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_162),
.B(n_6),
.C(n_10),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_256),
.Y(n_362)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_164),
.Y(n_304)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_304),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_307),
.B(n_310),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_261),
.A2(n_166),
.B(n_159),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_312),
.B(n_331),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_254),
.A2(n_199),
.B1(n_152),
.B2(n_200),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_313),
.A2(n_315),
.B1(n_326),
.B2(n_330),
.Y(n_394)
);

NOR2x1_ASAP7_75t_L g406 ( 
.A(n_322),
.B(n_338),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_276),
.A2(n_158),
.B(n_181),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_324),
.A2(n_346),
.B(n_226),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_253),
.A2(n_199),
.B1(n_152),
.B2(n_200),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_256),
.B(n_176),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_231),
.C(n_250),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_290),
.A2(n_137),
.B1(n_196),
.B2(n_155),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_247),
.B(n_151),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_334),
.B(n_351),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_253),
.A2(n_137),
.B1(n_182),
.B2(n_201),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_335),
.A2(n_345),
.B1(n_353),
.B2(n_354),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_240),
.B(n_160),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_342),
.Y(n_403)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_291),
.A2(n_178),
.B1(n_202),
.B2(n_184),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_271),
.A2(n_176),
.B(n_188),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_266),
.B(n_201),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_349),
.B(n_363),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_286),
.B(n_160),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_240),
.A2(n_188),
.B1(n_13),
.B2(n_16),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_299),
.A2(n_188),
.B1(n_11),
.B2(n_13),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_237),
.B(n_230),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_355),
.B(n_303),
.Y(n_405)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_270),
.Y(n_358)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_358),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_229),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_360),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_255),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_362),
.B(n_267),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_262),
.B(n_302),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_278),
.B(n_292),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_365),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_225),
.B(n_260),
.Y(n_365)
);

INVx13_ASAP7_75t_L g366 ( 
.A(n_344),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_366),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g367 ( 
.A(n_311),
.B(n_249),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_367),
.B(n_368),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_347),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_356),
.A2(n_233),
.B1(n_284),
.B2(n_298),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_369),
.A2(n_373),
.B(n_397),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_370),
.B(n_317),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_347),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_371),
.B(n_377),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_314),
.Y(n_372)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_356),
.A2(n_233),
.B1(n_273),
.B2(n_231),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_306),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_375),
.B(n_387),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_350),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_365),
.Y(n_378)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_306),
.Y(n_379)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_379),
.Y(n_422)
);

INVx13_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_381),
.Y(n_431)
);

AND2x6_ASAP7_75t_L g382 ( 
.A(n_322),
.B(n_283),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_382),
.B(n_404),
.Y(n_417)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_332),
.A2(n_273),
.B1(n_264),
.B2(n_295),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_384),
.A2(n_385),
.B1(n_392),
.B2(n_326),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_336),
.A2(n_264),
.B1(n_279),
.B2(n_251),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_341),
.Y(n_386)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_386),
.Y(n_428)
);

OA21x2_ASAP7_75t_L g387 ( 
.A1(n_312),
.A2(n_250),
.B(n_277),
.Y(n_387)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_321),
.Y(n_389)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_389),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_309),
.B(n_255),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_390),
.B(n_391),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_348),
.B(n_238),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_348),
.A2(n_241),
.B1(n_295),
.B2(n_267),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_393),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_396),
.B(n_399),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_338),
.A2(n_275),
.B1(n_227),
.B2(n_277),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_362),
.B(n_227),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_341),
.Y(n_400)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_400),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_226),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_405),
.B(n_410),
.Y(n_440)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_308),
.Y(n_407)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_407),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_408),
.A2(n_409),
.B1(n_323),
.B2(n_335),
.Y(n_419)
);

INVx11_ASAP7_75t_L g409 ( 
.A(n_360),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_339),
.B(n_303),
.Y(n_410)
);

OAI22x1_ASAP7_75t_SL g411 ( 
.A1(n_322),
.A2(n_239),
.B1(n_234),
.B2(n_303),
.Y(n_411)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_411),
.A2(n_342),
.B(n_346),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_339),
.B(n_239),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_412),
.B(n_413),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_320),
.B(n_239),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_380),
.A2(n_315),
.B1(n_324),
.B2(n_338),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_415),
.A2(n_420),
.B1(n_423),
.B2(n_376),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_419),
.A2(n_442),
.B(n_406),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_380),
.A2(n_363),
.B1(n_340),
.B2(n_329),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_380),
.A2(n_329),
.B1(n_325),
.B2(n_310),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_424),
.A2(n_444),
.B1(n_448),
.B2(n_394),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_388),
.Y(n_425)
);

INVx13_ASAP7_75t_L g472 ( 
.A(n_425),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_388),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_427),
.B(n_441),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_398),
.B(n_350),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_434),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_327),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_406),
.A2(n_320),
.B(n_342),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_395),
.A2(n_313),
.B1(n_330),
.B2(n_354),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_386),
.Y(n_446)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_446),
.Y(n_461)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_447),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_395),
.A2(n_353),
.B1(n_359),
.B2(n_357),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_403),
.C(n_370),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_378),
.B(n_357),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_452),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_376),
.B(n_333),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_451),
.B(n_396),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_383),
.B(n_343),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_453),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_455),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_435),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_457),
.B(n_474),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_458),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_377),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_459),
.B(n_463),
.Y(n_500)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_418),
.B(n_367),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_460),
.B(n_481),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_452),
.B(n_401),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_430),
.B(n_404),
.Y(n_464)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_464),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_437),
.B(n_399),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_465),
.B(n_450),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_466),
.Y(n_495)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_428),
.Y(n_468)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_468),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_425),
.B(n_391),
.Y(n_469)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_469),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_440),
.B(n_333),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_470),
.B(n_475),
.Y(n_504)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_428),
.Y(n_471)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_471),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_476),
.C(n_478),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_445),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_371),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_437),
.B(n_406),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_403),
.C(n_379),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_445),
.B(n_387),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_479),
.A2(n_480),
.B(n_441),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_445),
.A2(n_408),
.B(n_395),
.Y(n_480)
);

AND2x6_ASAP7_75t_L g481 ( 
.A(n_417),
.B(n_382),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_486),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_427),
.B(n_368),
.Y(n_483)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_483),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_439),
.B(n_390),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_484),
.B(n_489),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_434),
.B(n_375),
.C(n_387),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_485),
.B(n_490),
.C(n_444),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g486 ( 
.A(n_417),
.B(n_411),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_421),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_431),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_488),
.A2(n_423),
.B1(n_416),
.B2(n_426),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_422),
.B(n_343),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_420),
.B(n_387),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_494),
.B(n_509),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_483),
.B(n_432),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_496),
.B(n_501),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_499),
.A2(n_503),
.B1(n_516),
.B2(n_526),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_456),
.B(n_432),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_490),
.A2(n_416),
.B1(n_426),
.B2(n_415),
.Y(n_503)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_507),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_456),
.B(n_464),
.Y(n_508)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_508),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_473),
.B(n_422),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_454),
.B(n_448),
.Y(n_512)
);

CKINVDCx14_ASAP7_75t_R g536 ( 
.A(n_512),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_514),
.A2(n_518),
.B(n_472),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_454),
.B(n_414),
.Y(n_515)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_515),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_479),
.A2(n_477),
.B1(n_466),
.B2(n_485),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_469),
.B(n_414),
.Y(n_517)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_517),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_480),
.A2(n_441),
.B(n_442),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_519),
.B(n_458),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_457),
.B(n_443),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_520),
.B(n_521),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_482),
.B(n_443),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_478),
.B(n_447),
.C(n_446),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_477),
.C(n_455),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_468),
.B(n_453),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_523),
.B(n_524),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_461),
.B(n_438),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_487),
.B(n_436),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_528),
.B(n_538),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_520),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_529),
.B(n_537),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_530),
.B(n_540),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_495),
.A2(n_477),
.B1(n_479),
.B2(n_481),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_531),
.A2(n_514),
.B1(n_496),
.B2(n_498),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_533),
.A2(n_547),
.B(n_526),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_509),
.B(n_465),
.C(n_476),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_534),
.B(n_545),
.C(n_555),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_407),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_522),
.B(n_472),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_504),
.B(n_438),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_500),
.B(n_314),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_541),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_500),
.B(n_316),
.Y(n_542)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_542),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_513),
.B(n_374),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_543),
.B(n_554),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_492),
.B(n_462),
.C(n_471),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_499),
.A2(n_486),
.B1(n_424),
.B2(n_394),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_546),
.A2(n_549),
.B1(n_551),
.B2(n_505),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_510),
.A2(n_467),
.B(n_462),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_525),
.A2(n_433),
.B1(n_384),
.B2(n_402),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_524),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_513),
.B(n_467),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_492),
.B(n_461),
.C(n_429),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_519),
.B(n_429),
.C(n_436),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_556),
.B(n_545),
.C(n_555),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_501),
.B(n_389),
.Y(n_557)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_557),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_507),
.Y(n_558)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_558),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_562),
.B(n_574),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_538),
.Y(n_563)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_563),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_556),
.B(n_516),
.C(n_497),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_564),
.B(n_567),
.Y(n_601)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_527),
.Y(n_565)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_565),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_550),
.B(n_511),
.C(n_494),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_536),
.A2(n_503),
.B1(n_525),
.B2(n_512),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_568),
.A2(n_582),
.B1(n_553),
.B2(n_552),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_535),
.Y(n_571)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_571),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_528),
.B(n_518),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_572),
.B(n_578),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_550),
.B(n_511),
.C(n_491),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_575),
.A2(n_460),
.B1(n_433),
.B2(n_502),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_576),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_546),
.A2(n_498),
.B1(n_505),
.B2(n_493),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_577),
.A2(n_549),
.B1(n_558),
.B2(n_527),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_530),
.B(n_491),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_534),
.B(n_515),
.C(n_517),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_580),
.B(n_583),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_533),
.B(n_521),
.C(n_493),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_532),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_584),
.B(n_585),
.Y(n_593)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_532),
.Y(n_585)
);

CKINVDCx16_ASAP7_75t_R g586 ( 
.A(n_569),
.Y(n_586)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_586),
.Y(n_610)
);

NAND3xp33_ASAP7_75t_L g587 ( 
.A(n_570),
.B(n_548),
.C(n_508),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_587),
.A2(n_574),
.B1(n_581),
.B2(n_561),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_562),
.B(n_531),
.C(n_547),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_SL g624 ( 
.A(n_589),
.B(n_597),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_590),
.A2(n_600),
.B1(n_564),
.B2(n_566),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_591),
.A2(n_596),
.B1(n_305),
.B2(n_319),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_580),
.B(n_548),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_592),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_568),
.A2(n_551),
.B1(n_553),
.B2(n_552),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_560),
.B(n_539),
.C(n_544),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_560),
.B(n_539),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_598),
.B(n_604),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_566),
.B(n_544),
.C(n_502),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_599),
.B(n_393),
.C(n_337),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_559),
.B(n_523),
.Y(n_603)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_603),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_578),
.B(n_506),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_600),
.A2(n_565),
.B1(n_579),
.B2(n_575),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_608),
.B(n_623),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_602),
.A2(n_576),
.B(n_583),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_612),
.A2(n_615),
.B(n_617),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_598),
.B(n_597),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_613),
.B(n_619),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_603),
.B(n_573),
.Y(n_614)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_614),
.Y(n_632)
);

CKINVDCx14_ASAP7_75t_R g616 ( 
.A(n_593),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_616),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_602),
.A2(n_577),
.B(n_572),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_618),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_596),
.A2(n_567),
.B(n_506),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_607),
.A2(n_402),
.B1(n_409),
.B2(n_392),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_620),
.B(n_622),
.Y(n_641)
);

XNOR2x1_ASAP7_75t_L g621 ( 
.A(n_604),
.B(n_385),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_621),
.B(n_591),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_589),
.B(n_337),
.C(n_305),
.Y(n_623)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_626),
.B(n_621),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_624),
.B(n_606),
.C(n_605),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_627),
.Y(n_650)
);

CKINVDCx16_ASAP7_75t_R g628 ( 
.A(n_619),
.Y(n_628)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_628),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_611),
.B(n_599),
.C(n_601),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_630),
.B(n_622),
.C(n_623),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_SL g634 ( 
.A1(n_626),
.A2(n_608),
.B(n_594),
.C(n_617),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_634),
.A2(n_625),
.B(n_614),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_609),
.B(n_588),
.Y(n_635)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_635),
.Y(n_651)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_638),
.B(n_639),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_611),
.B(n_595),
.Y(n_640)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_640),
.A2(n_316),
.B(n_358),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_SL g642 ( 
.A1(n_637),
.A2(n_612),
.B(n_618),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_642),
.A2(n_648),
.B(n_652),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_645),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_646),
.B(n_649),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_636),
.B(n_610),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_647),
.B(n_632),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_630),
.B(n_595),
.C(n_361),
.Y(n_648)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_627),
.B(n_352),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_631),
.A2(n_319),
.B(n_361),
.Y(n_652)
);

XOR2xp5_ASAP7_75t_L g658 ( 
.A(n_653),
.B(n_639),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_654),
.B(n_657),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_SL g657 ( 
.A1(n_650),
.A2(n_629),
.B1(n_633),
.B2(n_641),
.Y(n_657)
);

XOR2xp5_ASAP7_75t_L g666 ( 
.A(n_658),
.B(n_661),
.Y(n_666)
);

AOI322xp5_ASAP7_75t_L g659 ( 
.A1(n_643),
.A2(n_629),
.A3(n_634),
.B1(n_352),
.B2(n_361),
.C1(n_381),
.C2(n_366),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_SL g665 ( 
.A1(n_659),
.A2(n_352),
.B1(n_234),
.B2(n_308),
.Y(n_665)
);

XOR2xp5_ASAP7_75t_L g661 ( 
.A(n_646),
.B(n_634),
.Y(n_661)
);

AO21x1_ASAP7_75t_L g662 ( 
.A1(n_656),
.A2(n_651),
.B(n_649),
.Y(n_662)
);

AOI322xp5_ASAP7_75t_L g667 ( 
.A1(n_662),
.A2(n_661),
.A3(n_660),
.B1(n_658),
.B2(n_644),
.C1(n_366),
.C2(n_381),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_655),
.A2(n_634),
.B(n_648),
.Y(n_664)
);

XOR2xp5_ASAP7_75t_L g668 ( 
.A(n_664),
.B(n_665),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_667),
.A2(n_669),
.B(n_660),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_663),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g670 ( 
.A(n_668),
.B(n_663),
.C(n_666),
.Y(n_670)
);

OAI32xp33_ASAP7_75t_SL g672 ( 
.A1(n_670),
.A2(n_671),
.A3(n_644),
.B1(n_236),
.B2(n_318),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_672),
.A2(n_317),
.B(n_318),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_673),
.B(n_328),
.C(n_236),
.Y(n_674)
);

XOR2xp5_ASAP7_75t_L g675 ( 
.A(n_674),
.B(n_328),
.Y(n_675)
);


endmodule