module real_jpeg_6781_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_0),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_0),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_0),
.A2(n_208),
.B1(n_278),
.B2(n_281),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_0),
.A2(n_84),
.B1(n_86),
.B2(n_208),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_0),
.A2(n_143),
.B1(n_208),
.B2(n_422),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_1),
.A2(n_58),
.B1(n_154),
.B2(n_157),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_1),
.A2(n_58),
.B1(n_361),
.B2(n_363),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_1),
.A2(n_58),
.B1(n_383),
.B2(n_404),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_2),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_2),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_2),
.Y(n_245)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_2),
.Y(n_255)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_2),
.Y(n_266)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_3),
.Y(n_132)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_3),
.Y(n_146)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_3),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_3),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_3),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_4),
.A2(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_4),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_4),
.A2(n_88),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_4),
.A2(n_88),
.B1(n_299),
.B2(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_4),
.A2(n_88),
.B1(n_183),
.B2(n_307),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_5),
.A2(n_46),
.B1(n_48),
.B2(n_51),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_5),
.A2(n_51),
.B1(n_211),
.B2(n_333),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_5),
.A2(n_51),
.B1(n_403),
.B2(n_404),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_5),
.A2(n_51),
.B1(n_416),
.B2(n_419),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_6),
.A2(n_173),
.B1(n_176),
.B2(n_179),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_6),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_6),
.B(n_194),
.C(n_198),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_6),
.B(n_73),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_6),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_6),
.B(n_118),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_6),
.B(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_8),
.Y(n_518)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_9),
.Y(n_103)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_9),
.Y(n_110)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_9),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_10),
.A2(n_182),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_10),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_10),
.A2(n_186),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_10),
.A2(n_186),
.B1(n_290),
.B2(n_292),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_10),
.A2(n_186),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_12),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_12),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_12),
.A2(n_93),
.B1(n_105),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_12),
.A2(n_93),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_13),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_13),
.Y(n_115)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_13),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_14),
.A2(n_142),
.B1(n_143),
.B2(n_147),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_14),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_14),
.A2(n_142),
.B1(n_297),
.B2(n_299),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_14),
.A2(n_120),
.B1(n_142),
.B2(n_383),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_14),
.A2(n_142),
.B1(n_409),
.B2(n_412),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_15),
.A2(n_192),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_15),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_15),
.A2(n_231),
.B1(n_250),
.B2(n_252),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_15),
.A2(n_231),
.B1(n_305),
.B2(n_324),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_15),
.A2(n_55),
.B1(n_143),
.B2(n_231),
.Y(n_438)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_17),
.Y(n_520)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_516),
.B(n_519),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_162),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_160),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_133),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_23),
.B(n_133),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_122),
.B2(n_123),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_59),
.C(n_94),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_26),
.B(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_45),
.B1(n_52),
.B2(n_54),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_27),
.A2(n_52),
.B1(n_54),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_27),
.A2(n_45),
.B1(n_52),
.B2(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_27),
.A2(n_374),
.B(n_421),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_27),
.A2(n_36),
.B1(n_421),
.B2(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_28),
.A2(n_372),
.B(n_373),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_28),
.B(n_375),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_31),
.Y(n_350)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_33),
.Y(n_129)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_36),
.B(n_179),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_36)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_37),
.Y(n_352)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_40),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_40),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_40),
.Y(n_411)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_41),
.Y(n_326)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_43),
.Y(n_305)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_43),
.Y(n_414)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_52),
.A2(n_438),
.B(n_460),
.Y(n_470)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_53),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_53),
.B(n_141),
.Y(n_459)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_59),
.A2(n_94),
.B1(n_95),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_83),
.B1(n_89),
.B2(n_90),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_60),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_60),
.A2(n_83),
.B1(n_89),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_60),
.A2(n_89),
.B1(n_323),
.B2(n_380),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_60),
.A2(n_89),
.B1(n_408),
.B2(n_415),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_73),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_66),
.Y(n_287)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_72),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_73),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_73),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

AOI22x1_ASAP7_75t_L g439 ( 
.A1(n_73),
.A2(n_125),
.B1(n_328),
.B2(n_440),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_73),
.A2(n_125),
.B1(n_153),
.B2(n_448),
.Y(n_447)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_79),
.B2(n_82),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_75),
.Y(n_309)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_77),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_78),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_78),
.Y(n_192)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_79),
.Y(n_404)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_81),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_81),
.Y(n_234)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_81),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_81),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_81),
.Y(n_383)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_SL g284 ( 
.A1(n_86),
.A2(n_179),
.B(n_285),
.Y(n_284)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_89),
.B(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_89),
.A2(n_323),
.B(n_327),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_94),
.B(n_139),
.C(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_94),
.A2(n_95),
.B1(n_150),
.B2(n_151),
.Y(n_505)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_117),
.B(n_119),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_96),
.A2(n_172),
.B(n_180),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_96),
.A2(n_117),
.B1(n_230),
.B2(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_96),
.A2(n_180),
.B(n_277),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_96),
.A2(n_117),
.B1(n_382),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_97),
.B(n_181),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_97),
.A2(n_118),
.B1(n_402),
.B2(n_405),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_97),
.A2(n_118),
.B1(n_405),
.B2(n_426),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_97),
.A2(n_118),
.B1(n_426),
.B2(n_451),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_98)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_99),
.Y(n_403)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_102),
.Y(n_281)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_103),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_107),
.A2(n_230),
.B(n_235),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_114),
.B2(n_116),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_113),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g298 ( 
.A(n_113),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_113),
.Y(n_299)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_114),
.Y(n_243)
);

BUFx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g365 ( 
.A(n_115),
.Y(n_365)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_115),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_117),
.A2(n_235),
.B(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_118),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_119),
.Y(n_451)
);

INVx5_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_125),
.A2(n_284),
.B(n_288),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_125),
.B(n_328),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_125),
.A2(n_288),
.B(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.C(n_148),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_511)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_138),
.A2(n_139),
.B1(n_505),
.B2(n_506),
.Y(n_504)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_148),
.A2(n_149),
.B1(n_510),
.B2(n_511),
.Y(n_509)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g344 ( 
.A1(n_154),
.A2(n_345),
.A3(n_350),
.B1(n_351),
.B2(n_353),
.Y(n_344)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_499),
.B(n_513),
.Y(n_163)
);

OAI311xp33_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_386),
.A3(n_475),
.B1(n_493),
.C1(n_494),
.Y(n_164)
);

AOI21x1_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_338),
.B(n_385),
.Y(n_165)
);

AO21x1_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_314),
.B(n_337),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_271),
.B(n_313),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_238),
.B(n_270),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_203),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_170),
.B(n_203),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_189),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_171),
.A2(n_189),
.B1(n_190),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_171),
.Y(n_268)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_179),
.A2(n_213),
.B(n_221),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_179),
.B(n_354),
.Y(n_353)
);

OAI21xp33_ASAP7_75t_SL g372 ( 
.A1(n_179),
.A2(n_346),
.B(n_353),
.Y(n_372)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_201),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_227),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_204),
.B(n_228),
.C(n_237),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_213),
.B(n_221),
.Y(n_204)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_205),
.Y(n_262)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_213),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_213),
.A2(n_392),
.B1(n_395),
.B2(n_397),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_213),
.A2(n_254),
.B(n_397),
.Y(n_427)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_224),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_214),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_214),
.A2(n_296),
.B1(n_332),
.B2(n_335),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_214),
.A2(n_360),
.B1(n_434),
.B2(n_435),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_222),
.Y(n_358)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_225),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_236),
.B2(n_237),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_259),
.B(n_269),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_247),
.B(n_258),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_246),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_245),
.Y(n_396)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_245),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_257),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_257),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_254),
.B(n_256),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_250),
.Y(n_334)
);

INVx8_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_251),
.Y(n_400)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_254),
.Y(n_335)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_256),
.A2(n_295),
.B(n_300),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_267),
.Y(n_269)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_273),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_293),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_282),
.B2(n_283),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_282),
.C(n_293),
.Y(n_315)
);

INVx3_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI32xp33_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_304),
.A3(n_306),
.B1(n_308),
.B2(n_310),
.Y(n_303)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_290),
.B(n_352),
.Y(n_351)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_303),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_303),
.Y(n_320)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_311),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_315),
.B(n_316),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_321),
.B2(n_336),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_320),
.C(n_336),
.Y(n_339)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_321),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_329),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_330),
.C(n_331),
.Y(n_366)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_326),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_326),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_332),
.Y(n_357)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_339),
.B(n_340),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_369),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.Y(n_341)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_342),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_355),
.B2(n_356),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_344),
.B(n_355),
.Y(n_471)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_349),
.Y(n_354)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_354),
.Y(n_422)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx6_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_366),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_366),
.B(n_367),
.C(n_369),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_371),
.B1(n_378),
.B2(n_384),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_370),
.B(n_379),
.C(n_381),
.Y(n_484)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_378),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_381),
.Y(n_378)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_380),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_461),
.Y(n_386)
);

A2O1A1Ixp33_ASAP7_75t_SL g494 ( 
.A1(n_387),
.A2(n_461),
.B(n_495),
.C(n_498),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_441),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_388),
.B(n_441),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_423),
.C(n_429),
.Y(n_388)
);

FAx1_ASAP7_75t_SL g474 ( 
.A(n_389),
.B(n_423),
.CI(n_429),
.CON(n_474),
.SN(n_474)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_406),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_390),
.B(n_407),
.C(n_420),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_401),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_391),
.B(n_401),
.Y(n_467)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_392),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_420),
.Y(n_406)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_408),
.Y(n_440)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_415),
.Y(n_448)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_424),
.A2(n_425),
.B1(n_427),
.B2(n_428),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_427),
.Y(n_455)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_427),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_427),
.A2(n_428),
.B1(n_457),
.B2(n_458),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_427),
.A2(n_455),
.B(n_458),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_436),
.C(n_439),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_430),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_433),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_431),
.B(n_433),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_436),
.A2(n_437),
.B1(n_439),
.B2(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_439),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_442),
.B(n_445),
.C(n_453),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_445),
.B1(n_453),
.B2(n_454),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_449),
.B(n_452),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_447),
.B(n_450),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_452),
.B(n_504),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_452),
.B(n_502),
.C(n_504),
.Y(n_512)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_474),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_462),
.B(n_474),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_467),
.C(n_468),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_463),
.A2(n_464),
.B1(n_467),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_468),
.B(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_471),
.C(n_472),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_469),
.A2(n_470),
.B1(n_472),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_472),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g522 ( 
.A(n_474),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_488),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_477),
.A2(n_496),
.B(n_497),
.Y(n_495)
);

NOR2x1_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_485),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_485),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_482),
.C(n_484),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_491),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_482),
.A2(n_483),
.B1(n_484),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_484),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_490),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_508),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_507),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_501),
.B(n_507),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_505),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_508),
.A2(n_514),
.B(n_515),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_509),
.B(n_512),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_509),
.B(n_512),
.Y(n_515)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

BUFx4f_ASAP7_75t_SL g516 ( 
.A(n_517),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_517),
.B(n_520),
.Y(n_519)
);

INVx13_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);


endmodule