module fake_jpeg_23162_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_41),
.Y(n_55)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_26),
.B1(n_22),
.B2(n_30),
.Y(n_52)
);

INVx2_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_21),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_38),
.B1(n_26),
.B2(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_56),
.B1(n_54),
.B2(n_60),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_40),
.B(n_18),
.C(n_29),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_46),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_68),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_15),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_78),
.Y(n_92)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_88),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_84),
.B(n_98),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_38),
.B1(n_58),
.B2(n_49),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_97),
.B1(n_78),
.B2(n_74),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_51),
.B(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_89),
.Y(n_109)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_61),
.B1(n_44),
.B2(n_20),
.Y(n_111)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_68),
.B(n_48),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_37),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_73),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_64),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_65),
.A2(n_44),
.B1(n_60),
.B2(n_20),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_0),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_43),
.B1(n_67),
.B2(n_29),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_71),
.B1(n_69),
.B2(n_73),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_111),
.B1(n_113),
.B2(n_117),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_71),
.C(n_73),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_108),
.C(n_110),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_116),
.B(n_28),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_62),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_66),
.C(n_64),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_24),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_82),
.A2(n_84),
.B1(n_79),
.B2(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_24),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_1),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_67),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_97),
.B1(n_96),
.B2(n_98),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_87),
.B(n_98),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_122),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_43),
.B1(n_16),
.B2(n_28),
.Y(n_123)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_16),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_37),
.C(n_80),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_131),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_43),
.C(n_28),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_134),
.A2(n_113),
.B1(n_102),
.B2(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_19),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_135),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_134),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_SL g138 ( 
.A1(n_130),
.A2(n_116),
.A3(n_107),
.B1(n_102),
.B2(n_117),
.C1(n_99),
.C2(n_14),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_138),
.A2(n_132),
.B(n_128),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_107),
.B1(n_116),
.B2(n_29),
.Y(n_140)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_19),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_19),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_125),
.C(n_126),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_154),
.C(n_161),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_146),
.B1(n_145),
.B2(n_150),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_125),
.C(n_119),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_155),
.A2(n_159),
.B(n_136),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_121),
.B(n_120),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_157),
.B(n_142),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_135),
.B(n_118),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_121),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_163),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_162),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_127),
.C(n_23),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_23),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_165),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_143),
.C(n_139),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_169),
.C(n_173),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_142),
.C(n_149),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_172),
.B(n_153),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_136),
.B(n_3),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_174),
.A2(n_2),
.B(n_3),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_158),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_168),
.C(n_167),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_178),
.B(n_167),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g179 ( 
.A1(n_171),
.A2(n_2),
.B(n_3),
.C(n_5),
.Y(n_179)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_178),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_181),
.Y(n_183)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_166),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_188),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_189),
.B(n_179),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_5),
.C(n_6),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_193),
.Y(n_196)
);

NOR2xp67_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_182),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_6),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_7),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_195),
.A2(n_190),
.B(n_9),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_186),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_8),
.C(n_10),
.Y(n_199)
);

AOI21x1_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_199),
.B(n_10),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_196),
.Y(n_201)
);


endmodule