module fake_aes_8679_n_708 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_708);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_708;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g78 ( .A(n_19), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_36), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_7), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_10), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_39), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_46), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_43), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_47), .Y(n_85) );
BUFx3_ASAP7_75t_L g86 ( .A(n_29), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_2), .Y(n_87) );
INVxp33_ASAP7_75t_L g88 ( .A(n_33), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_13), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_30), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_28), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_68), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_64), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_72), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_11), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_2), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_61), .Y(n_97) );
BUFx2_ASAP7_75t_L g98 ( .A(n_6), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_42), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_17), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_70), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_21), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_37), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_74), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_9), .Y(n_105) );
INVxp33_ASAP7_75t_L g106 ( .A(n_44), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_21), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_75), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_71), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_32), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_54), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_50), .Y(n_112) );
INVxp33_ASAP7_75t_SL g113 ( .A(n_15), .Y(n_113) );
CKINVDCx14_ASAP7_75t_R g114 ( .A(n_38), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_12), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_11), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_8), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_59), .B(n_18), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_73), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_10), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_1), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_76), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_65), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_34), .Y(n_124) );
INVxp33_ASAP7_75t_SL g125 ( .A(n_66), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_58), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_80), .B(n_0), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_98), .B(n_0), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_84), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_93), .Y(n_136) );
NOR2xp67_ASAP7_75t_L g137 ( .A(n_85), .B(n_1), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_85), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_90), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_80), .B(n_3), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_90), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_112), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_91), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_115), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_92), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_86), .B(n_27), .Y(n_147) );
AND3x1_ASAP7_75t_L g148 ( .A(n_81), .B(n_3), .C(n_4), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_86), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_116), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_120), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_92), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_97), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_88), .B(n_4), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_97), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_81), .B(n_5), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_108), .Y(n_157) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_87), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_87), .B(n_5), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_108), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_109), .Y(n_161) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_109), .A2(n_35), .B(n_77), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_119), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_119), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_123), .Y(n_165) );
OR2x2_ASAP7_75t_L g166 ( .A(n_89), .B(n_6), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_114), .Y(n_167) );
NOR2xp33_ASAP7_75t_SL g168 ( .A(n_82), .B(n_40), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_123), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_89), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_128), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_128), .Y(n_172) );
OR2x2_ASAP7_75t_L g173 ( .A(n_131), .B(n_78), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_158), .B(n_96), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_149), .Y(n_175) );
AO22x2_ASAP7_75t_L g176 ( .A1(n_128), .A2(n_121), .B1(n_95), .B2(n_102), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_167), .B(n_106), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_128), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_167), .B(n_126), .Y(n_180) );
OAI21xp33_ASAP7_75t_L g181 ( .A1(n_127), .A2(n_100), .B(n_95), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_131), .B(n_121), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_128), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_158), .B(n_96), .Y(n_184) );
OR2x2_ASAP7_75t_L g185 ( .A(n_144), .B(n_107), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_144), .B(n_100), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_152), .Y(n_187) );
BUFx2_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_152), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_136), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_170), .A2(n_151), .B1(n_154), .B2(n_132), .Y(n_191) );
INVx5_ASAP7_75t_L g192 ( .A(n_147), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_127), .B(n_103), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_134), .B(n_102), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_142), .Y(n_196) );
OA22x2_ASAP7_75t_L g197 ( .A1(n_132), .A2(n_117), .B1(n_105), .B2(n_124), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_152), .B(n_124), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_154), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_160), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_160), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_134), .B(n_117), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g203 ( .A(n_168), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_135), .B(n_110), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_135), .B(n_99), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_149), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_149), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_160), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_149), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_130), .B(n_104), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_149), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_149), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_130), .B(n_125), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_139), .B(n_113), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_160), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_139), .B(n_122), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_161), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_161), .Y(n_218) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_166), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_147), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_145), .B(n_169), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_169), .B(n_111), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_161), .Y(n_223) );
AND2x6_ASAP7_75t_L g224 ( .A(n_161), .B(n_118), .Y(n_224) );
NAND3xp33_ASAP7_75t_L g225 ( .A(n_145), .B(n_101), .C(n_94), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_153), .B(n_7), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_130), .B(n_41), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_153), .B(n_8), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_165), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_157), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_155), .B(n_164), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_157), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_219), .Y(n_234) );
OR2x6_ASAP7_75t_L g235 ( .A(n_188), .B(n_166), .Y(n_235) );
CKINVDCx6p67_ASAP7_75t_R g236 ( .A(n_190), .Y(n_236) );
INVx5_ASAP7_75t_L g237 ( .A(n_198), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_184), .B(n_166), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_219), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_222), .B(n_130), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_222), .B(n_130), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_222), .B(n_165), .Y(n_242) );
AND3x2_ASAP7_75t_SL g243 ( .A(n_203), .B(n_148), .C(n_163), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_184), .B(n_140), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_207), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_227), .Y(n_246) );
NOR2xp33_ASAP7_75t_R g247 ( .A(n_190), .B(n_168), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_221), .B(n_165), .Y(n_248) );
OR2x6_ASAP7_75t_SL g249 ( .A(n_196), .B(n_140), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_227), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_207), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_220), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_196), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_212), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_191), .Y(n_255) );
AND3x1_ASAP7_75t_L g256 ( .A(n_186), .B(n_159), .C(n_156), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_224), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_174), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_176), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_176), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_176), .Y(n_261) );
INVx2_ASAP7_75t_SL g262 ( .A(n_174), .Y(n_262) );
BUFx12f_ASAP7_75t_L g263 ( .A(n_174), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_224), .Y(n_264) );
INVxp67_ASAP7_75t_L g265 ( .A(n_232), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_220), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_182), .B(n_148), .Y(n_267) );
BUFx10_ASAP7_75t_L g268 ( .A(n_180), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_195), .B(n_164), .Y(n_269) );
OR2x6_ASAP7_75t_L g270 ( .A(n_197), .B(n_173), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_195), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_195), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_202), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_220), .B(n_157), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_202), .B(n_155), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_185), .B(n_156), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_202), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_177), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_212), .Y(n_279) );
NAND2xp33_ASAP7_75t_SL g280 ( .A(n_214), .B(n_159), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_220), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_199), .Y(n_282) );
OR2x6_ASAP7_75t_L g283 ( .A(n_197), .B(n_137), .Y(n_283) );
BUFx8_ASAP7_75t_L g284 ( .A(n_224), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_180), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_171), .B(n_143), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_213), .B(n_137), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_172), .B(n_179), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_187), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_198), .Y(n_290) );
OR2x6_ASAP7_75t_L g291 ( .A(n_183), .B(n_163), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_189), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_198), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_192), .Y(n_294) );
INVx3_ASAP7_75t_SL g295 ( .A(n_198), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_216), .Y(n_296) );
INVx2_ASAP7_75t_SL g297 ( .A(n_213), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_198), .B(n_163), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_193), .B(n_143), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_200), .Y(n_300) );
BUFx12f_ASAP7_75t_L g301 ( .A(n_224), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_295), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_263), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_265), .B(n_225), .Y(n_304) );
OAI22xp33_ASAP7_75t_L g305 ( .A1(n_235), .A2(n_229), .B1(n_204), .B2(n_205), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_265), .Y(n_306) );
BUFx10_ASAP7_75t_L g307 ( .A(n_238), .Y(n_307) );
CKINVDCx8_ASAP7_75t_R g308 ( .A(n_253), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_244), .B(n_194), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_271), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_278), .B(n_194), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_295), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_290), .Y(n_313) );
INVx3_ASAP7_75t_SL g314 ( .A(n_258), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_296), .B(n_224), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_288), .A2(n_269), .B(n_275), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_288), .A2(n_210), .B(n_192), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_260), .Y(n_318) );
INVx5_ASAP7_75t_L g319 ( .A(n_237), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_278), .B(n_217), .Y(n_320) );
INVx3_ASAP7_75t_SL g321 ( .A(n_235), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_272), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_234), .A2(n_181), .B1(n_133), .B2(n_138), .C(n_129), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_238), .B(n_208), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_273), .Y(n_325) );
BUFx12f_ASAP7_75t_L g326 ( .A(n_235), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_290), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_262), .B(n_210), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_301), .B(n_129), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_292), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_237), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_269), .A2(n_192), .B(n_218), .Y(n_332) );
BUFx12f_ASAP7_75t_L g333 ( .A(n_282), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_289), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_291), .Y(n_335) );
OAI22xp33_ASAP7_75t_L g336 ( .A1(n_276), .A2(n_129), .B1(n_133), .B2(n_146), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_300), .Y(n_337) );
NAND2x1p5_ASAP7_75t_L g338 ( .A(n_237), .B(n_192), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_245), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_281), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_251), .Y(n_341) );
BUFx12f_ASAP7_75t_L g342 ( .A(n_267), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_291), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_291), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_239), .B(n_226), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_275), .B(n_230), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_277), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_248), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_256), .B(n_297), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_L g350 ( .A1(n_270), .A2(n_201), .B(n_215), .C(n_223), .Y(n_350) );
CKINVDCx16_ASAP7_75t_R g351 ( .A(n_247), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_246), .B(n_133), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_236), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_248), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_334), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_316), .A2(n_261), .B1(n_259), .B2(n_250), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_348), .B(n_270), .Y(n_357) );
BUFx12f_ASAP7_75t_L g358 ( .A(n_326), .Y(n_358) );
INVxp33_ASAP7_75t_L g359 ( .A(n_349), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_340), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_306), .A2(n_255), .B1(n_267), .B2(n_285), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_334), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_354), .B(n_270), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_321), .B(n_240), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_349), .A2(n_280), .B1(n_283), .B2(n_268), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_337), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_340), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_309), .B(n_268), .Y(n_368) );
NAND3x1_ASAP7_75t_L g369 ( .A(n_321), .B(n_243), .C(n_249), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_326), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_340), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_340), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_335), .B(n_257), .Y(n_373) );
CKINVDCx11_ASAP7_75t_R g374 ( .A(n_308), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_311), .A2(n_283), .B1(n_287), .B2(n_284), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_336), .A2(n_283), .B1(n_286), .B2(n_143), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_337), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_340), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_309), .B(n_304), .Y(n_379) );
NAND3xp33_ASAP7_75t_SL g380 ( .A(n_308), .B(n_247), .C(n_353), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_317), .A2(n_286), .B(n_242), .Y(n_381) );
OR2x2_ASAP7_75t_SL g382 ( .A(n_351), .B(n_243), .Y(n_382) );
OAI211xp5_ASAP7_75t_L g383 ( .A1(n_350), .A2(n_242), .B(n_240), .C(n_241), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_324), .B(n_241), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_349), .A2(n_287), .B1(n_299), .B2(n_138), .C(n_141), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g386 ( .A1(n_305), .A2(n_298), .B(n_299), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_318), .A2(n_284), .B1(n_264), .B2(n_293), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_304), .B(n_293), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_376), .A2(n_335), .B1(n_343), .B2(n_344), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_355), .Y(n_390) );
OAI211xp5_ASAP7_75t_L g391 ( .A1(n_375), .A2(n_323), .B(n_353), .C(n_303), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g393 ( .A1(n_375), .A2(n_303), .B(n_320), .C(n_352), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_368), .A2(n_304), .B1(n_324), .B2(n_322), .C(n_325), .Y(n_394) );
OAI211xp5_ASAP7_75t_L g395 ( .A1(n_365), .A2(n_318), .B(n_345), .C(n_344), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_368), .B(n_343), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_379), .A2(n_342), .B1(n_333), .B2(n_329), .Y(n_397) );
AO21x2_ASAP7_75t_L g398 ( .A1(n_356), .A2(n_315), .B(n_228), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_381), .A2(n_332), .B(n_330), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_384), .B(n_310), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_379), .A2(n_342), .B1(n_333), .B2(n_329), .Y(n_401) );
OAI21x1_ASAP7_75t_L g402 ( .A1(n_360), .A2(n_331), .B(n_162), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_362), .Y(n_403) );
NAND3xp33_ASAP7_75t_L g404 ( .A(n_386), .B(n_157), .C(n_228), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_362), .Y(n_405) );
OAI21x1_ASAP7_75t_L g406 ( .A1(n_360), .A2(n_331), .B(n_162), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g407 ( .A1(n_376), .A2(n_307), .B1(n_329), .B2(n_312), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_366), .Y(n_408) );
OR2x6_ASAP7_75t_L g409 ( .A(n_366), .B(n_329), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_358), .A2(n_307), .B1(n_312), .B2(n_302), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_357), .A2(n_314), .B1(n_307), .B2(n_328), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_357), .A2(n_314), .B1(n_328), .B2(n_347), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_377), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_384), .B(n_346), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_377), .Y(n_415) );
AOI211xp5_ASAP7_75t_L g416 ( .A1(n_359), .A2(n_328), .B(n_141), .C(n_138), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_356), .Y(n_417) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_405), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_405), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_394), .A2(n_369), .B1(n_386), .B2(n_363), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_409), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_405), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_415), .B(n_363), .Y(n_423) );
NOR2x1_ASAP7_75t_L g424 ( .A(n_409), .B(n_380), .Y(n_424) );
OAI31xp33_ASAP7_75t_L g425 ( .A1(n_393), .A2(n_383), .A3(n_361), .B(n_364), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_415), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_415), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_390), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_390), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
OAI321xp33_ASAP7_75t_L g431 ( .A1(n_389), .A2(n_385), .A3(n_387), .B1(n_388), .B2(n_369), .C(n_364), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_392), .B(n_330), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_403), .Y(n_433) );
AOI33xp33_ASAP7_75t_L g434 ( .A1(n_397), .A2(n_141), .A3(n_146), .B1(n_382), .B2(n_233), .B3(n_231), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_403), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_408), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_408), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_413), .B(n_360), .Y(n_438) );
INVx5_ASAP7_75t_L g439 ( .A(n_409), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_413), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_389), .A2(n_388), .B1(n_373), .B2(n_146), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_417), .B(n_367), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_417), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_402), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_396), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g446 ( .A(n_401), .B(n_382), .C(n_373), .D(n_298), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_414), .B(n_373), .Y(n_447) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_404), .A2(n_378), .B(n_367), .Y(n_448) );
NOR2xp33_ASAP7_75t_R g449 ( .A(n_414), .B(n_374), .Y(n_449) );
OAI221xp5_ASAP7_75t_SL g450 ( .A1(n_395), .A2(n_370), .B1(n_358), .B2(n_341), .C(n_339), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_400), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_404), .B(n_373), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_409), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_428), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_428), .Y(n_455) );
NAND4xp25_ASAP7_75t_L g456 ( .A(n_425), .B(n_412), .C(n_391), .D(n_416), .Y(n_456) );
OAI33xp33_ASAP7_75t_L g457 ( .A1(n_446), .A2(n_9), .A3(n_12), .B1(n_13), .B2(n_14), .B3(n_15), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_430), .Y(n_458) );
AND4x1_ASAP7_75t_L g459 ( .A(n_425), .B(n_358), .C(n_416), .D(n_411), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_430), .Y(n_460) );
AOI33xp33_ASAP7_75t_L g461 ( .A1(n_451), .A2(n_407), .A3(n_396), .B1(n_410), .B2(n_18), .B3(n_19), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_439), .B(n_372), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_436), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g464 ( .A1(n_446), .A2(n_409), .B1(n_399), .B2(n_157), .C(n_162), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_451), .B(n_157), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_432), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_426), .B(n_398), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_436), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_453), .B(n_398), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_426), .B(n_398), .Y(n_470) );
OAI221xp5_ASAP7_75t_L g471 ( .A1(n_420), .A2(n_157), .B1(n_162), .B2(n_339), .C(n_341), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_418), .B(n_14), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_427), .B(n_162), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_445), .B(n_16), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_432), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_419), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_437), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_418), .B(n_16), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_422), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_449), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_437), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_440), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_422), .A2(n_372), .B(n_378), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_419), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_420), .A2(n_378), .B1(n_367), .B2(n_371), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_429), .B(n_17), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_440), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_429), .B(n_20), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_445), .B(n_20), .Y(n_489) );
INVx3_ASAP7_75t_L g490 ( .A(n_422), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_419), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_441), .A2(n_147), .B1(n_313), .B2(n_327), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_429), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_427), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_450), .B(n_175), .C(n_178), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_433), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_439), .B(n_302), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_433), .B(n_406), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_433), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_431), .A2(n_402), .B(n_406), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_435), .Y(n_501) );
OAI22xp5_ASAP7_75t_SL g502 ( .A1(n_441), .A2(n_302), .B1(n_312), .B2(n_371), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_435), .Y(n_503) );
NOR2xp33_ASAP7_75t_R g504 ( .A(n_480), .B(n_439), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_494), .Y(n_505) );
NOR2xp33_ASAP7_75t_R g506 ( .A(n_479), .B(n_439), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_479), .Y(n_507) );
INVxp33_ASAP7_75t_L g508 ( .A(n_502), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_457), .B(n_431), .C(n_450), .Y(n_509) );
BUFx2_ASAP7_75t_L g510 ( .A(n_490), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_496), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_493), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_466), .B(n_423), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_496), .Y(n_514) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_472), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_454), .Y(n_516) );
NAND2xp33_ASAP7_75t_R g517 ( .A(n_490), .B(n_472), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_467), .B(n_443), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_467), .B(n_443), .Y(n_519) );
INVx2_ASAP7_75t_SL g520 ( .A(n_490), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_459), .B(n_447), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_475), .B(n_423), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_499), .B(n_501), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_499), .B(n_435), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_476), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_470), .B(n_442), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_455), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_476), .Y(n_528) );
OAI221xp5_ASAP7_75t_SL g529 ( .A1(n_461), .A2(n_434), .B1(n_447), .B2(n_452), .C(n_421), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_470), .B(n_442), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_484), .Y(n_531) );
BUFx2_ASAP7_75t_L g532 ( .A(n_484), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_458), .B(n_423), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_460), .B(n_438), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_503), .B(n_452), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_491), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_491), .B(n_442), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_463), .B(n_448), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_468), .B(n_438), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_477), .B(n_438), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_481), .B(n_432), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_482), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_456), .A2(n_421), .B1(n_453), .B2(n_439), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_498), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_487), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_498), .B(n_448), .Y(n_546) );
OAI21xp33_ASAP7_75t_L g547 ( .A1(n_461), .A2(n_424), .B(n_453), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_478), .B(n_453), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_478), .B(n_448), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_474), .B(n_424), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_469), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_469), .B(n_448), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_489), .B(n_439), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_486), .B(n_439), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_464), .A2(n_444), .B(n_371), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_486), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_469), .B(n_444), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_488), .B(n_444), .Y(n_558) );
NOR2x1_ASAP7_75t_L g559 ( .A(n_488), .B(n_372), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_465), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_485), .B(n_462), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_473), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_526), .B(n_485), .Y(n_563) );
NOR4xp25_ASAP7_75t_SL g564 ( .A(n_517), .B(n_471), .C(n_462), .D(n_500), .Y(n_564) );
OAI21xp33_ASAP7_75t_SL g565 ( .A1(n_508), .A2(n_492), .B(n_473), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_526), .B(n_497), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_505), .B(n_483), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_530), .B(n_497), .Y(n_568) );
AOI21xp33_ASAP7_75t_L g569 ( .A1(n_508), .A2(n_495), .B(n_175), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_515), .B(n_518), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_542), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_532), .Y(n_572) );
OR2x6_ASAP7_75t_L g573 ( .A(n_507), .B(n_372), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_544), .B(n_211), .Y(n_574) );
A2O1A1O1Ixp25_ASAP7_75t_L g575 ( .A1(n_547), .A2(n_22), .B(n_23), .C(n_24), .D(n_25), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_509), .A2(n_147), .B1(n_175), .B2(n_372), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_518), .B(n_175), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_519), .B(n_206), .Y(n_578) );
AOI31xp33_ASAP7_75t_L g579 ( .A1(n_543), .A2(n_338), .A3(n_31), .B(n_45), .Y(n_579) );
AOI22xp5_ASAP7_75t_SL g580 ( .A1(n_521), .A2(n_372), .B1(n_312), .B2(n_302), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_532), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_542), .Y(n_582) );
AOI322xp5_ASAP7_75t_L g583 ( .A1(n_556), .A2(n_209), .A3(n_206), .B1(n_211), .B2(n_178), .C1(n_233), .C2(n_231), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_555), .A2(n_302), .B(n_312), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_530), .B(n_26), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_550), .A2(n_147), .B1(n_209), .B2(n_327), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_516), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_527), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_545), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_533), .B(n_48), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_512), .Y(n_591) );
AND2x4_ASAP7_75t_SL g592 ( .A(n_537), .B(n_331), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_531), .Y(n_593) );
OAI21xp33_ASAP7_75t_L g594 ( .A1(n_552), .A2(n_274), .B(n_279), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_519), .B(n_147), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_512), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_523), .Y(n_597) );
NAND3xp33_ASAP7_75t_L g598 ( .A(n_529), .B(n_274), .C(n_319), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_513), .B(n_49), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_553), .A2(n_147), .B1(n_313), .B2(n_327), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_522), .B(n_51), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_523), .Y(n_602) );
AOI211xp5_ASAP7_75t_SL g603 ( .A1(n_504), .A2(n_52), .B(n_53), .C(n_55), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_535), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_561), .B(n_319), .C(n_254), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_554), .A2(n_147), .B1(n_313), .B2(n_319), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_535), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_544), .B(n_56), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_524), .B(n_57), .Y(n_609) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_561), .A2(n_60), .B(n_62), .Y(n_610) );
INVx2_ASAP7_75t_SL g611 ( .A(n_506), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_524), .Y(n_612) );
INVx3_ASAP7_75t_SL g613 ( .A(n_520), .Y(n_613) );
NOR3xp33_ASAP7_75t_SL g614 ( .A(n_560), .B(n_63), .C(n_67), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_534), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_613), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_587), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_604), .B(n_546), .Y(n_618) );
AOI33xp33_ASAP7_75t_L g619 ( .A1(n_615), .A2(n_552), .A3(n_546), .B1(n_562), .B2(n_557), .B3(n_538), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_611), .B(n_510), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_570), .B(n_531), .Y(n_621) );
CKINVDCx16_ASAP7_75t_R g622 ( .A(n_566), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_588), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_589), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_579), .A2(n_559), .B(n_520), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_607), .B(n_549), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_571), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_565), .A2(n_548), .B1(n_551), .B2(n_549), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_582), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_597), .B(n_602), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_591), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_596), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_612), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_568), .B(n_557), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_567), .Y(n_635) );
INVx3_ASAP7_75t_L g636 ( .A(n_573), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_572), .Y(n_637) );
OAI21xp5_ASAP7_75t_L g638 ( .A1(n_575), .A2(n_538), .B(n_541), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_563), .B(n_551), .Y(n_639) );
XNOR2x2_ASAP7_75t_L g640 ( .A(n_605), .B(n_548), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_593), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_581), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_578), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_574), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g645 ( .A1(n_579), .A2(n_540), .B(n_539), .Y(n_645) );
XNOR2x2_ASAP7_75t_L g646 ( .A(n_585), .B(n_558), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_590), .A2(n_537), .B1(n_511), .B2(n_514), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_577), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_599), .A2(n_511), .B1(n_514), .B2(n_525), .Y(n_649) );
INVx3_ASAP7_75t_L g650 ( .A(n_573), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_573), .Y(n_651) );
INVxp67_ASAP7_75t_SL g652 ( .A(n_580), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_635), .B(n_525), .Y(n_653) );
NOR3xp33_ASAP7_75t_L g654 ( .A(n_652), .B(n_610), .C(n_569), .Y(n_654) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_637), .Y(n_655) );
INVxp67_ASAP7_75t_L g656 ( .A(n_616), .Y(n_656) );
AOI322xp5_ASAP7_75t_L g657 ( .A1(n_622), .A2(n_569), .A3(n_610), .B1(n_601), .B2(n_614), .C1(n_576), .C2(n_595), .Y(n_657) );
AOI221x1_ASAP7_75t_L g658 ( .A1(n_642), .A2(n_594), .B1(n_608), .B2(n_584), .C(n_598), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_619), .B(n_633), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_617), .Y(n_660) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_652), .A2(n_603), .B(n_592), .C(n_609), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_641), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_625), .A2(n_603), .B(n_583), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_623), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_628), .A2(n_595), .B1(n_528), .B2(n_536), .C(n_600), .Y(n_665) );
O2A1O1Ixp33_ASAP7_75t_L g666 ( .A1(n_620), .A2(n_564), .B(n_536), .C(n_528), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_651), .B(n_606), .Y(n_667) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_621), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_628), .B(n_564), .C(n_586), .Y(n_669) );
XOR2xp5_ASAP7_75t_L g670 ( .A(n_646), .B(n_69), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_624), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_641), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_618), .B(n_338), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_620), .A2(n_281), .B(n_266), .Y(n_674) );
CKINVDCx16_ASAP7_75t_R g675 ( .A(n_670), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_659), .B(n_619), .Y(n_676) );
INVx3_ASAP7_75t_L g677 ( .A(n_662), .Y(n_677) );
O2A1O1Ixp33_ASAP7_75t_L g678 ( .A1(n_666), .A2(n_645), .B(n_638), .C(n_651), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_655), .Y(n_679) );
OAI32xp33_ASAP7_75t_L g680 ( .A1(n_659), .A2(n_650), .A3(n_636), .B1(n_630), .B2(n_626), .Y(n_680) );
OAI311xp33_ASAP7_75t_L g681 ( .A1(n_663), .A2(n_647), .A3(n_650), .B1(n_636), .C1(n_649), .Y(n_681) );
AOI21xp33_ASAP7_75t_SL g682 ( .A1(n_661), .A2(n_663), .B(n_669), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_653), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_674), .A2(n_650), .B(n_636), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_656), .A2(n_648), .B1(n_639), .B2(n_643), .Y(n_685) );
AOI321xp33_ASAP7_75t_L g686 ( .A1(n_654), .A2(n_644), .A3(n_629), .B1(n_631), .B2(n_627), .C(n_632), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_653), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_660), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_667), .A2(n_634), .B1(n_644), .B2(n_640), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_657), .A2(n_252), .B(n_266), .C(n_281), .Y(n_690) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_668), .Y(n_691) );
AOI222xp33_ASAP7_75t_L g692 ( .A1(n_665), .A2(n_252), .B1(n_266), .B2(n_294), .C1(n_664), .C2(n_671), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_667), .A2(n_252), .B1(n_294), .B2(n_672), .Y(n_693) );
OAI321xp33_ASAP7_75t_L g694 ( .A1(n_673), .A2(n_294), .A3(n_669), .B1(n_663), .B2(n_666), .C(n_652), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_658), .Y(n_695) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_682), .B(n_695), .C(n_678), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_676), .B(n_691), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_679), .Y(n_698) );
A2O1A1Ixp33_ASAP7_75t_L g699 ( .A1(n_678), .A2(n_694), .B(n_689), .C(n_680), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_688), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_696), .B(n_675), .C(n_690), .Y(n_701) );
BUFx2_ASAP7_75t_L g702 ( .A(n_698), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_699), .A2(n_685), .B1(n_683), .B2(n_687), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_702), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_703), .Y(n_705) );
OAI222xp33_ASAP7_75t_L g706 ( .A1(n_705), .A2(n_697), .B1(n_701), .B2(n_700), .C1(n_681), .C2(n_684), .Y(n_706) );
AOI22xp5_ASAP7_75t_SL g707 ( .A1(n_706), .A2(n_704), .B1(n_677), .B2(n_686), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_707), .A2(n_692), .B(n_693), .Y(n_708) );
endmodule