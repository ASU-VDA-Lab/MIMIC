module fake_jpeg_7148_n_331 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_45),
.Y(n_56)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_52),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_48),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_23),
.B1(n_25),
.B2(n_17),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_60),
.Y(n_91)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_61),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_25),
.B(n_28),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_29),
.B(n_33),
.C(n_19),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_35),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_17),
.B1(n_24),
.B2(n_23),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_35),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_53),
.Y(n_78)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_73),
.Y(n_105)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_85),
.B1(n_54),
.B2(n_65),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_76),
.A2(n_87),
.B1(n_89),
.B2(n_94),
.Y(n_100)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_77),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_21),
.Y(n_124)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_47),
.B1(n_48),
.B2(n_58),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_54),
.B1(n_28),
.B2(n_60),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_24),
.B1(n_45),
.B2(n_18),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_86),
.B1(n_65),
.B2(n_20),
.Y(n_113)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_28),
.B1(n_45),
.B2(n_18),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_37),
.B1(n_18),
.B2(n_29),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_29),
.B1(n_33),
.B2(n_19),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_59),
.B(n_50),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_95),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_20),
.B1(n_33),
.B2(n_27),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_115),
.B(n_95),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_59),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_92),
.B1(n_82),
.B2(n_71),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_114),
.Y(n_140)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_108),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_111),
.B1(n_113),
.B2(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_117),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_20),
.B1(n_27),
.B2(n_50),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_56),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_56),
.B(n_51),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_120),
.Y(n_146)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_74),
.A2(n_63),
.B1(n_27),
.B2(n_41),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_51),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_51),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_21),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_124),
.B(n_82),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_126),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_89),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_128),
.A2(n_131),
.B(n_144),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_99),
.Y(n_160)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_87),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_135),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_154),
.Y(n_161)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_138),
.Y(n_184)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

OAI22x1_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_76),
.B1(n_86),
.B2(n_83),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_143),
.B1(n_149),
.B2(n_103),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_84),
.B1(n_85),
.B2(n_70),
.Y(n_143)
);

INVx2_ASAP7_75t_R g144 ( 
.A(n_122),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_84),
.B1(n_71),
.B2(n_79),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_145),
.A2(n_139),
.B1(n_131),
.B2(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_127),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_100),
.A2(n_97),
.B(n_73),
.C(n_51),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_157),
.B(n_112),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_97),
.B1(n_41),
.B2(n_32),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_106),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_116),
.B(n_106),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_21),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_21),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_41),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_159),
.B(n_163),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_21),
.Y(n_210)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_164),
.B(n_172),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_165),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_141),
.B1(n_134),
.B2(n_156),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_130),
.B(n_110),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_179),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_121),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_154),
.C(n_129),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_171),
.A2(n_185),
.B(n_190),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_150),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_177),
.Y(n_206)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_188),
.Y(n_205)
);

BUFx16f_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_127),
.Y(n_183)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_133),
.A2(n_122),
.B(n_112),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_117),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_107),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_136),
.A2(n_122),
.B1(n_119),
.B2(n_32),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

XOR2x2_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_142),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_210),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_202),
.B1(n_204),
.B2(n_216),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_162),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_198),
.B(n_207),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_208),
.C(n_214),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_141),
.B1(n_156),
.B2(n_137),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_164),
.B1(n_176),
.B2(n_191),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_162),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_155),
.C(n_128),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_163),
.A2(n_157),
.B1(n_138),
.B2(n_146),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_209),
.A2(n_178),
.B(n_175),
.C(n_161),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_119),
.C(n_21),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_171),
.A2(n_32),
.B1(n_31),
.B2(n_26),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_31),
.B1(n_26),
.B2(n_3),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_217),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_174),
.A2(n_31),
.B1(n_26),
.B2(n_3),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_218),
.B(n_168),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_175),
.A2(n_31),
.B1(n_26),
.B2(n_3),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_174),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_236),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_211),
.A2(n_180),
.B1(n_173),
.B2(n_165),
.Y(n_224)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

XNOR2x2_ASAP7_75t_SL g229 ( 
.A(n_199),
.B(n_182),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_229),
.B(n_199),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_189),
.C(n_182),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_239),
.C(n_214),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_196),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_232),
.A2(n_245),
.B(n_246),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_233),
.A2(n_216),
.B1(n_219),
.B2(n_204),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_213),
.A2(n_178),
.B(n_169),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_243),
.B(n_212),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_185),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_238),
.Y(n_249)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_186),
.C(n_184),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

BUFx24_ASAP7_75t_SL g241 ( 
.A(n_195),
.Y(n_241)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_184),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_218),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_203),
.B(n_199),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_177),
.B1(n_212),
.B2(n_217),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_206),
.B(n_167),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_251),
.C(n_253),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_233),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_202),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_233),
.B1(n_243),
.B2(n_230),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_239),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_266),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_209),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_263),
.C(n_265),
.Y(n_273)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_194),
.C(n_201),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_226),
.B1(n_223),
.B2(n_235),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_220),
.C(n_159),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_220),
.C(n_181),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_222),
.B(n_181),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_267),
.B(n_240),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_271),
.B1(n_279),
.B2(n_263),
.Y(n_285)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_233),
.B1(n_234),
.B2(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_215),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_277),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_9),
.C(n_4),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_0),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_283),
.B(n_12),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_10),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_282),
.B(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_10),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_288),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_293),
.B(n_7),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_250),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_26),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_247),
.C(n_250),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_291),
.C(n_281),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_281),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_253),
.C(n_267),
.Y(n_291)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_259),
.B(n_251),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_11),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_295),
.B(n_7),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_270),
.B1(n_278),
.B2(n_273),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_9),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_300),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_9),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_260),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_302),
.B(n_305),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_15),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_7),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_306),
.A2(n_307),
.B(n_308),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_2),
.B(n_4),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_5),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_312),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_305),
.A2(n_291),
.B(n_295),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_298),
.B(n_300),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_286),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_318),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_5),
.A3(n_6),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_2),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_322),
.B(n_315),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_303),
.C(n_15),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_14),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_324),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_16),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

NOR2x1_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_311),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_327),
.B1(n_322),
.B2(n_325),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_319),
.B(n_324),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_16),
.Y(n_331)
);


endmodule