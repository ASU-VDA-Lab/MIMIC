module fake_jpeg_27314_n_271 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_44),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_29),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_33),
.B1(n_17),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_54),
.B1(n_57),
.B2(n_59),
.Y(n_85)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_22),
.B1(n_27),
.B2(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_51),
.A2(n_41),
.B1(n_44),
.B2(n_34),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_27),
.B1(n_22),
.B2(n_23),
.Y(n_54)
);

NOR2x1_ASAP7_75t_R g56 ( 
.A(n_45),
.B(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_60),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_61),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_66),
.Y(n_92)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_28),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_43),
.B1(n_38),
.B2(n_40),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_71),
.A2(n_77),
.B1(n_80),
.B2(n_65),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_73),
.B(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_76),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_43),
.B1(n_38),
.B2(n_44),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_79),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_42),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_84),
.Y(n_104)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

CKINVDCx10_ASAP7_75t_R g83 ( 
.A(n_64),
.Y(n_83)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_28),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_41),
.B1(n_53),
.B2(n_50),
.Y(n_115)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_89),
.Y(n_108)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_96),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_35),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_90),
.B(n_91),
.Y(n_123)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_99),
.Y(n_125)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_111),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_72),
.C(n_85),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_77),
.C(n_74),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_16),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_116),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_32),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_74),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_93),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_53),
.B1(n_66),
.B2(n_82),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_85),
.A2(n_79),
.A3(n_72),
.B1(n_92),
.B2(n_71),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_30),
.C(n_18),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_130),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_124),
.B(n_126),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_86),
.B(n_77),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_103),
.B1(n_117),
.B2(n_116),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_134),
.B1(n_135),
.B2(n_55),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_88),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_83),
.B(n_82),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_101),
.B(n_109),
.Y(n_151)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_139),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_67),
.B1(n_61),
.B2(n_49),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_94),
.A2(n_49),
.B1(n_55),
.B2(n_41),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_30),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_142),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_107),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_104),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_141),
.B(n_32),
.Y(n_156)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_129),
.A2(n_100),
.B1(n_118),
.B2(n_110),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_150),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_100),
.B(n_98),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_152),
.B(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_151),
.A2(n_153),
.B(n_160),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_101),
.B(n_34),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_101),
.B(n_99),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_156),
.B(n_136),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_97),
.B1(n_107),
.B2(n_30),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_34),
.B(n_24),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_162),
.C(n_167),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_97),
.C(n_30),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_97),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_122),
.A2(n_0),
.B(n_1),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_165),
.B(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_121),
.A2(n_21),
.B1(n_34),
.B2(n_3),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_21),
.C(n_14),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_21),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_0),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_121),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_145),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_170),
.B(n_179),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_160),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_184),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_136),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_183),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_180),
.B(n_189),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_127),
.C(n_133),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_192),
.C(n_162),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_127),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_124),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

BUFx12_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_191),
.B(n_143),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_195),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

INVxp33_ASAP7_75t_SL g196 ( 
.A(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

OAI322xp33_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_169),
.A3(n_163),
.B1(n_168),
.B2(n_156),
.C1(n_167),
.C2(n_146),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_199),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_161),
.Y(n_198)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_148),
.A3(n_152),
.B1(n_149),
.B2(n_166),
.C1(n_157),
.C2(n_155),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_153),
.B1(n_151),
.B2(n_161),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_175),
.C(n_178),
.Y(n_219)
);

FAx1_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_148),
.CI(n_165),
.CON(n_202),
.SN(n_202)
);

A2O1A1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_202),
.A2(n_171),
.B(n_173),
.C(n_190),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_126),
.B1(n_164),
.B2(n_142),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_210),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_205),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_191),
.B(n_169),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_175),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_182),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_216),
.A2(n_202),
.B1(n_195),
.B2(n_206),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_211),
.C(n_134),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_209),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_226),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_223),
.B(n_224),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_192),
.C(n_191),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_176),
.C(n_187),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_203),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_229),
.A2(n_214),
.B(n_221),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_234),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_207),
.B1(n_204),
.B2(n_188),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_232),
.B1(n_1),
.B2(n_3),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_209),
.B1(n_198),
.B2(n_206),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_213),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_237),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_138),
.C(n_132),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_215),
.C(n_228),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_238),
.B(n_239),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_132),
.C(n_139),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_135),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_1),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_222),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_247),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_238),
.A2(n_227),
.B1(n_225),
.B2(n_228),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_246),
.B(n_248),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_227),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_249),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_250),
.B(n_251),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_234),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_236),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_253),
.A2(n_256),
.B(n_255),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_4),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_252),
.A2(n_247),
.B(n_243),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_257),
.A2(n_258),
.B(n_261),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_252),
.A2(n_4),
.B(n_5),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_260),
.B(n_5),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_254),
.A2(n_4),
.B(n_5),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_259),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_13),
.B(n_8),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

OAI311xp33_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_264),
.A3(n_9),
.B1(n_10),
.C1(n_13),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_268),
.B(n_6),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_269),
.C(n_6),
.Y(n_271)
);


endmodule