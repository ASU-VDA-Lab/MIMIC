module real_jpeg_4763_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_0),
.A2(n_259),
.B1(n_263),
.B2(n_265),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_0),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_0),
.B(n_277),
.C(n_281),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_0),
.B(n_106),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_0),
.B(n_232),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_0),
.B(n_89),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_0),
.B(n_355),
.Y(n_354)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_1),
.Y(n_183)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_1),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_1),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_1),
.Y(n_296)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_1),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_1),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_2),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_2),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_2),
.A2(n_122),
.B1(n_147),
.B2(n_151),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_2),
.A2(n_113),
.B1(n_122),
.B2(n_196),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_2),
.A2(n_122),
.B1(n_298),
.B2(n_435),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_3),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_3),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_3),
.A2(n_94),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_3),
.A2(n_94),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_4),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_4),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_4),
.Y(n_203)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_4),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_4),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g418 ( 
.A(n_4),
.Y(n_418)
);

BUFx5_ASAP7_75t_L g471 ( 
.A(n_4),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_5),
.A2(n_61),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_5),
.A2(n_61),
.B1(n_196),
.B2(n_235),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_5),
.A2(n_61),
.B1(n_401),
.B2(n_402),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_7),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_7),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_7),
.A2(n_245),
.B1(n_288),
.B2(n_292),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_7),
.A2(n_245),
.B1(n_259),
.B2(n_346),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_7),
.A2(n_120),
.B1(n_245),
.B2(n_447),
.Y(n_446)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_8),
.Y(n_520)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_9),
.Y(n_87)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_11),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_11),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_11),
.A2(n_202),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_11),
.A2(n_202),
.B1(n_298),
.B2(n_301),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_11),
.A2(n_175),
.B1(n_202),
.B2(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_12),
.Y(n_300)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_14),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_15),
.A2(n_127),
.B1(n_129),
.B2(n_133),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_15),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_15),
.A2(n_133),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_15),
.A2(n_133),
.B1(n_224),
.B2(n_228),
.Y(n_223)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_17),
.A2(n_196),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_17),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_17),
.A2(n_306),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_17),
.A2(n_306),
.B1(n_393),
.B2(n_394),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_17),
.A2(n_306),
.B1(n_470),
.B2(n_472),
.Y(n_469)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_18),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_18),
.A2(n_53),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_18),
.A2(n_53),
.B1(n_364),
.B2(n_368),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g449 ( 
.A1(n_18),
.A2(n_53),
.B1(n_68),
.B2(n_165),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_518),
.B(n_521),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_208),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_207),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_155),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_24),
.B(n_155),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_134),
.B2(n_135),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_62),
.C(n_95),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_27),
.A2(n_136),
.B1(n_137),
.B2(n_154),
.Y(n_135)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_27),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_27),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_51),
.B1(n_58),
.B2(n_60),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_28),
.A2(n_58),
.B1(n_60),
.B2(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_28),
.A2(n_242),
.B(n_247),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_28),
.A2(n_41),
.B1(n_242),
.B2(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_29),
.B(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_29),
.A2(n_442),
.B(n_443),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_41),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g422 ( 
.A(n_40),
.Y(n_422)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_41),
.B(n_265),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_41)
);

INVx6_ASAP7_75t_L g420 ( 
.A(n_42),
.Y(n_420)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g359 ( 
.A(n_44),
.Y(n_359)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_45),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_46),
.Y(n_128)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_46),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_46),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_46),
.Y(n_394)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_47),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_47),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_47),
.Y(n_425)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_48),
.Y(n_175)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_52),
.B(n_59),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_SL g442 ( 
.A1(n_54),
.A2(n_265),
.B(n_426),
.Y(n_442)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_58),
.A2(n_200),
.B(n_469),
.Y(n_488)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_59),
.B(n_201),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_62),
.A2(n_63),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_62),
.A2(n_63),
.B1(n_95),
.B2(n_96),
.Y(n_157)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_88),
.B(n_90),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_64),
.A2(n_258),
.B(n_266),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_64),
.A2(n_88),
.B1(n_305),
.B2(n_345),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_64),
.A2(n_266),
.B(n_345),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_64),
.A2(n_88),
.B1(n_449),
.B2(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_65),
.A2(n_89),
.B1(n_161),
.B2(n_168),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_65),
.A2(n_89),
.B1(n_161),
.B2(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_65),
.A2(n_89),
.B1(n_195),
.B2(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_65),
.B(n_267),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_77),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_71),
.B1(n_73),
.B2(n_75),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_69),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_69),
.Y(n_197)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_69),
.Y(n_308)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_70),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_70),
.Y(n_375)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_72),
.Y(n_280)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_77),
.A2(n_305),
.B(n_309),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_84),
.B2(n_86),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_82),
.Y(n_284)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_82),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_83),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_83),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_85),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_85),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_85),
.Y(n_229)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_85),
.Y(n_401)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_88),
.A2(n_309),
.B(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_89),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_90),
.Y(n_168)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_93),
.Y(n_270)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_93),
.Y(n_275)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_117),
.B1(n_125),
.B2(n_126),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_97),
.A2(n_125),
.B1(n_126),
.B2(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_97),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_97),
.A2(n_125),
.B1(n_172),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_97),
.A2(n_125),
.B1(n_392),
.B2(n_446),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_106),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_100),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_102),
.Y(n_239)
);

INVx6_ASAP7_75t_L g381 ( 
.A(n_103),
.Y(n_381)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_106),
.A2(n_118),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

AOI22x1_ASAP7_75t_L g474 ( 
.A1(n_106),
.A2(n_170),
.B1(n_396),
.B2(n_475),
.Y(n_474)
);

AO22x2_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B1(n_113),
.B2(n_115),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_112),
.Y(n_348)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_123),
.Y(n_447)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_125),
.B(n_358),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_125),
.A2(n_392),
.B(n_395),
.Y(n_391)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_127),
.Y(n_352)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_145),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_142),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_149),
.Y(n_473)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_150),
.Y(n_429)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_176),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_156),
.B(n_159),
.CI(n_176),
.CON(n_210),
.SN(n_210)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_159),
.A2(n_218),
.B(n_219),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_169),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_167),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_170),
.A2(n_351),
.B(n_357),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_170),
.B(n_396),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_170),
.A2(n_357),
.B(n_491),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI32xp33_ASAP7_75t_L g374 ( 
.A1(n_174),
.A2(n_354),
.A3(n_375),
.B1(n_376),
.B2(n_379),
.Y(n_374)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B(n_198),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_194),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_198),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_178),
.A2(n_194),
.B1(n_216),
.B2(n_458),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_187),
.B(n_189),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_179),
.A2(n_189),
.B1(n_223),
.B2(n_230),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_179),
.A2(n_287),
.B(n_294),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_179),
.A2(n_265),
.B(n_294),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_179),
.A2(n_231),
.B1(n_432),
.B2(n_433),
.Y(n_431)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_180),
.B(n_297),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_180),
.A2(n_295),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_180),
.A2(n_363),
.B1(n_400),
.B2(n_406),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_180),
.A2(n_434),
.B1(n_464),
.B2(n_465),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_183),
.Y(n_407)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_183),
.Y(n_466)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_193),
.Y(n_293)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_193),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_194),
.Y(n_458)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_248),
.B(n_517),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_210),
.B(n_211),
.Y(n_517)
);

BUFx24_ASAP7_75t_SL g526 ( 
.A(n_210),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.C(n_220),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_212),
.A2(n_213),
.B1(n_217),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_217),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_220),
.B(n_477),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_237),
.C(n_241),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_221),
.B(n_456),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_233),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_222),
.B(n_233),
.Y(n_485)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_223),
.Y(n_464)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_227),
.Y(n_291)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_228),
.Y(n_324)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_234),
.Y(n_462)
);

INVx4_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_237),
.B(n_241),
.Y(n_456)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_238),
.Y(n_475)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_247),
.Y(n_443)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI311xp33_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_452),
.A3(n_493),
.B1(n_511),
.C1(n_512),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_410),
.B(n_451),
.Y(n_251)
);

AO21x1_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_383),
.B(n_409),
.Y(n_252)
);

OAI21x1_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_339),
.B(n_382),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_312),
.B(n_338),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_285),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_256),
.B(n_285),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_271),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_257),
.A2(n_271),
.B1(n_272),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_257),
.Y(n_336)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

INVx5_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_SL g351 ( 
.A1(n_265),
.A2(n_352),
.B(n_353),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_265),
.B(n_427),
.Y(n_426)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_284),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_302),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_303),
.C(n_311),
.Y(n_340)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_287),
.Y(n_334)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx8_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_300),
.Y(n_318)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_300),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_310),
.B2(n_311),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp33_ASAP7_75t_SL g379 ( 
.A(n_307),
.B(n_380),
.Y(n_379)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_331),
.B(n_337),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_321),
.B(n_330),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_318),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_329),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_329),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_327),
.B(n_328),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_323),
.Y(n_333)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_328),
.A2(n_362),
.B(n_371),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_335),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_341),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_360),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_349),
.B2(n_350),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_344),
.B(n_349),
.C(n_360),
.Y(n_384)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_358),
.Y(n_396)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_374),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_361),
.B(n_374),
.Y(n_389)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx4_ASAP7_75t_SL g365 ( 
.A(n_366),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_384),
.B(n_385),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_387),
.B1(n_390),
.B2(n_408),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_389),
.C(n_408),
.Y(n_411)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_390),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_397),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_391),
.B(n_398),
.C(n_399),
.Y(n_436)
);

OAI32xp33_ASAP7_75t_L g416 ( 
.A1(n_394),
.A2(n_417),
.A3(n_419),
.B1(n_421),
.B2(n_426),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_400),
.Y(n_432)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_411),
.B(n_412),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_439),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_436),
.B1(n_437),
.B2(n_438),
.Y(n_413)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_414),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_416),
.B1(n_430),
.B2(n_431),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_416),
.B(n_430),
.Y(n_489)
);

INVx8_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_424),
.Y(n_423)
);

INVx6_ASAP7_75t_SL g424 ( 
.A(n_425),
.Y(n_424)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_436),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_436),
.B(n_437),
.C(n_439),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_444),
.B2(n_450),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_440),
.B(n_445),
.C(n_448),
.Y(n_502)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_444),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_445),
.B(n_448),
.Y(n_444)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_446),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_479),
.Y(n_452)
);

A2O1A1Ixp33_ASAP7_75t_SL g512 ( 
.A1(n_453),
.A2(n_479),
.B(n_513),
.C(n_516),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_476),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_454),
.B(n_476),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_457),
.C(n_459),
.Y(n_454)
);

FAx1_ASAP7_75t_SL g492 ( 
.A(n_455),
.B(n_457),
.CI(n_459),
.CON(n_492),
.SN(n_492)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_467),
.C(n_474),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_461),
.B(n_463),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_461),
.B(n_463),
.Y(n_501)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_467),
.A2(n_468),
.B1(n_474),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_474),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_492),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_480),
.B(n_492),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_485),
.C(n_486),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_481),
.A2(n_482),
.B1(n_485),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_485),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_504),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_489),
.C(n_490),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_487),
.A2(n_488),
.B1(n_490),
.B2(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_489),
.B(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_490),
.Y(n_499)
);

BUFx24_ASAP7_75t_SL g525 ( 
.A(n_492),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_494),
.B(n_506),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_495),
.A2(n_514),
.B(n_515),
.Y(n_513)
);

NOR2x1_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_503),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_503),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_500),
.C(n_502),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_509),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_501),
.B1(n_502),
.B2(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_502),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_507),
.B(n_508),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx13_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_520),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_523),
.Y(n_521)
);


endmodule