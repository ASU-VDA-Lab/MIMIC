module real_jpeg_17016_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_611;
wire n_221;
wire n_489;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_602;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_597;
wire n_42;
wire n_268;
wire n_313;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_2),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_2),
.Y(n_123)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_2),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_3),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_3),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_3),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_4),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_4),
.A2(n_116),
.B1(n_218),
.B2(n_222),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_4),
.A2(n_116),
.B1(n_338),
.B2(n_341),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g554 ( 
.A1(n_4),
.A2(n_116),
.B1(n_152),
.B2(n_555),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_5),
.A2(n_167),
.B1(n_171),
.B2(n_173),
.Y(n_166)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_5),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_5),
.A2(n_173),
.B1(n_315),
.B2(n_318),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_5),
.A2(n_99),
.B1(n_173),
.B2(n_546),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_SL g596 ( 
.A1(n_5),
.A2(n_173),
.B1(n_597),
.B2(n_602),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_6),
.B(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_6),
.A2(n_91),
.B(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_6),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_6),
.B(n_79),
.Y(n_411)
);

OAI32xp33_ASAP7_75t_L g414 ( 
.A1(n_6),
.A2(n_415),
.A3(n_417),
.B1(n_420),
.B2(n_422),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g433 ( 
.A1(n_6),
.A2(n_304),
.B1(n_338),
.B2(n_434),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_6),
.A2(n_103),
.B1(n_500),
.B2(n_505),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_7),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_7),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g456 ( 
.A(n_7),
.Y(n_456)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_7),
.Y(n_466)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_8),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_8),
.A2(n_38),
.B1(n_240),
.B2(n_244),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_8),
.A2(n_38),
.B1(n_300),
.B2(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_8),
.A2(n_38),
.B1(n_198),
.B2(n_440),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_9),
.A2(n_149),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_9),
.A2(n_160),
.B1(n_262),
.B2(n_267),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_9),
.A2(n_160),
.B1(n_392),
.B2(n_395),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g482 ( 
.A1(n_9),
.A2(n_160),
.B1(n_483),
.B2(n_485),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_10),
.Y(n_115)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_10),
.Y(n_129)
);

BUFx4f_ASAP7_75t_L g170 ( 
.A(n_10),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_11),
.A2(n_147),
.B1(n_152),
.B2(n_154),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_11),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_11),
.A2(n_154),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_11),
.A2(n_154),
.B1(n_386),
.B2(n_389),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_11),
.A2(n_154),
.B1(n_501),
.B2(n_503),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_12),
.A2(n_171),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_12),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_12),
.A2(n_184),
.B1(n_360),
.B2(n_363),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_12),
.A2(n_184),
.B1(n_291),
.B2(n_569),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g611 ( 
.A1(n_12),
.A2(n_184),
.B1(n_612),
.B2(n_613),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_21),
.B(n_23),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_14),
.A2(n_199),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_14),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_14),
.A2(n_230),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_14),
.A2(n_230),
.B1(n_296),
.B2(n_300),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_14),
.A2(n_230),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_16),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_16),
.Y(n_216)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_16),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_16),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_16),
.Y(n_388)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_16),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_16),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_17),
.A2(n_114),
.B1(n_125),
.B2(n_130),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_17),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_17),
.A2(n_130),
.B1(n_198),
.B2(n_203),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_17),
.A2(n_130),
.B1(n_249),
.B2(n_356),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g564 ( 
.A1(n_17),
.A2(n_130),
.B1(n_330),
.B2(n_565),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_18),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_18),
.A2(n_74),
.B1(n_222),
.B2(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_18),
.A2(n_74),
.B1(n_330),
.B2(n_333),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_18),
.A2(n_74),
.B1(n_407),
.B2(n_408),
.Y(n_406)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_19),
.Y(n_139)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_19),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_19),
.Y(n_153)
);

BUFx8_ASAP7_75t_L g159 ( 
.A(n_19),
.Y(n_159)
);

BUFx12f_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_622),
.B(n_626),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_538),
.B(n_615),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_378),
.B(n_533),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_307),
.C(n_347),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_253),
.B(n_282),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_29),
.B(n_253),
.C(n_535),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_161),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_30),
.B(n_162),
.C(n_225),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_81),
.C(n_131),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_31),
.A2(n_131),
.B1(n_132),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_31),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_42),
.B1(n_69),
.B2(n_79),
.Y(n_31)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_32),
.Y(n_270)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_34),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_35),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_37),
.Y(n_266)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_41),
.Y(n_436)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_42),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_42),
.A2(n_79),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

OAI21xp33_ASAP7_75t_SL g592 ( 
.A1(n_42),
.A2(n_79),
.B(n_593),
.Y(n_592)
);

OA21x2_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_51),
.B(n_58),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_50),
.Y(n_292)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_50),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g422 ( 
.A(n_51),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_55),
.Y(n_356)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_57),
.Y(n_142)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_57),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_63),
.B2(n_66),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_62),
.Y(n_317)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_65),
.Y(n_202)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_65),
.Y(n_397)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_69),
.Y(n_246)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_76),
.Y(n_416)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_77),
.Y(n_252)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_78),
.Y(n_571)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_80),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_80),
.A2(n_247),
.B1(n_261),
.B2(n_270),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_80),
.A2(n_247),
.B1(n_261),
.B2(n_289),
.Y(n_288)
);

OAI22x1_ASAP7_75t_L g336 ( 
.A1(n_80),
.A2(n_247),
.B1(n_248),
.B2(n_337),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_80),
.A2(n_247),
.B1(n_289),
.B2(n_433),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_80),
.A2(n_247),
.B1(n_355),
.B2(n_545),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_80),
.A2(n_247),
.B1(n_545),
.B2(n_568),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_81),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_102),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_82),
.B(n_102),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_90),
.B1(n_94),
.B2(n_98),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_95),
.Y(n_94)
);

AO21x2_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_134),
.B(n_140),
.Y(n_133)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_110),
.B1(n_120),
.B2(n_124),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_103),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_103),
.A2(n_124),
.B1(n_166),
.B2(n_234),
.Y(n_233)
);

AO21x1_ASAP7_75t_L g321 ( 
.A1(n_103),
.A2(n_181),
.B(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_103),
.A2(n_175),
.B1(n_399),
.B2(n_405),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_103),
.A2(n_426),
.B1(n_482),
.B2(n_500),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_105),
.Y(n_427)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_108),
.A2(n_190),
.B1(n_191),
.B2(n_194),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_109),
.Y(n_299)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_109),
.Y(n_470)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_111),
.A2(n_164),
.B1(n_295),
.B2(n_302),
.Y(n_294)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_114),
.Y(n_409)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_115),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_115),
.Y(n_407)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_115),
.Y(n_502)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_122),
.Y(n_302)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_123),
.Y(n_323)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_146),
.B1(n_155),
.B2(n_156),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_133),
.A2(n_155),
.B1(n_156),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_133),
.A2(n_146),
.B1(n_155),
.B2(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_133),
.A2(n_155),
.B1(n_239),
.B2(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_133),
.A2(n_155),
.B1(n_329),
.B2(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_133),
.A2(n_155),
.B1(n_371),
.B2(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_133),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_133),
.A2(n_155),
.B1(n_595),
.B2(n_596),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_133),
.A2(n_155),
.B1(n_596),
.B2(n_611),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_138),
.Y(n_603)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_139),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_139),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_139),
.Y(n_613)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_140),
.A2(n_562),
.B1(n_563),
.B2(n_564),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g623 ( 
.A1(n_140),
.A2(n_563),
.B(n_624),
.Y(n_623)
);

AO22x2_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_142),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_151),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx8_ASAP7_75t_L g612 ( 
.A(n_153),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_155),
.B(n_304),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_159),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_225),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_185),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_163),
.A2(n_186),
.B(n_206),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_174),
.B2(n_180),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_164),
.A2(n_295),
.B1(n_406),
.B2(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_164),
.A2(n_481),
.B1(n_489),
.B2(n_491),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_169),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_169),
.Y(n_504)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_170),
.Y(n_488)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_175),
.B(n_304),
.Y(n_498)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_176),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_206),
.Y(n_185)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_196),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_187),
.A2(n_207),
.B1(n_217),
.B2(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_R g357 ( 
.A1(n_187),
.A2(n_207),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_187),
.A2(n_207),
.B1(n_385),
.B2(n_391),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_187),
.A2(n_207),
.B1(n_391),
.B2(n_439),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_187),
.A2(n_207),
.B1(n_385),
.B2(n_473),
.Y(n_472)
);

OA21x2_ASAP7_75t_L g558 ( 
.A1(n_187),
.A2(n_207),
.B(n_359),
.Y(n_558)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_188),
.A2(n_277),
.B1(n_278),
.B2(n_281),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_188),
.A2(n_197),
.B1(n_277),
.B2(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_188),
.B(n_304),
.Y(n_508)
);

OAI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_188),
.A2(n_277),
.B1(n_278),
.B2(n_524),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_189),
.B(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_193),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_193),
.Y(n_484)
);

OAI22xp33_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_209),
.B1(n_211),
.B2(n_214),
.Y(n_208)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_202),
.Y(n_394)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_217),
.Y(n_206)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_207),
.Y(n_277)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_215),
.Y(n_280)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_221),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_221),
.Y(n_448)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_223),
.Y(n_421)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_224),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_224),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_237),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_226),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_233),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_227),
.A2(n_228),
.B1(n_233),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_229),
.Y(n_281)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_245),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_238),
.B(n_245),
.C(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_242),
.Y(n_332)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_243),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_243),
.Y(n_374)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_244),
.Y(n_372)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.C(n_259),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_254),
.B(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_259),
.Y(n_306)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_271),
.C(n_276),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_276),
.Y(n_285)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_305),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_283),
.B(n_305),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.C(n_287),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_284),
.B(n_530),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_286),
.B(n_287),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_293),
.C(n_303),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_288),
.B(n_518),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_293),
.A2(n_294),
.B1(n_303),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_302),
.Y(n_505)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_303),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_304),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_304),
.B(n_458),
.Y(n_457)
);

OAI21xp33_ASAP7_75t_SL g473 ( 
.A1(n_304),
.A2(n_457),
.B(n_474),
.Y(n_473)
);

A2O1A1O1Ixp25_ASAP7_75t_L g533 ( 
.A1(n_307),
.A2(n_347),
.B(n_534),
.C(n_536),
.D(n_537),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_346),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_308),
.B(n_346),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_309),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_326),
.B1(n_344),
.B2(n_345),
.Y(n_311)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_312),
.B(n_345),
.C(n_377),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_321),
.B1(n_324),
.B2(n_325),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_313),
.B(n_325),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_317),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_320),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_321),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_321),
.B(n_370),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_321),
.A2(n_370),
.B(n_375),
.Y(n_581)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_343),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_336),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_336),
.C(n_343),
.Y(n_349)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_335),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_337),
.Y(n_353)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_376),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_348),
.B(n_376),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_349),
.B(n_584),
.C(n_585),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_366),
.Y(n_350)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_351),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_357),
.B(n_365),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_357),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_365),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_365),
.A2(n_577),
.B1(n_580),
.B2(n_588),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_366),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_368),
.B1(n_369),
.B2(n_375),
.Y(n_366)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_367),
.Y(n_375)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_SL g373 ( 
.A(n_374),
.Y(n_373)
);

AOI21x1_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_528),
.B(n_532),
.Y(n_378)
);

OAI21x1_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_513),
.B(n_527),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_444),
.B(n_512),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_412),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_382),
.B(n_412),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_398),
.C(n_410),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_383),
.A2(n_384),
.B1(n_410),
.B2(n_411),
.Y(n_477)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_387),
.Y(n_390)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_398),
.B(n_477),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_399),
.Y(n_491)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_430),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_413),
.B(n_431),
.C(n_438),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_423),
.B1(n_428),
.B2(n_429),
.Y(n_413)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_414),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_414),
.B(n_429),
.Y(n_522)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_423),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_431),
.A2(n_432),
.B1(n_437),
.B2(n_438),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_439),
.Y(n_524)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

OAI21x1_ASAP7_75t_SL g444 ( 
.A1(n_445),
.A2(n_478),
.B(n_511),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_476),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_446),
.B(n_476),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_471),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_447),
.A2(n_471),
.B1(n_472),
.B2(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_447),
.Y(n_493)
);

OAI32xp33_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_449),
.A3(n_454),
.B1(n_457),
.B2(n_462),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_467),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx8_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_479),
.A2(n_494),
.B(n_510),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_492),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_480),
.B(n_492),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_495),
.A2(n_506),
.B(n_509),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_499),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_507),
.B(n_508),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_514),
.B(n_515),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_516),
.A2(n_517),
.B1(n_520),
.B2(n_521),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_516),
.B(n_523),
.C(n_525),
.Y(n_531)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_522),
.A2(n_523),
.B1(n_525),
.B2(n_526),
.Y(n_521)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_522),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_523),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_529),
.B(n_531),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_529),
.B(n_531),
.Y(n_532)
);

NOR3xp33_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_589),
.C(n_608),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_582),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_541),
.A2(n_618),
.B(n_619),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_SL g541 ( 
.A(n_542),
.B(n_575),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_542),
.B(n_575),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_559),
.Y(n_542)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_543),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_552),
.C(n_558),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_544),
.B(n_558),
.Y(n_578)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_552),
.A2(n_553),
.B1(n_560),
.B2(n_574),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_552),
.A2(n_553),
.B1(n_578),
.B2(n_579),
.Y(n_577)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_553),
.B(n_606),
.C(n_607),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_554),
.Y(n_562)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_558),
.A2(n_567),
.B1(n_572),
.B2(n_573),
.Y(n_566)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_558),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_558),
.B(n_561),
.C(n_573),
.Y(n_604)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_560),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_560),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_566),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_564),
.Y(n_595)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_567),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_568),
.Y(n_593)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx6_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_580),
.C(n_581),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_577),
.Y(n_588)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_578),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_581),
.B(n_587),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_586),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_583),
.B(n_586),
.Y(n_618)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

A2O1A1O1Ixp25_ASAP7_75t_L g616 ( 
.A1(n_590),
.A2(n_609),
.B(n_617),
.C(n_620),
.D(n_621),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_591),
.B(n_605),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_591),
.B(n_605),
.Y(n_620)
);

BUFx24_ASAP7_75t_SL g629 ( 
.A(n_591),
.Y(n_629)
);

FAx1_ASAP7_75t_L g591 ( 
.A(n_592),
.B(n_594),
.CI(n_604),
.CON(n_591),
.SN(n_591)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_592),
.B(n_594),
.C(n_604),
.Y(n_614)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_610),
.B(n_614),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_610),
.B(n_614),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_610),
.B(n_623),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_610),
.B(n_623),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_611),
.Y(n_625)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_625),
.Y(n_624)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);


endmodule