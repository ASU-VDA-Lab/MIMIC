module fake_jpeg_28510_n_535 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_535);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_535;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_3),
.B(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_54),
.Y(n_165)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_17),
.Y(n_55)
);

INVx5_ASAP7_75t_SL g149 ( 
.A(n_55),
.Y(n_149)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_7),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_57),
.B(n_68),
.Y(n_121)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_60),
.Y(n_170)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_64),
.Y(n_174)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_8),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_69),
.Y(n_175)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_48),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_80),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_18),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_101),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_88),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_23),
.B(n_8),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_100),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g101 ( 
.A(n_36),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_104),
.B(n_106),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_108),
.Y(n_154)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_107),
.B(n_18),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_55),
.A2(n_32),
.B1(n_41),
.B2(n_36),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_111),
.A2(n_117),
.B1(n_118),
.B2(n_123),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_57),
.A2(n_68),
.B1(n_37),
.B2(n_30),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_114),
.B(n_136),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_99),
.B1(n_105),
.B2(n_108),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_37),
.B1(n_30),
.B2(n_23),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_41),
.B1(n_49),
.B2(n_25),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_80),
.B(n_52),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_131),
.B(n_158),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_72),
.A2(n_29),
.B(n_43),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_54),
.A2(n_41),
.B1(n_52),
.B2(n_44),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_139),
.A2(n_142),
.B1(n_163),
.B2(n_171),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_98),
.A2(n_50),
.B1(n_26),
.B2(n_44),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_76),
.B(n_50),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_76),
.B(n_49),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_20),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_100),
.B(n_27),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_146),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_71),
.A2(n_31),
.B1(n_27),
.B2(n_40),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_74),
.B(n_13),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_167),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_70),
.A2(n_20),
.B1(n_25),
.B2(n_35),
.Y(n_171)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_176),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_177),
.B(n_178),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_179),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_167),
.A2(n_40),
.B1(n_31),
.B2(n_35),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_187),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_140),
.A2(n_82),
.B1(n_59),
.B2(n_88),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_181),
.A2(n_146),
.B1(n_127),
.B2(n_129),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_46),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_190),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_117),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_185),
.A2(n_195),
.B1(n_215),
.B2(n_141),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_121),
.A2(n_18),
.B1(n_29),
.B2(n_16),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_159),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_189),
.B(n_202),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_112),
.B(n_0),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_193),
.B(n_197),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_81),
.B1(n_75),
.B2(n_77),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

OA22x2_ASAP7_75t_SL g200 ( 
.A1(n_139),
.A2(n_84),
.B1(n_73),
.B2(n_18),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_200),
.A2(n_187),
.B1(n_228),
.B2(n_111),
.Y(n_246)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_201),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_138),
.B(n_18),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_203),
.B(n_213),
.Y(n_241)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_207),
.Y(n_260)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_154),
.B(n_29),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_209),
.B(n_151),
.Y(n_267)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_210),
.B(n_212),
.Y(n_270)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_149),
.B(n_46),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_134),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_119),
.Y(n_214)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_152),
.A2(n_29),
.B1(n_9),
.B2(n_10),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_124),
.A2(n_103),
.B(n_92),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_132),
.B(n_126),
.Y(n_244)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_217),
.B(n_220),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_133),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_219),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_159),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_148),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_222),
.Y(n_264)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_130),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_223),
.Y(n_236)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_224),
.Y(n_253)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_225),
.Y(n_268)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_130),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_116),
.Y(n_265)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_160),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_238),
.A2(n_156),
.B1(n_194),
.B2(n_214),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_243),
.A2(n_174),
.B1(n_160),
.B2(n_229),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_244),
.A2(n_257),
.B(n_132),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_SL g272 ( 
.A1(n_246),
.A2(n_247),
.B(n_200),
.C(n_191),
.Y(n_272)
);

OR2x4_ASAP7_75t_L g247 ( 
.A(n_204),
.B(n_29),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_141),
.B1(n_116),
.B2(n_129),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_184),
.B1(n_228),
.B2(n_200),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_180),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_250),
.B(n_267),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_218),
.A2(n_124),
.B(n_166),
.Y(n_257)
);

CKINVDCx12_ASAP7_75t_R g261 ( 
.A(n_196),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_SL g262 ( 
.A(n_203),
.B(n_204),
.C(n_216),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_183),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_271),
.A2(n_275),
.B1(n_284),
.B2(n_294),
.Y(n_315)
);

AOI32xp33_ASAP7_75t_L g314 ( 
.A1(n_272),
.A2(n_278),
.A3(n_299),
.B1(n_277),
.B2(n_287),
.Y(n_314)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_267),
.B(n_186),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_281),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_236),
.Y(n_325)
);

OAI22x1_ASAP7_75t_SL g278 ( 
.A1(n_246),
.A2(n_191),
.B1(n_143),
.B2(n_219),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_278),
.A2(n_297),
.B1(n_234),
.B2(n_256),
.Y(n_307)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_241),
.B(n_188),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_248),
.A2(n_174),
.B1(n_192),
.B2(n_199),
.Y(n_284)
);

O2A1O1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_244),
.A2(n_198),
.B(n_197),
.C(n_219),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_285),
.Y(n_318)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_286),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_295),
.B(n_300),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_264),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_288),
.B(n_293),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_206),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_289),
.B(n_290),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_201),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_233),
.B(n_176),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_292),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_205),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_237),
.B(n_227),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_257),
.A2(n_225),
.B1(n_224),
.B2(n_221),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_246),
.A2(n_226),
.B1(n_223),
.B2(n_166),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_251),
.Y(n_298)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_231),
.B(n_250),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_302),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_231),
.A2(n_151),
.B(n_126),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_231),
.A2(n_211),
.B(n_143),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_301),
.A2(n_249),
.B(n_263),
.Y(n_328)
);

AND2x2_ASAP7_75t_SL g302 ( 
.A(n_247),
.B(n_168),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_246),
.A2(n_242),
.B1(n_238),
.B2(n_266),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_303),
.A2(n_278),
.B1(n_271),
.B2(n_295),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_307),
.A2(n_326),
.B1(n_294),
.B2(n_284),
.Y(n_340)
);

OAI32xp33_ASAP7_75t_L g311 ( 
.A1(n_274),
.A2(n_258),
.A3(n_234),
.B1(n_236),
.B2(n_232),
.Y(n_311)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_311),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_274),
.B(n_261),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_316),
.C(n_329),
.Y(n_337)
);

XOR2x1_ASAP7_75t_L g353 ( 
.A(n_314),
.B(n_272),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_259),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_302),
.B1(n_301),
.B2(n_300),
.Y(n_335)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_320),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_283),
.A2(n_232),
.B1(n_249),
.B2(n_256),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_321),
.A2(n_328),
.B(n_298),
.Y(n_341)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_286),
.Y(n_323)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_325),
.B(n_327),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_302),
.A2(n_268),
.B1(n_253),
.B2(n_259),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_291),
.B(n_268),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_281),
.B(n_264),
.Y(n_329)
);

OA21x2_ASAP7_75t_L g331 ( 
.A1(n_285),
.A2(n_253),
.B(n_263),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_331),
.A2(n_318),
.B(n_285),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_230),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_302),
.C(n_289),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_326),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_334),
.B(n_339),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_335),
.A2(n_342),
.B1(n_354),
.B2(n_355),
.Y(n_388)
);

AO21x1_ASAP7_75t_L g365 ( 
.A1(n_336),
.A2(n_341),
.B(n_353),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_327),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_340),
.A2(n_347),
.B1(n_359),
.B2(n_315),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_317),
.A2(n_272),
.B1(n_283),
.B2(n_297),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_293),
.Y(n_343)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_343),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_346),
.B(n_309),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_307),
.A2(n_272),
.B1(n_275),
.B2(n_283),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_322),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_230),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_332),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_350),
.B(n_239),
.Y(n_390)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_304),
.Y(n_351)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_351),
.Y(n_379)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_352),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_333),
.A2(n_305),
.B1(n_315),
.B2(n_328),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_305),
.A2(n_272),
.B1(n_292),
.B2(n_280),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_313),
.B(n_290),
.Y(n_356)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_356),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_331),
.A2(n_314),
.B(n_324),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_357),
.A2(n_319),
.B(n_298),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_332),
.A2(n_272),
.B(n_279),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_358),
.A2(n_331),
.B(n_306),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_324),
.A2(n_273),
.B1(n_298),
.B2(n_251),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_288),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_360),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_308),
.B(n_235),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_361),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_312),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_363),
.B(n_364),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_308),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_366),
.A2(n_387),
.B1(n_342),
.B2(n_352),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_337),
.B(n_316),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_368),
.B(n_369),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_311),
.Y(n_369)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_309),
.C(n_306),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_375),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_371),
.A2(n_336),
.B(n_357),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_346),
.B(n_310),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_373),
.C(n_374),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_310),
.C(n_323),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_320),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_376),
.A2(n_336),
.B(n_357),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_319),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_380),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_355),
.B(n_330),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_382),
.Y(n_411)
);

AOI21xp33_ASAP7_75t_L g383 ( 
.A1(n_345),
.A2(n_196),
.B(n_153),
.Y(n_383)
);

OAI21xp33_ASAP7_75t_L g415 ( 
.A1(n_383),
.A2(n_153),
.B(n_351),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_239),
.C(n_252),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_384),
.B(n_361),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_334),
.A2(n_296),
.B1(n_240),
.B2(n_245),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_338),
.A2(n_296),
.B1(n_240),
.B2(n_245),
.Y(n_389)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_389),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_339),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_379),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_392),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_393),
.B(n_410),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_388),
.A2(n_347),
.B1(n_338),
.B2(n_334),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_394),
.A2(n_419),
.B1(n_365),
.B2(n_343),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g427 ( 
.A(n_396),
.Y(n_427)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_367),
.Y(n_398)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_399),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_377),
.B(n_349),
.Y(n_401)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_405),
.Y(n_423)
);

BUFx12_ASAP7_75t_L g403 ( 
.A(n_386),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_413),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_385),
.B(n_350),
.Y(n_404)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_376),
.A2(n_367),
.B(n_362),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_373),
.B(n_356),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_408),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_381),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_366),
.A2(n_342),
.B1(n_354),
.B2(n_335),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_409),
.A2(n_417),
.B1(n_418),
.B2(n_369),
.Y(n_421)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_371),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_412),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_374),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_362),
.A2(n_353),
.B(n_341),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_344),
.C(n_269),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_415),
.B(n_384),
.Y(n_422)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_378),
.A2(n_340),
.B1(n_353),
.B2(n_359),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_421),
.B(n_425),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_433),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_424),
.A2(n_431),
.B1(n_396),
.B2(n_418),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_363),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_419),
.A2(n_365),
.B1(n_344),
.B2(n_348),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_416),
.B(n_375),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_364),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_435),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_416),
.B(n_368),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_395),
.B(n_372),
.C(n_348),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_436),
.B(n_440),
.C(n_441),
.Y(n_445)
);

MAJx2_ASAP7_75t_L g452 ( 
.A(n_438),
.B(n_399),
.C(n_417),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_395),
.B(n_269),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_391),
.B(n_235),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_409),
.A2(n_245),
.B1(n_252),
.B2(n_208),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_402),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_432),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_446),
.Y(n_467)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_437),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_442),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_447),
.Y(n_469)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_420),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_448),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_432),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_449),
.A2(n_457),
.B1(n_404),
.B2(n_411),
.Y(n_465)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_428),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_461),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_431),
.A2(n_410),
.B(n_414),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_451),
.A2(n_454),
.B(n_391),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_452),
.B(n_422),
.Y(n_468)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_406),
.C(n_401),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_456),
.A2(n_458),
.B1(n_460),
.B2(n_462),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_429),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_430),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_424),
.A2(n_397),
.B1(n_412),
.B2(n_398),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_441),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

XOR2x1_ASAP7_75t_SL g464 ( 
.A(n_452),
.B(n_393),
.Y(n_464)
);

AOI21x1_ASAP7_75t_L g491 ( 
.A1(n_464),
.A2(n_474),
.B(n_11),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_466),
.Y(n_483)
);

FAx1_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_405),
.CI(n_421),
.CON(n_466),
.SN(n_466)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_473),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_440),
.C(n_436),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_472),
.C(n_478),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_445),
.B(n_434),
.C(n_435),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_460),
.A2(n_397),
.B1(n_443),
.B2(n_394),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_475),
.B(n_109),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_425),
.C(n_439),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_433),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_480),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_407),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_413),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_481),
.B(n_451),
.C(n_453),
.Y(n_484)
);

MAJx2_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_491),
.C(n_8),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_459),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_492),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_453),
.C(n_411),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_486),
.B(n_490),
.Y(n_504)
);

AND2x2_ASAP7_75t_SL g487 ( 
.A(n_464),
.B(n_403),
.Y(n_487)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_487),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_466),
.A2(n_403),
.B1(n_426),
.B2(n_392),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_488),
.A2(n_6),
.B(n_12),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_467),
.A2(n_477),
.B1(n_466),
.B2(n_470),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_489),
.A2(n_494),
.B1(n_9),
.B2(n_13),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_408),
.C(n_403),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_478),
.A2(n_85),
.B1(n_175),
.B2(n_11),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_46),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_4),
.Y(n_509)
);

NAND4xp25_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_473),
.C(n_468),
.D(n_476),
.Y(n_497)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_497),
.Y(n_516)
);

OAI32xp33_ASAP7_75t_L g498 ( 
.A1(n_488),
.A2(n_481),
.A3(n_479),
.B1(n_46),
.B2(n_42),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_505),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_46),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_499),
.B(n_501),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_487),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_493),
.Y(n_511)
);

NOR3xp33_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_10),
.C(n_13),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_503),
.A2(n_507),
.B(n_11),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_505),
.Y(n_518)
);

AOI21xp33_ASAP7_75t_L g507 ( 
.A1(n_482),
.A2(n_6),
.B(n_12),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_509),
.B(n_508),
.Y(n_514)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_510),
.Y(n_521)
);

AOI21xp33_ASAP7_75t_L g524 ( 
.A1(n_511),
.A2(n_514),
.B(n_518),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_504),
.B(n_486),
.C(n_496),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_513),
.A2(n_515),
.B(n_496),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_502),
.A2(n_484),
.B(n_493),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_519),
.B(n_520),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_516),
.A2(n_503),
.B(n_2),
.Y(n_520)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g522 ( 
.A1(n_512),
.A2(n_42),
.B(n_16),
.C(n_3),
.D(n_2),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_522),
.B(n_523),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_513),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_524),
.A2(n_517),
.B(n_518),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_526),
.A2(n_527),
.B(n_523),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_521),
.A2(n_512),
.B(n_2),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_529),
.A2(n_530),
.B(n_1),
.Y(n_531)
);

OAI311xp33_ASAP7_75t_L g530 ( 
.A1(n_525),
.A2(n_1),
.A3(n_16),
.B1(n_42),
.C1(n_528),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_531),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_1),
.B(n_16),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_16),
.B(n_42),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_42),
.Y(n_535)
);


endmodule