module fake_jpeg_10283_n_26 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_26);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_26;

wire n_21;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_17;
wire n_25;
wire n_15;

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_9),
.A2(n_6),
.B1(n_2),
.B2(n_4),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

NOR3xp33_ASAP7_75t_SL g21 ( 
.A(n_18),
.B(n_7),
.C(n_8),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_22),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_10),
.B(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_15),
.Y(n_25)
);

A2O1A1O1Ixp25_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_16),
.B(n_19),
.C(n_23),
.D(n_24),
.Y(n_26)
);


endmodule