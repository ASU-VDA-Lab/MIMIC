module fake_jpeg_19025_n_204 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_17),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_26),
.B1(n_19),
.B2(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_51),
.B1(n_33),
.B2(n_25),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_19),
.B1(n_26),
.B2(n_17),
.Y(n_51)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_29),
.C(n_36),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_74),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_33),
.B1(n_29),
.B2(n_37),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_67),
.B1(n_41),
.B2(n_45),
.Y(n_81)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_35),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_63),
.C(n_15),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_31),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_46),
.B1(n_47),
.B2(n_41),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_75),
.B1(n_68),
.B2(n_60),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_81),
.A2(n_27),
.B1(n_24),
.B2(n_23),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_42),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_93),
.B(n_28),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_34),
.Y(n_84)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_89),
.C(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_88),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_62),
.B(n_18),
.Y(n_88)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_34),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_42),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_91),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_55),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_112),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_107),
.B1(n_110),
.B2(n_76),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_84),
.C(n_78),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_79),
.C(n_96),
.Y(n_120)
);

OAI22x1_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_61),
.B1(n_64),
.B2(n_68),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_114),
.B1(n_82),
.B2(n_94),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_89),
.B(n_93),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_73),
.B1(n_69),
.B2(n_61),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_73),
.B(n_70),
.C(n_28),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_24),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_0),
.B(n_1),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_23),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_97),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_122),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_111),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_130),
.B1(n_114),
.B2(n_108),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_104),
.C(n_98),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_111),
.C(n_101),
.Y(n_137)
);

AOI221xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_111),
.B1(n_109),
.B2(n_117),
.C(n_113),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_136),
.C(n_135),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_132),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_92),
.B1(n_77),
.B2(n_83),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_85),
.Y(n_133)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_97),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_143),
.C(n_144),
.Y(n_155)
);

BUFx24_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_147),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_118),
.B1(n_106),
.B2(n_125),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_105),
.C(n_106),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_105),
.C(n_106),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_122),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_158),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_125),
.C(n_130),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_163),
.C(n_164),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_119),
.B1(n_121),
.B2(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_142),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_141),
.B1(n_163),
.B2(n_108),
.Y(n_172)
);

XNOR2x1_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_137),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_165),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_135),
.C(n_131),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_115),
.C(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_147),
.B(n_138),
.C(n_145),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_SL g179 ( 
.A(n_167),
.B(n_168),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_154),
.A2(n_138),
.B1(n_139),
.B2(n_148),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_172),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_173),
.A2(n_23),
.B(n_20),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_150),
.B1(n_151),
.B2(n_139),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_155),
.C(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_178),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_155),
.C(n_170),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_110),
.C(n_116),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_182),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_8),
.C(n_4),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_7),
.Y(n_189)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_167),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_184),
.A2(n_187),
.B1(n_4),
.B2(n_5),
.Y(n_193)
);

OAI321xp33_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_169),
.A3(n_168),
.B1(n_173),
.B2(n_6),
.C(n_7),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_8),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_0),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_190),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_7),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_9),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_191),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_4),
.C(n_5),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_192),
.Y(n_197)
);

AOI21x1_ASAP7_75t_L g198 ( 
.A1(n_193),
.A2(n_194),
.B(n_184),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_195),
.A3(n_192),
.B1(n_185),
.B2(n_13),
.C1(n_12),
.C2(n_10),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_199),
.A2(n_200),
.B(n_197),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_196),
.B(n_6),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_6),
.Y(n_202)
);

AOI221xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.C(n_193),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_10),
.C(n_12),
.Y(n_204)
);


endmodule