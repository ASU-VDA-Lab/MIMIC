module real_jpeg_13979_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_3),
.A2(n_62),
.B1(n_69),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_62),
.B1(n_69),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_71),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_7),
.A2(n_62),
.B1(n_69),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_7),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_47),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_8),
.A2(n_36),
.B1(n_37),
.B2(n_47),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_8),
.A2(n_47),
.B1(n_62),
.B2(n_69),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_11),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_80),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_11),
.A2(n_62),
.B1(n_69),
.B2(n_80),
.Y(n_142)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_13),
.A2(n_40),
.B1(n_62),
.B2(n_69),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_14),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_14),
.A2(n_45),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_14),
.B(n_57),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_75),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_14),
.A2(n_37),
.B(n_84),
.C(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_14),
.B(n_41),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_14),
.B(n_66),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_14),
.B(n_97),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_14),
.A2(n_28),
.B(n_31),
.C(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_15),
.A2(n_62),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_15),
.A2(n_36),
.B1(n_37),
.B2(n_68),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_16),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_16),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_16),
.A2(n_30),
.B1(n_62),
.B2(n_69),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_17),
.A2(n_45),
.B1(n_46),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_17),
.A2(n_28),
.B1(n_29),
.B2(n_56),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_17),
.A2(n_36),
.B1(n_37),
.B2(n_56),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_17),
.A2(n_56),
.B1(n_62),
.B2(n_69),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_129),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_128),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_104),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_22),
.B(n_104),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.C(n_93),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_23),
.B(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_58),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_42),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_25),
.B(n_42),
.C(n_58),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_38),
.B2(n_41),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_27),
.A2(n_35),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_28),
.A2(n_29),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_28),
.B(n_51),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_28),
.A2(n_33),
.A3(n_36),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_29),
.A2(n_45),
.A3(n_52),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_29),
.B(n_75),
.Y(n_150)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_31),
.A2(n_41),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_34),
.B(n_37),
.Y(n_151)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_35),
.A2(n_39),
.B1(n_99),
.B2(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_35),
.A2(n_137),
.B(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_36),
.A2(n_37),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_48),
.B1(n_54),
.B2(n_57),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_44),
.A2(n_49),
.B1(n_50),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_53)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_46),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_49),
.A2(n_50),
.B1(n_55),
.B2(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_72),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_59),
.A2(n_60),
.B1(n_72),
.B2(n_161),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_60)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_61),
.A2(n_66),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_61),
.A2(n_66),
.B1(n_67),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_61),
.A2(n_66),
.B1(n_142),
.B2(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_61),
.A2(n_66),
.B1(n_153),
.B2(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_61),
.A2(n_66),
.B1(n_75),
.B2(n_193),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_61),
.A2(n_66),
.B1(n_186),
.B2(n_193),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_69),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_62),
.B(n_195),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_65),
.A2(n_89),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_69),
.A2(n_75),
.B(n_85),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_72),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_76),
.B(n_93),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_88),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_88),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_82),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_81),
.A2(n_86),
.B1(n_145),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_97),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_82),
.A2(n_96),
.B1(n_97),
.B2(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_82),
.A2(n_97),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_82),
.A2(n_97),
.B1(n_172),
.B2(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.C(n_101),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_101),
.B(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_127),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_116),
.B1(n_125),
.B2(n_126),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_106),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_115),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_225),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_221),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_164),
.B(n_220),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_154),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_133),
.B(n_154),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_143),
.C(n_146),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_134),
.B(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_140),
.C(n_141),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_143),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_148),
.A2(n_149),
.B1(n_152),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_150),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_159),
.B2(n_163),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_155),
.B(n_160),
.C(n_162),
.Y(n_222)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_214),
.B(n_219),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_202),
.B(n_213),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_182),
.B(n_201),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_168),
.B(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_178),
.C(n_180),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_181),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_190),
.B(n_200),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_184),
.B(n_188),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_196),
.B(n_199),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_197),
.B(n_198),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_203),
.B(n_204),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_211),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_209),
.C(n_211),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_215),
.B(n_216),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_223),
.Y(n_225)
);


endmodule