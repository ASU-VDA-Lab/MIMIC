module fake_jpeg_11181_n_91 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_40),
.B1(n_34),
.B2(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_40),
.B1(n_37),
.B2(n_31),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_34),
.B1(n_24),
.B2(n_31),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_47),
.B1(n_27),
.B2(n_26),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_32),
.B1(n_27),
.B2(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_50),
.Y(n_58)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_55),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_0),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NAND2xp67_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_48),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_62),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_42),
.B(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_64),
.Y(n_71)
);

NOR3xp33_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_3),
.C(n_4),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_3),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_14),
.Y(n_67)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_67),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_51),
.B1(n_52),
.B2(n_12),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_74),
.B1(n_7),
.B2(n_8),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_5),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_51),
.B1(n_6),
.B2(n_7),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_5),
.C(n_6),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_77),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_22),
.C(n_15),
.Y(n_78)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

A2O1A1O1Ixp25_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_16),
.B(n_19),
.C(n_11),
.D(n_8),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_80),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_80),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_70),
.B(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_79),
.B(n_71),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_74),
.C(n_83),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_81),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_10),
.Y(n_91)
);


endmodule