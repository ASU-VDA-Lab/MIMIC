module fake_netlist_6_421_n_1800 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1800);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1800;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1737;
wire n_236;
wire n_653;
wire n_1464;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_13),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_98),
.Y(n_174)
);

BUFx10_ASAP7_75t_L g175 ( 
.A(n_79),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_53),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_63),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_3),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_41),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_123),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_3),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_55),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_33),
.Y(n_183)
);

BUFx8_ASAP7_75t_SL g184 ( 
.A(n_162),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_35),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_73),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_2),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_97),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_140),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_16),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_133),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_85),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_66),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_22),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_39),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_115),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_53),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_39),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_77),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_121),
.Y(n_201)
);

BUFx2_ASAP7_75t_SL g202 ( 
.A(n_163),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_117),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_141),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_82),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_84),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_50),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_143),
.Y(n_208)
);

BUFx8_ASAP7_75t_SL g209 ( 
.A(n_14),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_75),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_150),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_60),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_114),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_44),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_30),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_6),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_90),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_142),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_167),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_169),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_68),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_160),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_87),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_96),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_1),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_130),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_14),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_131),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_148),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_81),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_124),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_166),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_125),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_127),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_51),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_144),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_101),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_42),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_28),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_61),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_99),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_16),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_13),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_27),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_42),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_132),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_45),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_128),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_136),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_51),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_22),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_78),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_72),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_161),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_103),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_102),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_0),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_105),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_4),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_138),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_33),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_159),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_23),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_69),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_122),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_4),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_28),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_45),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_106),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_34),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_152),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_35),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_49),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_147),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_44),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_155),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_5),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_153),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_27),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_158),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_34),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_107),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_20),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_164),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_7),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_120),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_32),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_62),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_91),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_8),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_86),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_110),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_7),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_11),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_111),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_31),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_80),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_32),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_95),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_10),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_58),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_48),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_50),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_118),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_71),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_126),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_129),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_0),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_149),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_52),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_55),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_108),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_10),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_24),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_15),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_29),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_36),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_41),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_93),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_65),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_113),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_19),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_29),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_88),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_26),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_17),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_70),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_154),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_25),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_31),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_92),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_8),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_145),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_2),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_59),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_24),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_59),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_209),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_217),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_173),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_243),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_243),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_319),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_184),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_243),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_214),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_203),
.B(n_1),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_268),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_239),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_268),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_258),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_173),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_173),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_173),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_173),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_216),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_260),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_216),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_212),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_216),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_216),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_216),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_262),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_223),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_292),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_206),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_251),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_218),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_251),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_251),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_219),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_251),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_269),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_273),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_276),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_251),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_278),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_326),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_280),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_326),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_326),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_190),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_203),
.B(n_5),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_282),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_207),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_215),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_227),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_235),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_225),
.B(n_6),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_238),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_181),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_291),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_242),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_223),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_246),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_221),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_248),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_222),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_264),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_181),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_267),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_271),
.Y(n_405)
);

NOR2xp67_ASAP7_75t_L g406 ( 
.A(n_304),
.B(n_9),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_277),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_295),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_274),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_224),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_208),
.B(n_236),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_277),
.Y(n_412)
);

NAND2xp33_ASAP7_75t_R g413 ( 
.A(n_170),
.B(n_174),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_226),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_179),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_297),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_179),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_172),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_231),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_299),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_304),
.B(n_9),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_208),
.B(n_11),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_244),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_244),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_345),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_341),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_341),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_236),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_354),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g430 ( 
.A1(n_354),
.A2(n_252),
.B(n_284),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_211),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_211),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_355),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_367),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_355),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_369),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_340),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_344),
.B(n_171),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_356),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_403),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_413),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_356),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_344),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_357),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_372),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_347),
.B(n_171),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_357),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_359),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_170),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_174),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_342),
.B(n_229),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_359),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_347),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_360),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_361),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_399),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_361),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_362),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_362),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_350),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_406),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_343),
.B(n_229),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_350),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_363),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_363),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_366),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_348),
.B(n_261),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_401),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_368),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_368),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_365),
.B(n_397),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_353),
.Y(n_473)
);

BUFx8_ASAP7_75t_L g474 ( 
.A(n_349),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_370),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_373),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_377),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_346),
.B(n_306),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_381),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_410),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_382),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_414),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_383),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_384),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_419),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_415),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_415),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_339),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_417),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_417),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_423),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_422),
.B(n_189),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_407),
.B(n_180),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_424),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_352),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_423),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_339),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g500 ( 
.A1(n_424),
.A2(n_252),
.B(n_286),
.Y(n_500)
);

AO22x2_ASAP7_75t_L g501 ( 
.A1(n_442),
.A2(n_316),
.B1(n_308),
.B2(n_306),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_427),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_442),
.B(n_352),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_386),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_427),
.Y(n_505)
);

AND2x2_ASAP7_75t_SL g506 ( 
.A(n_428),
.B(n_308),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_447),
.A2(n_358),
.B1(n_420),
.B2(n_416),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_500),
.Y(n_508)
);

AND2x6_ASAP7_75t_L g509 ( 
.A(n_431),
.B(n_261),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_462),
.B(n_358),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_472),
.B(n_364),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_500),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_364),
.Y(n_513)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_500),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_500),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_427),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_472),
.B(n_261),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_454),
.Y(n_518)
);

BUFx4f_ASAP7_75t_L g519 ( 
.A(n_500),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_431),
.B(n_261),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_473),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_427),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_464),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_462),
.Y(n_524)
);

NAND3xp33_ASAP7_75t_L g525 ( 
.A(n_428),
.B(n_375),
.C(n_374),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_430),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_468),
.A2(n_316),
.B1(n_392),
.B2(n_421),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_427),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_433),
.Y(n_529)
);

NAND3xp33_ASAP7_75t_L g530 ( 
.A(n_451),
.B(n_375),
.C(n_374),
.Y(n_530)
);

AND3x2_ASAP7_75t_L g531 ( 
.A(n_444),
.B(n_294),
.C(n_288),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_436),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_455),
.Y(n_533)
);

NOR3xp33_ASAP7_75t_SL g534 ( 
.A(n_495),
.B(n_185),
.C(n_182),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_451),
.B(n_376),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_468),
.A2(n_430),
.B1(n_432),
.B2(n_431),
.Y(n_536)
);

NOR2x1p5_ASAP7_75t_L g537 ( 
.A(n_434),
.B(n_376),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_450),
.B(n_378),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_450),
.B(n_378),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_436),
.B(n_380),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_430),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_468),
.A2(n_330),
.B1(n_323),
.B2(n_318),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_464),
.B(n_176),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_433),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_468),
.B(n_431),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_444),
.B(n_454),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_432),
.B(n_261),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_433),
.Y(n_548)
);

CKINVDCx6p67_ASAP7_75t_R g549 ( 
.A(n_455),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_439),
.B(n_380),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_441),
.B(n_387),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_433),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_482),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_468),
.A2(n_338),
.B1(n_311),
.B2(n_409),
.Y(n_554)
);

OR2x6_ASAP7_75t_L g555 ( 
.A(n_461),
.B(n_202),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_468),
.B(n_387),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_468),
.B(n_395),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_468),
.B(n_395),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_433),
.Y(n_559)
);

BUFx4f_ASAP7_75t_L g560 ( 
.A(n_461),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_445),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_476),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_476),
.B(n_408),
.Y(n_563)
);

BUFx4f_ASAP7_75t_L g564 ( 
.A(n_497),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_SL g565 ( 
.A(n_441),
.B(n_408),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_477),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_430),
.A2(n_396),
.B1(n_405),
.B2(n_404),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_477),
.Y(n_568)
);

INVx6_ASAP7_75t_L g569 ( 
.A(n_474),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_445),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_432),
.B(n_416),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_478),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_497),
.B(n_420),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_432),
.B(n_310),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_430),
.A2(n_402),
.B1(n_400),
.B2(n_398),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_463),
.A2(n_393),
.B1(n_391),
.B2(n_390),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_452),
.B(n_310),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_463),
.A2(n_389),
.B1(n_388),
.B2(n_385),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_438),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_443),
.B(n_220),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_445),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_478),
.B(n_351),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_480),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_480),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_463),
.A2(n_310),
.B1(n_334),
.B2(n_332),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_485),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_445),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_485),
.B(n_234),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_443),
.B(n_263),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_437),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_452),
.B(n_310),
.Y(n_591)
);

AND2x6_ASAP7_75t_L g592 ( 
.A(n_452),
.B(n_310),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_446),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_445),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_449),
.B(n_232),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_463),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_479),
.A2(n_301),
.B1(n_312),
.B2(n_309),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_479),
.A2(n_265),
.B1(n_245),
.B2(n_247),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_479),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_488),
.B(n_177),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_449),
.B(n_180),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_425),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_457),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_448),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_496),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_453),
.B(n_186),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_456),
.B(n_186),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_467),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_448),
.Y(n_609)
);

INVxp33_ASAP7_75t_L g610 ( 
.A(n_488),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_456),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_474),
.A2(n_200),
.B1(n_188),
.B2(n_328),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_458),
.B(n_240),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_492),
.B(n_204),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_458),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_448),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_459),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_474),
.A2(n_188),
.B1(n_328),
.B2(n_322),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_469),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_460),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_496),
.B(n_205),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_448),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_496),
.B(n_210),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_470),
.B(n_241),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_471),
.B(n_191),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_471),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_435),
.B(n_249),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_L g628 ( 
.A(n_496),
.B(n_191),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_435),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_492),
.A2(n_333),
.B1(n_182),
.B2(n_327),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_496),
.B(n_213),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_489),
.B(n_228),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_L g633 ( 
.A(n_496),
.B(n_192),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_435),
.B(n_192),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_435),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_489),
.B(n_491),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_466),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_440),
.B(n_230),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_466),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_440),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_489),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_440),
.B(n_466),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_536),
.B(n_196),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_506),
.B(n_440),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_506),
.B(n_466),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_523),
.B(n_484),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_535),
.B(n_466),
.Y(n_647)
);

OAI221xp5_ASAP7_75t_L g648 ( 
.A1(n_504),
.A2(n_183),
.B1(n_331),
.B2(n_293),
.C(n_253),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_636),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_508),
.A2(n_512),
.B1(n_515),
.B2(n_542),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_538),
.B(n_481),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_538),
.B(n_481),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_539),
.B(n_481),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_511),
.B(n_503),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_526),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_641),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_542),
.A2(n_302),
.B1(n_178),
.B2(n_314),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_539),
.B(n_481),
.Y(n_658)
);

BUFx8_ASAP7_75t_L g659 ( 
.A(n_518),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_514),
.B(n_536),
.Y(n_660)
);

INVx8_ASAP7_75t_L g661 ( 
.A(n_546),
.Y(n_661)
);

BUFx6f_ASAP7_75t_SL g662 ( 
.A(n_602),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_514),
.B(n_483),
.Y(n_663)
);

AO22x1_ASAP7_75t_L g664 ( 
.A1(n_503),
.A2(n_550),
.B1(n_510),
.B2(n_563),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_634),
.B(n_483),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_526),
.B(n_483),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_596),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_526),
.Y(n_668)
);

NOR3xp33_ASAP7_75t_L g669 ( 
.A(n_565),
.B(n_467),
.C(n_487),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_519),
.A2(n_237),
.B(n_313),
.C(n_321),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_527),
.A2(n_298),
.B1(n_233),
.B2(n_259),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_519),
.B(n_196),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_526),
.B(n_279),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_541),
.B(n_196),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_543),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_525),
.B(n_563),
.C(n_530),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_541),
.B(n_287),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_541),
.B(n_527),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_571),
.B(n_474),
.C(n_193),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_541),
.B(n_289),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_513),
.B(n_196),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_524),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_611),
.B(n_307),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_554),
.A2(n_196),
.B1(n_329),
.B2(n_187),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_556),
.B(n_196),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_615),
.B(n_491),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_610),
.B(n_195),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_617),
.B(n_620),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_610),
.A2(n_498),
.B(n_493),
.C(n_491),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_554),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_540),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_626),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_SL g693 ( 
.A(n_569),
.B(n_557),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_558),
.B(n_196),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_545),
.B(n_250),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_585),
.A2(n_305),
.B1(n_193),
.B2(n_197),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_585),
.A2(n_305),
.B1(n_197),
.B2(n_200),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_560),
.B(n_490),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_599),
.B(n_493),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_532),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_550),
.B(n_201),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_521),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_507),
.B(n_254),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_551),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_595),
.A2(n_290),
.B1(n_272),
.B2(n_255),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_613),
.B(n_624),
.Y(n_706)
);

OAI221xp5_ASAP7_75t_L g707 ( 
.A1(n_598),
.A2(n_309),
.B1(n_303),
.B2(n_198),
.C(n_199),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_580),
.B(n_201),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_562),
.B(n_426),
.Y(n_709)
);

INVx6_ASAP7_75t_L g710 ( 
.A(n_602),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_555),
.A2(n_300),
.B1(n_256),
.B2(n_257),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_629),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_635),
.B(n_266),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_566),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_640),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_564),
.B(n_270),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_501),
.A2(n_315),
.B1(n_185),
.B2(n_187),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_568),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_572),
.B(n_426),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_583),
.B(n_426),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_589),
.B(n_320),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_584),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_574),
.B(n_564),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_586),
.B(n_429),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_587),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_627),
.B(n_281),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_567),
.B(n_283),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_517),
.B(n_429),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_567),
.B(n_285),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_601),
.B(n_606),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_632),
.Y(n_731)
);

A2O1A1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_588),
.A2(n_601),
.B(n_606),
.C(n_625),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_501),
.A2(n_335),
.B1(n_303),
.B2(n_312),
.Y(n_733)
);

AND3x1_ASAP7_75t_L g734 ( 
.A(n_534),
.B(n_195),
.C(n_315),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_587),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_632),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_501),
.A2(n_598),
.B1(n_575),
.B2(n_638),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_575),
.B(n_296),
.Y(n_738)
);

OR2x4_ASAP7_75t_L g739 ( 
.A(n_573),
.B(n_324),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_622),
.Y(n_740)
);

AND2x6_ASAP7_75t_SL g741 ( 
.A(n_546),
.B(n_499),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_642),
.B(n_320),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_505),
.B(n_322),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_582),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_588),
.B(n_171),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_638),
.A2(n_327),
.B1(n_194),
.B2(n_317),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_612),
.B(n_175),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_607),
.B(n_465),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_607),
.B(n_465),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_582),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_637),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_546),
.B(n_194),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_625),
.B(n_337),
.Y(n_753)
);

AND2x6_ASAP7_75t_SL g754 ( 
.A(n_555),
.B(n_337),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_574),
.Y(n_755)
);

AO221x1_ASAP7_75t_L g756 ( 
.A1(n_597),
.A2(n_175),
.B1(n_275),
.B2(n_325),
.C(n_324),
.Y(n_756)
);

INVx5_ASAP7_75t_L g757 ( 
.A(n_509),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_605),
.B(n_465),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_639),
.B(n_486),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_621),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_638),
.B(n_333),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_618),
.B(n_317),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_502),
.B(n_486),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_502),
.B(n_486),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_531),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_522),
.B(n_325),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_637),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_600),
.B(n_614),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_590),
.Y(n_769)
);

NAND3xp33_ASAP7_75t_SL g770 ( 
.A(n_534),
.B(n_336),
.C(n_335),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_638),
.A2(n_336),
.B1(n_325),
.B2(n_275),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_621),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_623),
.A2(n_475),
.B(n_275),
.C(n_175),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_579),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_623),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_603),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_639),
.B(n_475),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_516),
.B(n_475),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_600),
.B(n_12),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_516),
.B(n_165),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_529),
.B(n_157),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_600),
.A2(n_146),
.B1(n_139),
.B2(n_137),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_614),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_529),
.B(n_135),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_614),
.B(n_12),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_544),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_528),
.B(n_134),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_631),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_548),
.B(n_119),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_544),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_631),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_552),
.B(n_112),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_533),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_630),
.B(n_15),
.Y(n_794)
);

BUFx8_ASAP7_75t_L g795 ( 
.A(n_608),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_559),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_654),
.B(n_552),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_655),
.A2(n_581),
.B(n_570),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_732),
.A2(n_633),
.B(n_628),
.C(n_578),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_654),
.B(n_561),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_730),
.B(n_561),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_706),
.B(n_604),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_655),
.A2(n_581),
.B(n_570),
.Y(n_803)
);

BUFx12f_ASAP7_75t_L g804 ( 
.A(n_659),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_655),
.B(n_668),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_706),
.B(n_604),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_668),
.A2(n_609),
.B(n_616),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_699),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_668),
.B(n_619),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_666),
.A2(n_616),
.B(n_594),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_660),
.A2(n_643),
.B(n_753),
.C(n_701),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_678),
.A2(n_569),
.B1(n_537),
.B2(n_593),
.Y(n_812)
);

NOR2x1_ASAP7_75t_L g813 ( 
.A(n_676),
.B(n_553),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_673),
.A2(n_616),
.B(n_594),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_677),
.A2(n_616),
.B(n_594),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_687),
.B(n_549),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_646),
.B(n_576),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_701),
.A2(n_638),
.B1(n_577),
.B2(n_592),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_680),
.A2(n_594),
.B(n_576),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_674),
.A2(n_663),
.B(n_672),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_744),
.B(n_592),
.Y(n_821)
);

AOI21x1_ASAP7_75t_L g822 ( 
.A1(n_672),
.A2(n_592),
.B(n_591),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_691),
.B(n_569),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_643),
.A2(n_592),
.B1(n_591),
.B2(n_577),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_731),
.B(n_592),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_647),
.A2(n_547),
.B(n_520),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_664),
.B(n_17),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_650),
.A2(n_737),
.B1(n_750),
.B2(n_651),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_753),
.B(n_591),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_675),
.B(n_18),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_674),
.A2(n_591),
.B(n_577),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_740),
.A2(n_547),
.B(n_520),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_649),
.B(n_577),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_740),
.A2(n_547),
.B(n_520),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_644),
.A2(n_650),
.B(n_645),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_700),
.Y(n_836)
);

OAI21xp5_ASAP7_75t_L g837 ( 
.A1(n_665),
.A2(n_547),
.B(n_520),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_702),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_704),
.B(n_18),
.Y(n_839)
);

NOR2xp67_ASAP7_75t_L g840 ( 
.A(n_769),
.B(n_109),
.Y(n_840)
);

NOR2xp67_ASAP7_75t_L g841 ( 
.A(n_776),
.B(n_104),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_685),
.A2(n_520),
.B(n_509),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_708),
.B(n_509),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_685),
.A2(n_509),
.B(n_100),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_681),
.A2(n_509),
.B1(n_89),
.B2(n_83),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_783),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_737),
.A2(n_76),
.B1(n_74),
.B2(n_67),
.Y(n_847)
);

AOI21x1_ASAP7_75t_L g848 ( 
.A1(n_694),
.A2(n_64),
.B(n_20),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_694),
.A2(n_653),
.B(n_652),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_658),
.A2(n_19),
.B(n_21),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_731),
.B(n_736),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_708),
.B(n_721),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_682),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_727),
.A2(n_21),
.B(n_23),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_681),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_721),
.B(n_36),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_731),
.B(n_37),
.Y(n_857)
);

O2A1O1Ixp5_ASAP7_75t_L g858 ( 
.A1(n_748),
.A2(n_37),
.B(n_38),
.C(n_40),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_749),
.B(n_38),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_762),
.A2(n_58),
.B(n_43),
.C(n_46),
.Y(n_860)
);

AOI21x1_ASAP7_75t_L g861 ( 
.A1(n_695),
.A2(n_40),
.B(n_43),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_688),
.B(n_46),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_695),
.A2(n_47),
.B(n_48),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_671),
.A2(n_49),
.B(n_52),
.C(n_54),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_SL g865 ( 
.A1(n_670),
.A2(n_54),
.B(n_56),
.C(n_57),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_731),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_736),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_755),
.A2(n_56),
.B1(n_57),
.B2(n_736),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_727),
.A2(n_738),
.B(n_729),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_736),
.A2(n_760),
.B1(n_775),
.B2(n_788),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_758),
.A2(n_778),
.B(n_777),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_759),
.A2(n_763),
.B(n_764),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_762),
.A2(n_791),
.B(n_772),
.C(n_794),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_SL g874 ( 
.A(n_745),
.B(n_648),
.C(n_746),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_728),
.A2(n_757),
.B(n_726),
.Y(n_875)
);

BUFx8_ASAP7_75t_SL g876 ( 
.A(n_662),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_714),
.B(n_722),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_757),
.A2(n_726),
.B(n_686),
.Y(n_878)
);

NOR2x1_ASAP7_75t_L g879 ( 
.A(n_679),
.B(n_770),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_710),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_710),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_757),
.A2(n_725),
.B(n_767),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_692),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_757),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_794),
.A2(n_768),
.B(n_718),
.C(n_746),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_689),
.A2(n_712),
.B(n_715),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_735),
.A2(n_751),
.B(n_719),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_667),
.B(n_683),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_709),
.A2(n_724),
.B(n_720),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_742),
.A2(n_713),
.B(n_796),
.Y(n_890)
);

BUFx12f_ASAP7_75t_L g891 ( 
.A(n_659),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_657),
.B(n_710),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_723),
.B(n_771),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_713),
.B(n_705),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_786),
.A2(n_790),
.B(n_780),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_743),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_774),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_768),
.A2(n_703),
.B1(n_716),
.B2(n_761),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_693),
.B(n_789),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_766),
.B(n_733),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_781),
.A2(n_784),
.B(n_792),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_787),
.A2(n_789),
.B(n_716),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_793),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_703),
.A2(n_747),
.B(n_773),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_779),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_717),
.B(n_733),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_684),
.A2(n_771),
.B(n_711),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_661),
.Y(n_908)
);

CKINVDCx16_ASAP7_75t_R g909 ( 
.A(n_698),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_684),
.A2(n_782),
.B(n_765),
.Y(n_910)
);

BUFx8_ASAP7_75t_L g911 ( 
.A(n_662),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_717),
.B(n_697),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_739),
.A2(n_696),
.B(n_785),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_752),
.B(n_707),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_661),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_690),
.B(n_785),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_779),
.A2(n_661),
.B(n_690),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_756),
.B(n_734),
.Y(n_918)
);

NOR2x1p5_ASAP7_75t_SL g919 ( 
.A(n_754),
.B(n_669),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_795),
.A2(n_519),
.B(n_514),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_795),
.B(n_741),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_SL g922 ( 
.A1(n_732),
.A2(n_643),
.B(n_730),
.C(n_672),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_655),
.A2(n_519),
.B(n_514),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_732),
.A2(n_730),
.B(n_504),
.C(n_660),
.Y(n_924)
);

OAI22xp33_ASAP7_75t_L g925 ( 
.A1(n_730),
.A2(n_504),
.B1(n_660),
.B2(n_654),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_654),
.B(n_730),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_654),
.B(n_730),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_654),
.B(n_730),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_699),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_655),
.A2(n_519),
.B(n_514),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_655),
.A2(n_519),
.B(n_514),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_656),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_699),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_732),
.A2(n_730),
.B1(n_678),
.B2(n_660),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_654),
.A2(n_706),
.B1(n_701),
.B2(n_730),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_654),
.B(n_442),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_654),
.B(n_442),
.Y(n_937)
);

AND2x6_ASAP7_75t_L g938 ( 
.A(n_655),
.B(n_668),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_SL g939 ( 
.A(n_769),
.B(n_776),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_732),
.A2(n_654),
.B(n_701),
.C(n_753),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_699),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_732),
.A2(n_730),
.B(n_504),
.C(n_660),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_655),
.B(n_668),
.Y(n_943)
);

AOI21xp33_ASAP7_75t_L g944 ( 
.A1(n_701),
.A2(n_654),
.B(n_753),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_655),
.A2(n_519),
.B(n_514),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_731),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_699),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_655),
.B(n_668),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_655),
.A2(n_519),
.B(n_514),
.Y(n_949)
);

BUFx8_ASAP7_75t_L g950 ( 
.A(n_662),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_655),
.A2(n_519),
.B(n_514),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_654),
.B(n_442),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_655),
.A2(n_519),
.B(n_514),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_654),
.B(n_730),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_643),
.A2(n_660),
.B1(n_684),
.B2(n_654),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_732),
.A2(n_730),
.B(n_504),
.C(n_660),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_687),
.B(n_442),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_655),
.A2(n_519),
.B(n_514),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_732),
.A2(n_654),
.B(n_701),
.C(n_753),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_654),
.B(n_730),
.Y(n_960)
);

AO32x1_ASAP7_75t_L g961 ( 
.A1(n_671),
.A2(n_236),
.A3(n_208),
.B1(n_203),
.B2(n_712),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_655),
.B(n_668),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_655),
.A2(n_519),
.B(n_514),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_923),
.A2(n_931),
.B(n_930),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_895),
.A2(n_872),
.B(n_871),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_935),
.B(n_926),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_945),
.A2(n_951),
.B(n_949),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_957),
.B(n_817),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_936),
.B(n_937),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_927),
.A2(n_928),
.B1(n_960),
.B2(n_954),
.Y(n_970)
);

OAI21x1_ASAP7_75t_L g971 ( 
.A1(n_820),
.A2(n_886),
.B(n_887),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_940),
.A2(n_959),
.B(n_934),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_SL g973 ( 
.A1(n_811),
.A2(n_869),
.B(n_924),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_953),
.A2(n_958),
.B(n_963),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_922),
.A2(n_806),
.B(n_802),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_938),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_925),
.B(n_937),
.Y(n_977)
);

AOI21x1_ASAP7_75t_L g978 ( 
.A1(n_849),
.A2(n_902),
.B(n_800),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_955),
.A2(n_852),
.B1(n_944),
.B2(n_925),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_838),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_932),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_952),
.B(n_852),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_876),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_952),
.B(n_942),
.Y(n_984)
);

AOI221x1_ASAP7_75t_L g985 ( 
.A1(n_904),
.A2(n_827),
.B1(n_874),
.B2(n_918),
.C(n_913),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_810),
.A2(n_803),
.B(n_798),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_956),
.B(n_955),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_874),
.A2(n_914),
.B1(n_892),
.B2(n_898),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_932),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_808),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_875),
.A2(n_807),
.B(n_822),
.Y(n_991)
);

AOI21x1_ASAP7_75t_L g992 ( 
.A1(n_797),
.A2(n_878),
.B(n_801),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_889),
.A2(n_815),
.B(n_814),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_873),
.B(n_916),
.Y(n_994)
);

NAND2x1p5_ASAP7_75t_L g995 ( 
.A(n_880),
.B(n_881),
.Y(n_995)
);

AND2x2_ASAP7_75t_SL g996 ( 
.A(n_909),
.B(n_939),
.Y(n_996)
);

AOI21x1_ASAP7_75t_SL g997 ( 
.A1(n_856),
.A2(n_912),
.B(n_900),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_899),
.A2(n_826),
.B(n_882),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_905),
.B(n_885),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_884),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_929),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_901),
.A2(n_962),
.B(n_948),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_943),
.A2(n_962),
.B(n_948),
.Y(n_1003)
);

AO21x2_ASAP7_75t_L g1004 ( 
.A1(n_893),
.A2(n_835),
.B(n_829),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_804),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_908),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_L g1007 ( 
.A(n_907),
.B(n_827),
.C(n_914),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_910),
.A2(n_917),
.B(n_799),
.C(n_894),
.Y(n_1008)
);

NAND2xp33_ASAP7_75t_SL g1009 ( 
.A(n_880),
.B(n_881),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_828),
.B(n_906),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_896),
.B(n_859),
.Y(n_1011)
);

AO21x1_ASAP7_75t_L g1012 ( 
.A1(n_893),
.A2(n_854),
.B(n_847),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_836),
.B(n_809),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_938),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_933),
.Y(n_1015)
);

INVx1_ASAP7_75t_SL g1016 ( 
.A(n_897),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_846),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_816),
.B(n_830),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_938),
.B(n_877),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_819),
.A2(n_821),
.B(n_837),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_943),
.A2(n_805),
.B(n_843),
.Y(n_1021)
);

INVxp67_ASAP7_75t_SL g1022 ( 
.A(n_851),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_831),
.A2(n_870),
.B(n_833),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_938),
.B(n_888),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_SL g1025 ( 
.A1(n_920),
.A2(n_861),
.B(n_848),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_825),
.A2(n_842),
.B(n_884),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_812),
.B(n_813),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_908),
.B(n_915),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_879),
.A2(n_947),
.B1(n_941),
.B2(n_862),
.Y(n_1029)
);

AO21x1_ASAP7_75t_L g1030 ( 
.A1(n_863),
.A2(n_890),
.B(n_857),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_832),
.A2(n_834),
.B(n_825),
.Y(n_1031)
);

NAND2x1_ASAP7_75t_L g1032 ( 
.A(n_938),
.B(n_884),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_818),
.A2(n_844),
.B(n_858),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_866),
.B(n_867),
.Y(n_1034)
);

CKINVDCx6p67_ASAP7_75t_R g1035 ( 
.A(n_891),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_855),
.A2(n_860),
.B1(n_824),
.B2(n_857),
.Y(n_1036)
);

AND2x6_ASAP7_75t_L g1037 ( 
.A(n_884),
.B(n_866),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_867),
.B(n_946),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_824),
.A2(n_946),
.B(n_883),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_823),
.B(n_839),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_836),
.B(n_846),
.Y(n_1041)
);

BUFx12f_ASAP7_75t_L g1042 ( 
.A(n_911),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_823),
.B(n_853),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_839),
.B(n_840),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_845),
.A2(n_841),
.B(n_868),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_908),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_903),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_858),
.A2(n_850),
.B(n_864),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_865),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_908),
.B(n_919),
.Y(n_1050)
);

NAND2x1_ASAP7_75t_L g1051 ( 
.A(n_921),
.B(n_961),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_921),
.A2(n_911),
.B1(n_950),
.B2(n_961),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_961),
.B(n_950),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_895),
.A2(n_872),
.B(n_871),
.Y(n_1054)
);

AO31x2_ASAP7_75t_L g1055 ( 
.A1(n_940),
.A2(n_959),
.A3(n_934),
.B(n_828),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_895),
.A2(n_872),
.B(n_871),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_938),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_923),
.A2(n_668),
.B(n_655),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_957),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_957),
.B(n_817),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_880),
.B(n_655),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_908),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_895),
.A2(n_872),
.B(n_871),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_923),
.A2(n_668),
.B(n_655),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_957),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_923),
.A2(n_668),
.B(n_655),
.Y(n_1066)
);

INVx5_ASAP7_75t_L g1067 ( 
.A(n_938),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_935),
.A2(n_926),
.B1(n_928),
.B2(n_927),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_940),
.A2(n_959),
.B(n_934),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_957),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_852),
.A2(n_935),
.B(n_944),
.C(n_940),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_940),
.A2(n_959),
.B(n_934),
.Y(n_1072)
);

AO31x2_ASAP7_75t_L g1073 ( 
.A1(n_940),
.A2(n_959),
.A3(n_934),
.B(n_828),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_923),
.A2(n_668),
.B(n_655),
.Y(n_1074)
);

AO31x2_ASAP7_75t_L g1075 ( 
.A1(n_940),
.A2(n_959),
.A3(n_934),
.B(n_828),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_957),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_895),
.A2(n_872),
.B(n_871),
.Y(n_1077)
);

AO31x2_ASAP7_75t_L g1078 ( 
.A1(n_940),
.A2(n_959),
.A3(n_934),
.B(n_828),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_940),
.A2(n_959),
.B(n_934),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_895),
.A2(n_872),
.B(n_871),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_895),
.A2(n_872),
.B(n_871),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_895),
.A2(n_872),
.B(n_871),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_929),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_935),
.B(n_926),
.Y(n_1084)
);

INVx5_ASAP7_75t_L g1085 ( 
.A(n_938),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_923),
.A2(n_668),
.B(n_655),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_923),
.A2(n_668),
.B(n_655),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_895),
.A2(n_872),
.B(n_871),
.Y(n_1088)
);

AOI21x1_ASAP7_75t_SL g1089 ( 
.A1(n_918),
.A2(n_856),
.B(n_912),
.Y(n_1089)
);

AO21x2_ASAP7_75t_L g1090 ( 
.A1(n_869),
.A2(n_959),
.B(n_940),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_884),
.Y(n_1091)
);

AOI211x1_ASAP7_75t_L g1092 ( 
.A1(n_944),
.A2(n_854),
.B(n_927),
.C(n_926),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_936),
.B(n_937),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_895),
.A2(n_872),
.B(n_871),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_936),
.B(n_937),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_940),
.A2(n_959),
.B(n_934),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_884),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_923),
.A2(n_668),
.B(n_655),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_935),
.B(n_926),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_938),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_SL g1101 ( 
.A(n_935),
.B(n_852),
.C(n_523),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_957),
.B(n_817),
.Y(n_1102)
);

BUFx5_ASAP7_75t_L g1103 ( 
.A(n_938),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_895),
.A2(n_872),
.B(n_871),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_936),
.B(n_937),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_935),
.B(n_926),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_876),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_895),
.A2(n_872),
.B(n_871),
.Y(n_1108)
);

OAI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_982),
.A2(n_1095),
.B1(n_1093),
.B2(n_1105),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_969),
.A2(n_1007),
.B(n_1071),
.C(n_982),
.Y(n_1110)
);

BUFx8_ASAP7_75t_L g1111 ( 
.A(n_1042),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1101),
.B(n_1040),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_1016),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_987),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_976),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1028),
.B(n_1050),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_1017),
.Y(n_1117)
);

O2A1O1Ixp5_ASAP7_75t_L g1118 ( 
.A1(n_979),
.A2(n_1012),
.B(n_1048),
.C(n_1079),
.Y(n_1118)
);

INVx5_ASAP7_75t_L g1119 ( 
.A(n_1067),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1028),
.B(n_1050),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_980),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1001),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_990),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_1041),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_L g1125 ( 
.A(n_1047),
.B(n_981),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1015),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_989),
.Y(n_1127)
);

AO32x1_ASAP7_75t_L g1128 ( 
.A1(n_979),
.A2(n_1049),
.A3(n_1036),
.B1(n_1068),
.B2(n_970),
.Y(n_1128)
);

INVx5_ASAP7_75t_L g1129 ( 
.A(n_1067),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_970),
.B(n_1068),
.Y(n_1130)
);

NOR2xp67_ASAP7_75t_L g1131 ( 
.A(n_1044),
.B(n_1018),
.Y(n_1131)
);

OR2x6_ASAP7_75t_L g1132 ( 
.A(n_995),
.B(n_976),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_988),
.A2(n_977),
.B(n_1045),
.C(n_1008),
.Y(n_1133)
);

OA21x2_ASAP7_75t_L g1134 ( 
.A1(n_985),
.A2(n_1069),
.B(n_972),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_966),
.B(n_1084),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_1016),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1084),
.B(n_1099),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_SL g1138 ( 
.A1(n_1048),
.A2(n_1096),
.B(n_1079),
.C(n_972),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1083),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_973),
.A2(n_1096),
.B(n_1069),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_977),
.A2(n_1072),
.B(n_1106),
.C(n_1099),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1072),
.A2(n_975),
.B(n_987),
.Y(n_1142)
);

CKINVDCx11_ASAP7_75t_R g1143 ( 
.A(n_1107),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_1006),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1106),
.A2(n_984),
.B1(n_1092),
.B2(n_999),
.Y(n_1145)
);

NAND2xp33_ASAP7_75t_L g1146 ( 
.A(n_1103),
.B(n_1067),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_1006),
.B(n_1046),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_1059),
.B(n_1065),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_968),
.B(n_1060),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_984),
.A2(n_1081),
.B(n_965),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_994),
.A2(n_1036),
.B1(n_1102),
.B2(n_1010),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1010),
.A2(n_1065),
.B1(n_1070),
.B2(n_1076),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1014),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1031),
.A2(n_964),
.B(n_967),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1059),
.B(n_1070),
.Y(n_1155)
);

BUFx2_ASAP7_75t_SL g1156 ( 
.A(n_1046),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1054),
.A2(n_1080),
.B(n_1077),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1076),
.B(n_996),
.Y(n_1158)
);

BUFx12f_ASAP7_75t_L g1159 ( 
.A(n_1005),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1046),
.Y(n_1160)
);

OR2x6_ASAP7_75t_L g1161 ( 
.A(n_995),
.B(n_1014),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1027),
.A2(n_1090),
.B1(n_1013),
.B2(n_1030),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1011),
.A2(n_1029),
.B(n_1033),
.C(n_1002),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_983),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1043),
.B(n_1062),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1056),
.A2(n_1108),
.B(n_1094),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1062),
.B(n_1022),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1062),
.B(n_1057),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1067),
.B(n_1085),
.Y(n_1169)
);

AOI221x1_ASAP7_75t_L g1170 ( 
.A1(n_1053),
.A2(n_1033),
.B1(n_1023),
.B2(n_974),
.C(n_1025),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1057),
.B(n_1100),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_1053),
.Y(n_1172)
);

CKINVDCx8_ASAP7_75t_R g1173 ( 
.A(n_1037),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1063),
.A2(n_1082),
.B(n_1088),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1024),
.B(n_1019),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1034),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1055),
.B(n_1075),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1035),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1038),
.Y(n_1179)
);

BUFx2_ASAP7_75t_SL g1180 ( 
.A(n_1085),
.Y(n_1180)
);

INVx3_ASAP7_75t_SL g1181 ( 
.A(n_1037),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1019),
.Y(n_1182)
);

OR2x6_ASAP7_75t_L g1183 ( 
.A(n_1100),
.B(n_1061),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1073),
.B(n_1075),
.Y(n_1184)
);

AND2x2_ASAP7_75t_SL g1185 ( 
.A(n_1052),
.B(n_1024),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1051),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1090),
.B(n_1078),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1000),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1000),
.Y(n_1189)
);

BUFx12f_ASAP7_75t_L g1190 ( 
.A(n_1061),
.Y(n_1190)
);

BUFx4f_ASAP7_75t_SL g1191 ( 
.A(n_1037),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1075),
.B(n_1078),
.Y(n_1192)
);

INVx3_ASAP7_75t_SL g1193 ( 
.A(n_1037),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1078),
.B(n_1004),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1085),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1104),
.A2(n_1087),
.B(n_1098),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1091),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1085),
.A2(n_1039),
.B1(n_1032),
.B2(n_1003),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1097),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1058),
.A2(n_1074),
.B1(n_1064),
.B2(n_1066),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1097),
.B(n_1026),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1086),
.A2(n_1020),
.B(n_971),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1103),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1020),
.A2(n_1021),
.B1(n_978),
.B2(n_992),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_SL g1205 ( 
.A1(n_1089),
.A2(n_997),
.B(n_993),
.C(n_1004),
.Y(n_1205)
);

CKINVDCx8_ASAP7_75t_R g1206 ( 
.A(n_1009),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_1103),
.Y(n_1207)
);

CKINVDCx8_ASAP7_75t_R g1208 ( 
.A(n_1103),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1103),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_998),
.B(n_991),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_986),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_969),
.B(n_1093),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_976),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_969),
.B(n_1093),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1006),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_973),
.A2(n_1008),
.B(n_972),
.Y(n_1216)
);

BUFx10_ASAP7_75t_L g1217 ( 
.A(n_983),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_973),
.A2(n_1008),
.B(n_972),
.Y(n_1218)
);

INVx4_ASAP7_75t_L g1219 ( 
.A(n_1006),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_973),
.A2(n_1008),
.B(n_972),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_968),
.B(n_1102),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1028),
.B(n_908),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_980),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_980),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1006),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1041),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_968),
.B(n_1102),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_980),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1028),
.B(n_908),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_976),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_973),
.A2(n_1008),
.B(n_972),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_969),
.B(n_1093),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_968),
.B(n_1102),
.Y(n_1233)
);

OR2x6_ASAP7_75t_L g1234 ( 
.A(n_995),
.B(n_661),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1041),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1016),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_969),
.A2(n_935),
.B1(n_926),
.B2(n_928),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_980),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1041),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_968),
.B(n_1102),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_969),
.A2(n_944),
.B(n_959),
.C(n_940),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1041),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_968),
.B(n_1102),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1028),
.B(n_908),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_983),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1041),
.Y(n_1246)
);

AOI21xp33_ASAP7_75t_SL g1247 ( 
.A1(n_996),
.A2(n_467),
.B(n_455),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_968),
.B(n_1102),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_980),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1016),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_1107),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_969),
.A2(n_852),
.B1(n_1095),
.B2(n_1093),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_980),
.Y(n_1253)
);

AO22x1_ASAP7_75t_L g1254 ( 
.A1(n_969),
.A2(n_852),
.B1(n_1095),
.B2(n_1093),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1228),
.Y(n_1255)
);

NAND2x1p5_ASAP7_75t_L g1256 ( 
.A(n_1119),
.B(n_1129),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1110),
.B(n_1135),
.Y(n_1257)
);

AO21x1_ASAP7_75t_L g1258 ( 
.A1(n_1241),
.A2(n_1140),
.B(n_1130),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1135),
.B(n_1137),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1143),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1236),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1252),
.A2(n_1214),
.B1(n_1212),
.B2(n_1232),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1136),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1251),
.Y(n_1264)
);

OAI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1212),
.A2(n_1232),
.B1(n_1109),
.B2(n_1237),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1254),
.B(n_1137),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1113),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1250),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1237),
.B(n_1221),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1253),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1119),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1185),
.A2(n_1140),
.B1(n_1112),
.B2(n_1131),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1227),
.A2(n_1240),
.B1(n_1233),
.B2(n_1248),
.Y(n_1273)
);

BUFx2_ASAP7_75t_R g1274 ( 
.A(n_1178),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1121),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_1111),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1243),
.B(n_1149),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1136),
.Y(n_1278)
);

CKINVDCx9p33_ASAP7_75t_R g1279 ( 
.A(n_1149),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1119),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1216),
.A2(n_1218),
.B1(n_1220),
.B2(n_1231),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1164),
.Y(n_1282)
);

CKINVDCx11_ASAP7_75t_R g1283 ( 
.A(n_1159),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1129),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1124),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1158),
.A2(n_1216),
.B1(n_1218),
.B2(n_1220),
.Y(n_1286)
);

BUFx4f_ASAP7_75t_SL g1287 ( 
.A(n_1111),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1226),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1114),
.A2(n_1130),
.B1(n_1141),
.B2(n_1152),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1155),
.Y(n_1290)
);

NOR2x1_ASAP7_75t_R g1291 ( 
.A(n_1245),
.B(n_1222),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1223),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1231),
.A2(n_1172),
.B1(n_1151),
.B2(n_1152),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1182),
.B(n_1176),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1114),
.A2(n_1133),
.B1(n_1148),
.B2(n_1246),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1181),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1195),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_1217),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1224),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1196),
.A2(n_1157),
.B(n_1174),
.Y(n_1300)
);

INVxp33_ASAP7_75t_L g1301 ( 
.A(n_1165),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1196),
.A2(n_1166),
.B(n_1150),
.Y(n_1302)
);

BUFx4f_ASAP7_75t_SL g1303 ( 
.A(n_1217),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1187),
.B(n_1175),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1235),
.A2(n_1206),
.B1(n_1247),
.B2(n_1127),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1125),
.A2(n_1242),
.B1(n_1239),
.B2(n_1151),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1238),
.Y(n_1307)
);

INVx6_ASAP7_75t_L g1308 ( 
.A(n_1190),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1127),
.A2(n_1117),
.B1(n_1162),
.B2(n_1241),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1249),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1156),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1123),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1145),
.B(n_1116),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1222),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1117),
.Y(n_1315)
);

BUFx8_ASAP7_75t_L g1316 ( 
.A(n_1229),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1195),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1179),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1195),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1122),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1229),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1170),
.A2(n_1150),
.B(n_1118),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1126),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1116),
.A2(n_1120),
.B1(n_1134),
.B2(n_1145),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1207),
.B(n_1201),
.Y(n_1325)
);

BUFx2_ASAP7_75t_SL g1326 ( 
.A(n_1173),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1139),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1120),
.B(n_1134),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1197),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1208),
.Y(n_1330)
);

NAND2x1p5_ASAP7_75t_L g1331 ( 
.A(n_1207),
.B(n_1201),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1191),
.A2(n_1180),
.B1(n_1138),
.B2(n_1146),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1177),
.B(n_1184),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1193),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1192),
.B(n_1118),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_1199),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1198),
.A2(n_1142),
.B1(n_1234),
.B2(n_1186),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1188),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1189),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1192),
.B(n_1194),
.Y(n_1340)
);

OA21x2_ASAP7_75t_L g1341 ( 
.A1(n_1154),
.A2(n_1202),
.B(n_1163),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1194),
.A2(n_1244),
.B1(n_1234),
.B2(n_1167),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1234),
.A2(n_1161),
.B1(n_1132),
.B2(n_1183),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1144),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_1169),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1144),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1244),
.Y(n_1347)
);

AOI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1202),
.A2(n_1204),
.B(n_1200),
.Y(n_1348)
);

BUFx12f_ASAP7_75t_L g1349 ( 
.A(n_1160),
.Y(n_1349)
);

AO21x1_ASAP7_75t_SL g1350 ( 
.A1(n_1128),
.A2(n_1205),
.B(n_1200),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1171),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1128),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1171),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1128),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1211),
.A2(n_1183),
.B1(n_1168),
.B2(n_1132),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1210),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1147),
.A2(n_1115),
.B1(n_1213),
.B2(n_1230),
.Y(n_1357)
);

CKINVDCx11_ASAP7_75t_R g1358 ( 
.A(n_1160),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1160),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1203),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1183),
.A2(n_1161),
.B1(n_1132),
.B2(n_1153),
.Y(n_1361)
);

AO21x1_ASAP7_75t_L g1362 ( 
.A1(n_1219),
.A2(n_1209),
.B(n_1161),
.Y(n_1362)
);

AO21x2_ASAP7_75t_L g1363 ( 
.A1(n_1153),
.A2(n_1213),
.B(n_1230),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1215),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1215),
.Y(n_1365)
);

INVx3_ASAP7_75t_SL g1366 ( 
.A(n_1225),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1225),
.Y(n_1367)
);

NOR2x1_ASAP7_75t_R g1368 ( 
.A(n_1178),
.B(n_769),
.Y(n_1368)
);

BUFx10_ASAP7_75t_L g1369 ( 
.A(n_1164),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1251),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1214),
.A2(n_1093),
.B1(n_1095),
.B2(n_969),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1335),
.B(n_1333),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1335),
.B(n_1333),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1348),
.A2(n_1302),
.B(n_1300),
.Y(n_1374)
);

INVxp67_ASAP7_75t_SL g1375 ( 
.A(n_1281),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1282),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1356),
.B(n_1328),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1356),
.B(n_1328),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1340),
.B(n_1304),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1325),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1340),
.B(n_1304),
.Y(n_1381)
);

BUFx4f_ASAP7_75t_SL g1382 ( 
.A(n_1370),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1322),
.B(n_1352),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1341),
.A2(n_1289),
.B(n_1258),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1325),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1325),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1352),
.B(n_1354),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1354),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1259),
.B(n_1257),
.Y(n_1389)
);

AO31x2_ASAP7_75t_L g1390 ( 
.A1(n_1258),
.A2(n_1309),
.A3(n_1313),
.B(n_1362),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1331),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1257),
.B(n_1259),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1318),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1350),
.B(n_1286),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1265),
.A2(n_1266),
.B(n_1306),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1371),
.B(n_1262),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1275),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1292),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1299),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1271),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1307),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1310),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1324),
.A2(n_1362),
.B(n_1343),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1312),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1350),
.B(n_1293),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1318),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1295),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1269),
.B(n_1294),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1256),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1272),
.A2(n_1256),
.B(n_1360),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1255),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1270),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1337),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1320),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1361),
.A2(n_1355),
.B(n_1284),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1363),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1290),
.B(n_1301),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1323),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1363),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1327),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1277),
.B(n_1342),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1278),
.B(n_1330),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1261),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1338),
.B(n_1339),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1271),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1271),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1271),
.B(n_1280),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1268),
.Y(n_1428)
);

AO21x2_ASAP7_75t_L g1429 ( 
.A1(n_1344),
.A2(n_1359),
.B(n_1365),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1357),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1416),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1417),
.B(n_1268),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1417),
.B(n_1263),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1372),
.B(n_1273),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1372),
.B(n_1288),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1372),
.B(n_1288),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1373),
.B(n_1267),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1373),
.B(n_1267),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1417),
.B(n_1315),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1392),
.B(n_1285),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1380),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1396),
.A2(n_1305),
.B1(n_1334),
.B2(n_1326),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1429),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1373),
.B(n_1351),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1396),
.A2(n_1332),
.B(n_1329),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1392),
.B(n_1389),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1392),
.B(n_1285),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1379),
.B(n_1381),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1380),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1388),
.B(n_1330),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1389),
.B(n_1330),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1408),
.B(n_1351),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1393),
.Y(n_1453)
);

INVx4_ASAP7_75t_L g1454 ( 
.A(n_1427),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1380),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1379),
.B(n_1351),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1379),
.B(n_1353),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1416),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1423),
.Y(n_1459)
);

OAI33xp33_ASAP7_75t_L g1460 ( 
.A1(n_1422),
.A2(n_1346),
.A3(n_1311),
.B1(n_1334),
.B2(n_1260),
.B3(n_1264),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1393),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1413),
.A2(n_1298),
.B1(n_1326),
.B2(n_1314),
.Y(n_1462)
);

NOR2x1_ASAP7_75t_L g1463 ( 
.A(n_1395),
.B(n_1296),
.Y(n_1463)
);

NAND2x1p5_ASAP7_75t_L g1464 ( 
.A(n_1410),
.B(n_1280),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1377),
.B(n_1378),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1408),
.B(n_1264),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1381),
.B(n_1345),
.Y(n_1467)
);

INVxp67_ASAP7_75t_L g1468 ( 
.A(n_1423),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1408),
.B(n_1364),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1428),
.Y(n_1470)
);

OAI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1375),
.A2(n_1296),
.B1(n_1260),
.B2(n_1308),
.C(n_1321),
.Y(n_1471)
);

INVx2_ASAP7_75t_SL g1472 ( 
.A(n_1429),
.Y(n_1472)
);

INVxp67_ASAP7_75t_SL g1473 ( 
.A(n_1428),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1381),
.B(n_1377),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1429),
.Y(n_1475)
);

OAI221xp5_ASAP7_75t_L g1476 ( 
.A1(n_1375),
.A2(n_1308),
.B1(n_1347),
.B2(n_1314),
.C(n_1321),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1380),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1377),
.B(n_1345),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1386),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1383),
.B(n_1367),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1377),
.B(n_1364),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1406),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1377),
.B(n_1280),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1422),
.B(n_1346),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1432),
.B(n_1406),
.Y(n_1485)
);

NAND4xp25_ASAP7_75t_L g1486 ( 
.A(n_1445),
.B(n_1421),
.C(n_1413),
.D(n_1406),
.Y(n_1486)
);

OA211x2_ASAP7_75t_L g1487 ( 
.A1(n_1462),
.A2(n_1421),
.B(n_1279),
.C(n_1395),
.Y(n_1487)
);

NOR3xp33_ASAP7_75t_L g1488 ( 
.A(n_1460),
.B(n_1407),
.C(n_1430),
.Y(n_1488)
);

OAI21xp33_ASAP7_75t_L g1489 ( 
.A1(n_1442),
.A2(n_1407),
.B(n_1394),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1474),
.B(n_1387),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1439),
.B(n_1395),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1443),
.A2(n_1374),
.B(n_1384),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1474),
.B(n_1448),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1448),
.B(n_1387),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1433),
.B(n_1395),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1442),
.A2(n_1430),
.B1(n_1382),
.B2(n_1308),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1446),
.B(n_1395),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1465),
.B(n_1387),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1465),
.B(n_1378),
.Y(n_1499)
);

NAND3xp33_ASAP7_75t_L g1500 ( 
.A(n_1463),
.B(n_1412),
.C(n_1411),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1451),
.B(n_1401),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1465),
.B(n_1378),
.Y(n_1502)
);

NOR3xp33_ASAP7_75t_L g1503 ( 
.A(n_1471),
.B(n_1415),
.C(n_1425),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1435),
.B(n_1401),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_L g1505 ( 
.A(n_1463),
.B(n_1411),
.C(n_1412),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1476),
.A2(n_1394),
.B(n_1405),
.Y(n_1506)
);

NAND4xp25_ASAP7_75t_L g1507 ( 
.A(n_1466),
.B(n_1404),
.C(n_1399),
.D(n_1398),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1465),
.B(n_1378),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1435),
.B(n_1402),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1436),
.B(n_1402),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1436),
.B(n_1459),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1437),
.B(n_1394),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1484),
.A2(n_1415),
.B(n_1410),
.Y(n_1513)
);

OAI221xp5_ASAP7_75t_SL g1514 ( 
.A1(n_1434),
.A2(n_1405),
.B1(n_1440),
.B2(n_1447),
.C(n_1468),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1469),
.B(n_1402),
.Y(n_1515)
);

OAI211xp5_ASAP7_75t_SL g1516 ( 
.A1(n_1470),
.A2(n_1404),
.B(n_1399),
.C(n_1398),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1437),
.B(n_1402),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1438),
.B(n_1416),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1438),
.B(n_1397),
.Y(n_1519)
);

NAND3xp33_ASAP7_75t_L g1520 ( 
.A(n_1453),
.B(n_1386),
.C(n_1391),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1444),
.B(n_1416),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1452),
.A2(n_1382),
.B1(n_1308),
.B2(n_1336),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1461),
.B(n_1397),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1434),
.B(n_1397),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1473),
.B(n_1420),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1444),
.B(n_1416),
.Y(n_1526)
);

AOI211xp5_ASAP7_75t_L g1527 ( 
.A1(n_1450),
.A2(n_1405),
.B(n_1291),
.C(n_1403),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1467),
.B(n_1419),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1443),
.B(n_1414),
.C(n_1418),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1467),
.B(n_1419),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1483),
.B(n_1376),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1483),
.B(n_1385),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1456),
.B(n_1420),
.Y(n_1533)
);

OAI21xp33_ASAP7_75t_L g1534 ( 
.A1(n_1450),
.A2(n_1384),
.B(n_1424),
.Y(n_1534)
);

OAI22x1_ASAP7_75t_SL g1535 ( 
.A1(n_1454),
.A2(n_1276),
.B1(n_1370),
.B2(n_1282),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_R g1536 ( 
.A(n_1481),
.B(n_1276),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1498),
.B(n_1472),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1525),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1523),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1528),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1528),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1497),
.B(n_1390),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1521),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1530),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1495),
.B(n_1482),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1521),
.Y(n_1546)
);

NAND2x1p5_ASAP7_75t_L g1547 ( 
.A(n_1492),
.B(n_1454),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1498),
.B(n_1472),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1526),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1491),
.B(n_1390),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1493),
.B(n_1475),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1529),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1515),
.B(n_1390),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1526),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1533),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1485),
.B(n_1480),
.Y(n_1556)
);

NOR2x1_ASAP7_75t_L g1557 ( 
.A(n_1500),
.B(n_1454),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1494),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1493),
.B(n_1475),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1490),
.B(n_1454),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1494),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1499),
.B(n_1431),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1499),
.B(n_1431),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1529),
.Y(n_1564)
);

INVxp67_ASAP7_75t_SL g1565 ( 
.A(n_1500),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1504),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1502),
.B(n_1431),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1502),
.B(n_1458),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1509),
.B(n_1510),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1524),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1517),
.B(n_1480),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1492),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1518),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1501),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1492),
.Y(n_1575)
);

INVx4_ASAP7_75t_L g1576 ( 
.A(n_1492),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1508),
.B(n_1518),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1519),
.B(n_1479),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1560),
.B(n_1512),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1560),
.B(n_1567),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1538),
.B(n_1512),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1538),
.B(n_1511),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1558),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1558),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1545),
.B(n_1534),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1557),
.Y(n_1586)
);

INVxp67_ASAP7_75t_L g1587 ( 
.A(n_1556),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1545),
.B(n_1534),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1570),
.B(n_1456),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1553),
.B(n_1505),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1570),
.B(n_1457),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1561),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1557),
.B(n_1536),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1560),
.B(n_1513),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1553),
.B(n_1505),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1567),
.B(n_1527),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1567),
.B(n_1527),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1539),
.B(n_1457),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1556),
.B(n_1298),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1540),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1539),
.B(n_1507),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1574),
.B(n_1489),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1561),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1541),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1574),
.B(n_1489),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1555),
.B(n_1488),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1555),
.B(n_1503),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1541),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1544),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1567),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1550),
.B(n_1496),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1544),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1564),
.B(n_1542),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1567),
.B(n_1532),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1547),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1552),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1571),
.B(n_1303),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1606),
.B(n_1566),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1583),
.Y(n_1619)
);

A2O1A1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1593),
.A2(n_1565),
.B(n_1552),
.C(n_1506),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1600),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1600),
.Y(n_1622)
);

OAI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1611),
.A2(n_1565),
.B(n_1564),
.Y(n_1623)
);

AO21x1_ASAP7_75t_L g1624 ( 
.A1(n_1616),
.A2(n_1576),
.B(n_1550),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1583),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1584),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1596),
.B(n_1568),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1601),
.B(n_1602),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1605),
.B(n_1566),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1607),
.B(n_1542),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1587),
.B(n_1616),
.Y(n_1631)
);

O2A1O1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1586),
.A2(n_1486),
.B(n_1522),
.C(n_1514),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1584),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1596),
.B(n_1568),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1592),
.Y(n_1635)
);

NOR2x1p5_ASAP7_75t_L g1636 ( 
.A(n_1597),
.B(n_1535),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1592),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1582),
.B(n_1537),
.Y(n_1638)
);

NOR3xp33_ASAP7_75t_L g1639 ( 
.A(n_1599),
.B(n_1520),
.C(n_1516),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1617),
.B(n_1287),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1613),
.B(n_1578),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1603),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1604),
.Y(n_1643)
);

AOI32xp33_ASAP7_75t_L g1644 ( 
.A1(n_1597),
.A2(n_1551),
.A3(n_1559),
.B1(n_1548),
.B2(n_1537),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1581),
.B(n_1537),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1604),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1610),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1613),
.B(n_1548),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1594),
.A2(n_1487),
.B1(n_1531),
.B2(n_1483),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1608),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1615),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1580),
.B(n_1568),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1580),
.B(n_1568),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1586),
.Y(n_1654)
);

AOI21xp33_ASAP7_75t_L g1655 ( 
.A1(n_1590),
.A2(n_1571),
.B(n_1578),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1614),
.B(n_1568),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1585),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1614),
.B(n_1577),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1608),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1594),
.B(n_1577),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1623),
.A2(n_1535),
.B(n_1590),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1657),
.B(n_1595),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1628),
.B(n_1283),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1618),
.B(n_1579),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1627),
.B(n_1610),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1640),
.B(n_1283),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1639),
.B(n_1579),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1630),
.B(n_1620),
.Y(n_1668)
);

BUFx2_ASAP7_75t_L g1669 ( 
.A(n_1654),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1654),
.B(n_1615),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1631),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1619),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1658),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1627),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1636),
.B(n_1595),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1647),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1619),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1629),
.B(n_1632),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1658),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1625),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1625),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1634),
.B(n_1615),
.Y(n_1682)
);

NOR2xp67_ASAP7_75t_SL g1683 ( 
.A(n_1647),
.B(n_1311),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1621),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1634),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1621),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1655),
.B(n_1369),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1649),
.A2(n_1487),
.B1(n_1585),
.B2(n_1588),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1622),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1626),
.Y(n_1690)
);

OAI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1644),
.A2(n_1588),
.B1(n_1547),
.B2(n_1598),
.C(n_1591),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1638),
.B(n_1369),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1624),
.A2(n_1483),
.B1(n_1478),
.B2(n_1612),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1660),
.B(n_1577),
.Y(n_1694)
);

INVx3_ASAP7_75t_SL g1695 ( 
.A(n_1641),
.Y(n_1695)
);

CKINVDCx16_ASAP7_75t_R g1696 ( 
.A(n_1660),
.Y(n_1696)
);

OAI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1678),
.A2(n_1641),
.B1(n_1648),
.B2(n_1642),
.C(n_1651),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1672),
.Y(n_1698)
);

NAND2x1_ASAP7_75t_L g1699 ( 
.A(n_1683),
.B(n_1651),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1695),
.B(n_1642),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1672),
.Y(n_1701)
);

NOR2x1_ASAP7_75t_SL g1702 ( 
.A(n_1662),
.B(n_1652),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1676),
.Y(n_1703)
);

OAI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1661),
.A2(n_1651),
.B1(n_1645),
.B2(n_1626),
.C(n_1643),
.Y(n_1704)
);

OAI21xp33_ASAP7_75t_L g1705 ( 
.A1(n_1668),
.A2(n_1635),
.B(n_1633),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1669),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1677),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1695),
.B(n_1656),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1677),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1680),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1663),
.B(n_1369),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1695),
.B(n_1669),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1688),
.A2(n_1696),
.B1(n_1667),
.B2(n_1675),
.Y(n_1713)
);

AOI221xp5_ASAP7_75t_L g1714 ( 
.A1(n_1671),
.A2(n_1624),
.B1(n_1633),
.B2(n_1659),
.C(n_1635),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1696),
.A2(n_1656),
.B1(n_1653),
.B2(n_1652),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1674),
.B(n_1653),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1687),
.A2(n_1659),
.B1(n_1650),
.B2(n_1646),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1683),
.Y(n_1718)
);

NAND2xp33_ASAP7_75t_SL g1719 ( 
.A(n_1662),
.B(n_1336),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1680),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_SL g1721 ( 
.A(n_1685),
.B(n_1547),
.C(n_1637),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1692),
.B(n_1637),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1706),
.B(n_1712),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1713),
.A2(n_1691),
.B1(n_1679),
.B2(n_1673),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1703),
.B(n_1705),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1708),
.B(n_1673),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_SL g1727 ( 
.A(n_1718),
.B(n_1274),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1711),
.B(n_1666),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1719),
.B(n_1664),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1699),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1702),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1700),
.B(n_1679),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1715),
.B(n_1676),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1698),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1722),
.B(n_1665),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1701),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1707),
.Y(n_1737)
);

INVxp67_ASAP7_75t_L g1738 ( 
.A(n_1697),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1709),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1717),
.B(n_1665),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1716),
.B(n_1670),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1710),
.Y(n_1742)
);

OAI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1738),
.A2(n_1704),
.B1(n_1714),
.B2(n_1697),
.C(n_1693),
.Y(n_1743)
);

OAI32xp33_ASAP7_75t_L g1744 ( 
.A1(n_1731),
.A2(n_1704),
.A3(n_1720),
.B1(n_1690),
.B2(n_1681),
.Y(n_1744)
);

OAI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1724),
.A2(n_1721),
.B1(n_1690),
.B2(n_1681),
.C(n_1694),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1741),
.B(n_1729),
.Y(n_1746)
);

OAI222xp33_ASAP7_75t_L g1747 ( 
.A1(n_1731),
.A2(n_1670),
.B1(n_1682),
.B2(n_1684),
.C1(n_1686),
.C2(n_1689),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1733),
.A2(n_1682),
.B1(n_1670),
.B2(n_1689),
.Y(n_1748)
);

OAI21xp33_ASAP7_75t_L g1749 ( 
.A1(n_1733),
.A2(n_1740),
.B(n_1741),
.Y(n_1749)
);

AOI322xp5_ASAP7_75t_L g1750 ( 
.A1(n_1725),
.A2(n_1682),
.A3(n_1670),
.B1(n_1686),
.B2(n_1684),
.C1(n_1650),
.C2(n_1646),
.Y(n_1750)
);

NOR4xp25_ASAP7_75t_L g1751 ( 
.A(n_1723),
.B(n_1643),
.C(n_1622),
.D(n_1612),
.Y(n_1751)
);

AOI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1727),
.A2(n_1682),
.B1(n_1609),
.B2(n_1547),
.Y(n_1752)
);

AO21x1_ASAP7_75t_L g1753 ( 
.A1(n_1734),
.A2(n_1576),
.B(n_1609),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1723),
.B(n_1548),
.Y(n_1754)
);

NOR3xp33_ASAP7_75t_L g1755 ( 
.A(n_1749),
.B(n_1732),
.C(n_1728),
.Y(n_1755)
);

NAND3xp33_ASAP7_75t_L g1756 ( 
.A(n_1743),
.B(n_1726),
.C(n_1736),
.Y(n_1756)
);

XNOR2x1_ASAP7_75t_L g1757 ( 
.A(n_1746),
.B(n_1730),
.Y(n_1757)
);

NOR3xp33_ASAP7_75t_L g1758 ( 
.A(n_1744),
.B(n_1735),
.C(n_1737),
.Y(n_1758)
);

NOR2x1_ASAP7_75t_SL g1759 ( 
.A(n_1754),
.B(n_1742),
.Y(n_1759)
);

OAI211xp5_ASAP7_75t_SL g1760 ( 
.A1(n_1750),
.A2(n_1745),
.B(n_1748),
.C(n_1752),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1751),
.B(n_1742),
.Y(n_1761)
);

NOR2x1_ASAP7_75t_L g1762 ( 
.A(n_1747),
.B(n_1734),
.Y(n_1762)
);

NAND2x1_ASAP7_75t_SL g1763 ( 
.A(n_1753),
.B(n_1739),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1746),
.B(n_1739),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_SL g1765 ( 
.A1(n_1743),
.A2(n_1576),
.B1(n_1477),
.B2(n_1441),
.Y(n_1765)
);

AOI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1743),
.A2(n_1368),
.B(n_1366),
.C(n_1572),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1759),
.B(n_1562),
.Y(n_1767)
);

OAI221xp5_ASAP7_75t_SL g1768 ( 
.A1(n_1758),
.A2(n_1427),
.B1(n_1575),
.B2(n_1572),
.C(n_1589),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1762),
.A2(n_1576),
.B(n_1429),
.Y(n_1769)
);

AOI221xp5_ASAP7_75t_L g1770 ( 
.A1(n_1760),
.A2(n_1575),
.B1(n_1572),
.B2(n_1551),
.C(n_1559),
.Y(n_1770)
);

INVxp67_ASAP7_75t_SL g1771 ( 
.A(n_1763),
.Y(n_1771)
);

NOR3x1_ASAP7_75t_L g1772 ( 
.A(n_1756),
.B(n_1455),
.C(n_1449),
.Y(n_1772)
);

OAI221xp5_ASAP7_75t_L g1773 ( 
.A1(n_1755),
.A2(n_1575),
.B1(n_1464),
.B2(n_1543),
.C(n_1409),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1767),
.B(n_1757),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1771),
.Y(n_1775)
);

NOR2xp67_ASAP7_75t_L g1776 ( 
.A(n_1769),
.B(n_1761),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1772),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1770),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1768),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1773),
.A2(n_1765),
.B1(n_1764),
.B2(n_1766),
.Y(n_1780)
);

NAND5xp2_ASAP7_75t_L g1781 ( 
.A(n_1780),
.B(n_1358),
.C(n_1464),
.D(n_1551),
.E(n_1559),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1774),
.A2(n_1358),
.B1(n_1429),
.B2(n_1349),
.Y(n_1782)
);

NOR2xp67_ASAP7_75t_L g1783 ( 
.A(n_1775),
.B(n_1349),
.Y(n_1783)
);

INVxp33_ASAP7_75t_L g1784 ( 
.A(n_1779),
.Y(n_1784)
);

AOI31xp33_ASAP7_75t_L g1785 ( 
.A1(n_1777),
.A2(n_1400),
.A3(n_1464),
.B(n_1366),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1784),
.Y(n_1786)
);

NOR3xp33_ASAP7_75t_L g1787 ( 
.A(n_1783),
.B(n_1776),
.C(n_1778),
.Y(n_1787)
);

INVxp33_ASAP7_75t_SL g1788 ( 
.A(n_1782),
.Y(n_1788)
);

AOI22x1_ASAP7_75t_L g1789 ( 
.A1(n_1786),
.A2(n_1785),
.B1(n_1781),
.B2(n_1280),
.Y(n_1789)
);

OR3x1_ASAP7_75t_L g1790 ( 
.A(n_1789),
.B(n_1788),
.C(n_1787),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1790),
.A2(n_1554),
.B1(n_1546),
.B2(n_1549),
.C(n_1543),
.Y(n_1791)
);

AOI21x1_ASAP7_75t_L g1792 ( 
.A1(n_1790),
.A2(n_1563),
.B(n_1562),
.Y(n_1792)
);

NOR3xp33_ASAP7_75t_L g1793 ( 
.A(n_1792),
.B(n_1426),
.C(n_1425),
.Y(n_1793)
);

INVxp67_ASAP7_75t_SL g1794 ( 
.A(n_1791),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1794),
.A2(n_1418),
.B(n_1414),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1793),
.A2(n_1569),
.B(n_1549),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1795),
.B(n_1543),
.Y(n_1797)
);

AOI222xp33_ASAP7_75t_L g1798 ( 
.A1(n_1797),
.A2(n_1796),
.B1(n_1297),
.B2(n_1317),
.C1(n_1319),
.C2(n_1316),
.Y(n_1798)
);

OAI221xp5_ASAP7_75t_R g1799 ( 
.A1(n_1798),
.A2(n_1543),
.B1(n_1316),
.B2(n_1573),
.C(n_1569),
.Y(n_1799)
);

AOI211xp5_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1297),
.B(n_1317),
.C(n_1319),
.Y(n_1800)
);


endmodule