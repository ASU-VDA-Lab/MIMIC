module real_jpeg_17003_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_0),
.B(n_28),
.Y(n_27)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_0),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_0),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_0),
.B(n_146),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_0),
.B(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_1),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_2),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_2),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_2),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_2),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_2),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_2),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_2),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_2),
.B(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_3),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_3),
.Y(n_236)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_3),
.Y(n_350)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_4),
.Y(n_102)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_4),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_4),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_4),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_33),
.Y(n_32)
);

NAND2x1_ASAP7_75t_SL g73 ( 
.A(n_5),
.B(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_5),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_5),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_5),
.B(n_50),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g227 ( 
.A(n_5),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_5),
.B(n_257),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_6),
.Y(n_187)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_6),
.Y(n_231)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_7),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_7),
.Y(n_329)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_7),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_8),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_8),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_8),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_8),
.B(n_48),
.Y(n_188)
);

NAND2x1_ASAP7_75t_L g189 ( 
.A(n_8),
.B(n_190),
.Y(n_189)
);

AOI22x1_ASAP7_75t_SL g268 ( 
.A1(n_8),
.A2(n_12),
.B1(n_254),
.B2(n_269),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_8),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_9),
.B(n_78),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_9),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_9),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_9),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_9),
.B(n_74),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_9),
.B(n_50),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_9),
.B(n_52),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_10),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_10),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_10),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_10),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_10),
.B(n_392),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_10),
.Y(n_403)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_11),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_11),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_12),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_12),
.B(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_12),
.B(n_235),
.Y(n_234)
);

AOI31xp33_ASAP7_75t_L g291 ( 
.A1(n_12),
.A2(n_268),
.A3(n_292),
.B(n_295),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_12),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_12),
.B(n_190),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_12),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_12),
.B(n_52),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_13),
.B(n_33),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_13),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_13),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_13),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_13),
.B(n_174),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g222 ( 
.A(n_13),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_13),
.B(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_13),
.B(n_186),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_14),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_14),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_15),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_15),
.B(n_75),
.Y(n_96)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

BUFx8_ASAP7_75t_L g142 ( 
.A(n_16),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_204),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_202),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_157),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_22),
.B(n_157),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_92),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_68),
.C(n_85),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_25),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_42),
.C(n_54),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_26),
.B(n_42),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_27),
.B(n_37),
.C(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_30),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_37),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_32),
.Y(n_133)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_36),
.Y(n_149)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.C(n_51),
.Y(n_42)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_43),
.B(n_166),
.Y(n_165)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_47),
.A2(n_51),
.B1(n_66),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_47),
.Y(n_167)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_50),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_51),
.Y(n_66)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_56),
.C(n_62),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_53),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_54),
.B(n_454),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_55),
.A2(n_56),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_55),
.B(n_214),
.C(n_218),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_62),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_62),
.A2(n_67),
.B1(n_97),
.B2(n_98),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_65),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_98),
.C(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_68),
.B(n_85),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_77),
.C(n_80),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_69),
.B(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.C(n_76),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_70),
.B(n_76),
.Y(n_182)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

XOR2x1_ASAP7_75t_L g181 ( 
.A(n_73),
.B(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_77),
.A2(n_80),
.B1(n_81),
.B2(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_77),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_79),
.Y(n_249)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_87),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_81),
.B(n_90),
.C(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_84),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_88),
.B(n_185),
.C(n_188),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_89),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_128),
.B1(n_155),
.B2(n_156),
.Y(n_92)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

XNOR2x2_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_108),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_103),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_110),
.B(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.C(n_123),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_136),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_134),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_134),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_138),
.B(n_266),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_150),
.B2(n_154),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_163),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_158),
.B(n_160),
.Y(n_463)
);

XNOR2x1_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_163),
.B(n_463),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_183),
.C(n_198),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_164),
.B(n_452),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_181),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_165),
.B(n_168),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.C(n_178),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_169),
.A2(n_178),
.B1(n_179),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_169),
.Y(n_261)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_173),
.B(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_178),
.B(n_322),
.C(n_326),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_178),
.A2(n_179),
.B1(n_322),
.B2(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_181),
.B(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_183),
.B(n_199),
.Y(n_452)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.C(n_192),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_184),
.B(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_185),
.B(n_188),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_189),
.B(n_193),
.Y(n_275)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_192),
.A2(n_193),
.B1(n_303),
.B2(n_304),
.Y(n_429)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_193),
.B(n_300),
.C(n_303),
.Y(n_299)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_196),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g325 ( 
.A(n_197),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AO21x2_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_443),
.B(n_467),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_336),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_282),
.C(n_310),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_209),
.B(n_283),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_262),
.Y(n_209)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_210),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_245),
.C(n_259),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_211),
.B(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_220),
.C(n_232),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_SL g332 ( 
.A(n_213),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_218),
.Y(n_219)
);

XNOR2x1_ASAP7_75t_L g333 ( 
.A(n_220),
.B(n_233),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_227),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_221),
.B(n_227),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_230),
.Y(n_298)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_241),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_234),
.A2(n_237),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_234),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_237),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_237),
.A2(n_319),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_237),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_240),
.Y(n_381)
);

XOR2x2_ASAP7_75t_SL g316 ( 
.A(n_241),
.B(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_259),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_252),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_253),
.C(n_273),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.C(n_250),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_247),
.A2(n_250),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

XNOR2x2_ASAP7_75t_SL g344 ( 
.A(n_247),
.B(n_345),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_288),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_250),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_258),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_262)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_271),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_264),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.C(n_270),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_308),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_270),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_271)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_272),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_272),
.Y(n_448)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_274),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_277),
.Y(n_449)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_278),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_280),
.Y(n_458)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.C(n_307),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_284),
.B(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_286),
.B(n_307),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.C(n_299),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_291),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_289),
.B(n_346),
.C(n_351),
.Y(n_369)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx2_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_300),
.B(n_429),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

XNOR2x1_ASAP7_75t_SL g376 ( 
.A(n_301),
.B(n_302),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_301),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_301),
.A2(n_397),
.B1(n_398),
.B2(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_334),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_334),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.C(n_332),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_312),
.B(n_441),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_315),
.B(n_332),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.C(n_330),
.Y(n_315)
);

XOR2x1_ASAP7_75t_L g433 ( 
.A(n_316),
.B(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_321),
.B(n_331),
.Y(n_434)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_322),
.Y(n_372)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XOR2x2_ASAP7_75t_L g370 ( 
.A(n_326),
.B(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND3xp33_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_338),
.C(n_339),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_340),
.A2(n_437),
.B(n_442),
.Y(n_339)
);

AOI21x1_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_423),
.B(n_436),
.Y(n_340)
);

OAI21x1_ASAP7_75t_SL g341 ( 
.A1(n_342),
.A2(n_382),
.B(n_422),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_367),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_343),
.B(n_367),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_352),
.C(n_360),
.Y(n_343)
);

XOR2x1_ASAP7_75t_L g416 ( 
.A(n_344),
.B(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_351),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_352),
.A2(n_353),
.B1(n_360),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_354),
.B(n_357),
.Y(n_387)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_360),
.Y(n_418)
);

AO22x1_ASAP7_75t_SL g360 ( 
.A1(n_361),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.Y(n_360)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_361),
.Y(n_365)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_364),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_365),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_407),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_373),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_369),
.B(n_370),
.C(n_373),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g431 ( 
.A(n_374),
.B(n_376),
.C(n_377),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

AOI21x1_ASAP7_75t_SL g382 ( 
.A1(n_383),
.A2(n_415),
.B(n_421),
.Y(n_382)
);

OAI21x1_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_399),
.B(n_414),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_396),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_396),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_386),
.B(n_390),
.C(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_398),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_406),
.B(n_413),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_404),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_403),
.B(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_419),
.Y(n_415)
);

NOR2xp67_ASAP7_75t_SL g421 ( 
.A(n_416),
.B(n_419),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_435),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_424),
.B(n_435),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_432),
.B2(n_433),
.Y(n_424)
);

INVxp33_ASAP7_75t_SL g425 ( 
.A(n_426),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_428),
.B1(n_430),
.B2(n_431),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_427),
.Y(n_439)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_432),
.C(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_440),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_440),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_461),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_457),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_457),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_450),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_446),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.C(n_449),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_451),
.A2(n_453),
.B1(n_455),
.B2(n_456),
.Y(n_450)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_451),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_453),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_453),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_455),
.B(n_465),
.C(n_466),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.C(n_460),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_461),
.A2(n_468),
.B(n_469),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_464),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_462),
.B(n_464),
.Y(n_469)
);


endmodule