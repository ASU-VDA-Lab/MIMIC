module fake_jpeg_644_n_194 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_194);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_29),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_0),
.Y(n_63)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_74),
.Y(n_84)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_78),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_3),
.Y(n_78)
);

AND2x4_ASAP7_75t_SL g80 ( 
.A(n_73),
.B(n_57),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_77),
.B(n_71),
.C(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_89),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_73),
.B(n_74),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_77),
.B(n_71),
.C(n_61),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_103),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_80),
.B1(n_73),
.B2(n_67),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_60),
.B1(n_58),
.B2(n_65),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_50),
.Y(n_131)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_69),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_56),
.Y(n_107)
);

XNOR2x1_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_80),
.B(n_56),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_34),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_26),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_61),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_115),
.B1(n_118),
.B2(n_129),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_71),
.B1(n_79),
.B2(n_67),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_131),
.B1(n_45),
.B2(n_43),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_55),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_119),
.C(n_65),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_68),
.B1(n_52),
.B2(n_54),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_63),
.C(n_68),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_24),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_119),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_63),
.B1(n_54),
.B2(n_60),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_108),
.B1(n_96),
.B2(n_110),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_93),
.A2(n_50),
.B1(n_60),
.B2(n_64),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_3),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_4),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_121),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_134),
.C(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_140),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_64),
.B1(n_58),
.B2(n_70),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_131),
.B1(n_114),
.B2(n_13),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_70),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_139),
.C(n_143),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_48),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_4),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_37),
.Y(n_157)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_116),
.B(n_47),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_6),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_147),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_7),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_8),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_149),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_8),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_42),
.C(n_40),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_152),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_9),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_154),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_9),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_157),
.B1(n_145),
.B2(n_150),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_151),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_164),
.B1(n_15),
.B2(n_16),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_151),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_39),
.B(n_36),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C1(n_18),
.C2(n_19),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_25),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_173),
.B1(n_175),
.B2(n_165),
.Y(n_179)
);

NAND2xp67_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_137),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_172),
.A2(n_170),
.B(n_160),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_168),
.A2(n_139),
.B1(n_134),
.B2(n_20),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_178),
.C(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_28),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_166),
.A3(n_168),
.B1(n_157),
.B2(n_159),
.C1(n_161),
.C2(n_164),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_184),
.B(n_176),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_183),
.C(n_158),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_162),
.C(n_167),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_186),
.C(n_187),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_176),
.Y(n_187)
);

AO22x1_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_180),
.B1(n_22),
.B2(n_21),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_30),
.B(n_32),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_189),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_21),
.Y(n_194)
);


endmodule