module fake_aes_3652_n_472 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_472);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_472;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_73;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g69 ( .A(n_63), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_49), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_35), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_8), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_19), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_26), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_36), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_3), .Y(n_76) );
INVxp33_ASAP7_75t_SL g77 ( .A(n_16), .Y(n_77) );
BUFx2_ASAP7_75t_L g78 ( .A(n_31), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_62), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_37), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_14), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_13), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_22), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_38), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_65), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_15), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_47), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_57), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_30), .Y(n_89) );
CKINVDCx14_ASAP7_75t_R g90 ( .A(n_13), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_43), .Y(n_91) );
CKINVDCx14_ASAP7_75t_R g92 ( .A(n_41), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_50), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_25), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_42), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_1), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_51), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_46), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_64), .Y(n_99) );
INVxp33_ASAP7_75t_L g100 ( .A(n_21), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_78), .Y(n_101) );
INVx3_ASAP7_75t_L g102 ( .A(n_79), .Y(n_102) );
OA21x2_ASAP7_75t_L g103 ( .A1(n_69), .A2(n_0), .B(n_1), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_69), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_78), .B(n_0), .Y(n_105) );
OAI21x1_ASAP7_75t_L g106 ( .A1(n_79), .A2(n_32), .B(n_67), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_79), .Y(n_107) );
AND2x4_ASAP7_75t_L g108 ( .A(n_80), .B(n_2), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_70), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_80), .B(n_2), .Y(n_110) );
INVx3_ASAP7_75t_L g111 ( .A(n_87), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_87), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_87), .Y(n_113) );
OR2x2_ASAP7_75t_L g114 ( .A(n_100), .B(n_3), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_71), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_97), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_97), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_71), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_90), .B(n_4), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_90), .B(n_4), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_72), .B(n_5), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_97), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_108), .B(n_72), .Y(n_123) );
AND2x6_ASAP7_75t_L g124 ( .A(n_108), .B(n_74), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g125 ( .A(n_101), .B(n_91), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_107), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_107), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_102), .Y(n_128) );
INVx4_ASAP7_75t_SL g129 ( .A(n_108), .Y(n_129) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_108), .B(n_74), .Y(n_130) );
AND2x6_ASAP7_75t_L g131 ( .A(n_108), .B(n_75), .Y(n_131) );
INVx2_ASAP7_75t_SL g132 ( .A(n_108), .Y(n_132) );
AND2x6_ASAP7_75t_L g133 ( .A(n_119), .B(n_75), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_119), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_104), .B(n_92), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_104), .B(n_91), .Y(n_136) );
INVx4_ASAP7_75t_L g137 ( .A(n_103), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_116), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_116), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_104), .B(n_86), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_116), .Y(n_141) );
INVx4_ASAP7_75t_L g142 ( .A(n_103), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_107), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_107), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_126), .Y(n_145) );
OAI22xp5_ASAP7_75t_SL g146 ( .A1(n_130), .A2(n_77), .B1(n_82), .B2(n_114), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_128), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_130), .A2(n_120), .B1(n_119), .B2(n_103), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_134), .A2(n_110), .B(n_114), .C(n_105), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_126), .Y(n_150) );
INVx5_ASAP7_75t_L g151 ( .A(n_124), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_129), .B(n_120), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_127), .Y(n_153) );
AND3x2_ASAP7_75t_SL g154 ( .A(n_133), .B(n_122), .C(n_112), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_133), .A2(n_120), .B1(n_115), .B2(n_118), .Y(n_156) );
INVx1_ASAP7_75t_SL g157 ( .A(n_129), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_143), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_128), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_137), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_137), .Y(n_161) );
NAND2x1p5_ASAP7_75t_L g162 ( .A(n_123), .B(n_103), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_129), .B(n_114), .Y(n_163) );
BUFx12f_ASAP7_75t_L g164 ( .A(n_133), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_135), .B(n_110), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_133), .A2(n_103), .B1(n_109), .B2(n_118), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_124), .B(n_109), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_124), .B(n_115), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_143), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_124), .B(n_115), .Y(n_171) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_151), .B(n_128), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_164), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_164), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_149), .A2(n_125), .B(n_132), .C(n_121), .Y(n_176) );
NAND3xp33_ASAP7_75t_L g177 ( .A(n_167), .B(n_137), .C(n_142), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_145), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_164), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
AOI22xp33_ASAP7_75t_SL g181 ( .A1(n_146), .A2(n_133), .B1(n_124), .B2(n_131), .Y(n_181) );
OR2x6_ASAP7_75t_L g182 ( .A(n_163), .B(n_123), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_160), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_160), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_160), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_151), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_146), .A2(n_133), .B1(n_131), .B2(n_124), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_151), .B(n_129), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_151), .B(n_129), .Y(n_191) );
INVx2_ASAP7_75t_SL g192 ( .A(n_151), .Y(n_192) );
BUFx2_ASAP7_75t_L g193 ( .A(n_163), .Y(n_193) );
CKINVDCx6p67_ASAP7_75t_R g194 ( .A(n_151), .Y(n_194) );
CKINVDCx6p67_ASAP7_75t_R g195 ( .A(n_163), .Y(n_195) );
INVx5_ASAP7_75t_L g196 ( .A(n_152), .Y(n_196) );
INVx1_ASAP7_75t_SL g197 ( .A(n_153), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_156), .A2(n_131), .B1(n_124), .B2(n_123), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_156), .B(n_123), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_199), .B(n_166), .Y(n_200) );
INVx3_ASAP7_75t_SL g201 ( .A(n_195), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_173), .Y(n_202) );
OAI21x1_ASAP7_75t_L g203 ( .A1(n_177), .A2(n_106), .B(n_165), .Y(n_203) );
OAI221xp5_ASAP7_75t_L g204 ( .A1(n_181), .A2(n_148), .B1(n_136), .B2(n_169), .C(n_168), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_173), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_178), .Y(n_206) );
NAND2x1_ASAP7_75t_L g207 ( .A(n_186), .B(n_153), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_176), .A2(n_132), .B(n_171), .C(n_169), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_178), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_199), .B(n_140), .Y(n_210) );
AO31x2_ASAP7_75t_L g211 ( .A1(n_180), .A2(n_142), .A3(n_113), .B(n_117), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_195), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_183), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_197), .B(n_140), .Y(n_214) );
INVx6_ASAP7_75t_L g215 ( .A(n_196), .Y(n_215) );
INVx6_ASAP7_75t_L g216 ( .A(n_196), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_187), .A2(n_131), .B1(n_171), .B2(n_140), .Y(n_217) );
CKINVDCx8_ASAP7_75t_R g218 ( .A(n_174), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_183), .Y(n_219) );
AOI221xp5_ASAP7_75t_L g220 ( .A1(n_180), .A2(n_140), .B1(n_81), .B2(n_155), .C(n_170), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_213), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_200), .A2(n_198), .B1(n_190), .B2(n_182), .Y(n_222) );
OR2x2_ASAP7_75t_L g223 ( .A(n_205), .B(n_190), .Y(n_223) );
AO31x2_ASAP7_75t_L g224 ( .A1(n_208), .A2(n_117), .A3(n_122), .B(n_113), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_213), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_214), .A2(n_198), .B1(n_210), .B2(n_209), .Y(n_226) );
NAND3xp33_ASAP7_75t_L g227 ( .A(n_204), .B(n_177), .C(n_220), .Y(n_227) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_203), .A2(n_106), .B(n_117), .Y(n_228) );
OAI211xp5_ASAP7_75t_L g229 ( .A1(n_218), .A2(n_73), .B(n_96), .C(n_76), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_205), .B(n_155), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_209), .Y(n_231) );
AOI22xp33_ASAP7_75t_SL g232 ( .A1(n_212), .A2(n_174), .B1(n_175), .B2(n_196), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_202), .A2(n_196), .B1(n_193), .B2(n_182), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_206), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_219), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_203), .A2(n_185), .B(n_184), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_215), .A2(n_196), .B1(n_182), .B2(n_131), .Y(n_237) );
OAI22xp5_ASAP7_75t_SL g238 ( .A1(n_218), .A2(n_182), .B1(n_84), .B2(n_154), .Y(n_238) );
OAI211xp5_ASAP7_75t_L g239 ( .A1(n_217), .A2(n_76), .B(n_84), .C(n_102), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_231), .Y(n_240) );
NAND3xp33_ASAP7_75t_L g241 ( .A(n_227), .B(n_116), .C(n_207), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_221), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_221), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_222), .A2(n_216), .B1(n_215), .B2(n_201), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_231), .Y(n_245) );
AOI221xp5_ASAP7_75t_L g246 ( .A1(n_229), .A2(n_102), .B1(n_111), .B2(n_117), .C(n_112), .Y(n_246) );
OAI22xp33_ASAP7_75t_L g247 ( .A1(n_222), .A2(n_201), .B1(n_212), .B2(n_215), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_221), .Y(n_248) );
INVx1_ASAP7_75t_SL g249 ( .A(n_235), .Y(n_249) );
OR2x2_ASAP7_75t_L g250 ( .A(n_223), .B(n_211), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_225), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_234), .Y(n_252) );
AOI21x1_ASAP7_75t_L g253 ( .A1(n_236), .A2(n_207), .B(n_106), .Y(n_253) );
NOR2x1_ASAP7_75t_R g254 ( .A(n_235), .B(n_175), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_234), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_225), .Y(n_256) );
OAI22xp33_ASAP7_75t_L g257 ( .A1(n_226), .A2(n_216), .B1(n_215), .B2(n_175), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_238), .A2(n_216), .B1(n_131), .B2(n_179), .Y(n_258) );
OAI33xp33_ASAP7_75t_L g259 ( .A1(n_226), .A2(n_99), .A3(n_85), .B1(n_88), .B2(n_93), .B3(n_95), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_240), .B(n_225), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_250), .B(n_230), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_240), .B(n_224), .Y(n_262) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_259), .A2(n_239), .B1(n_227), .B2(n_83), .C(n_85), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_245), .Y(n_264) );
AND2x2_ASAP7_75t_SL g265 ( .A(n_254), .B(n_223), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_245), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_252), .B(n_230), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_242), .Y(n_268) );
O2A1O1Ixp5_ASAP7_75t_L g269 ( .A1(n_247), .A2(n_219), .B(n_122), .C(n_112), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_252), .B(n_224), .Y(n_270) );
OR2x2_ASAP7_75t_L g271 ( .A(n_249), .B(n_211), .Y(n_271) );
AOI33xp33_ASAP7_75t_L g272 ( .A1(n_255), .A2(n_93), .A3(n_95), .B1(n_98), .B2(n_99), .B3(n_122), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_242), .Y(n_273) );
INVx5_ASAP7_75t_L g274 ( .A(n_243), .Y(n_274) );
AND2x4_ASAP7_75t_SL g275 ( .A(n_244), .B(n_233), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_257), .A2(n_238), .B1(n_216), .B2(n_232), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_255), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_243), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_248), .B(n_224), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_248), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_258), .A2(n_111), .B1(n_237), .B2(n_103), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_249), .A2(n_228), .B1(n_154), .B2(n_170), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_246), .A2(n_111), .B1(n_98), .B2(n_112), .C(n_113), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_241), .A2(n_228), .B(n_157), .Y(n_284) );
NAND5xp2_ASAP7_75t_SL g285 ( .A(n_254), .B(n_89), .C(n_94), .D(n_7), .E(n_8), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_251), .B(n_211), .Y(n_286) );
OAI33xp33_ASAP7_75t_L g287 ( .A1(n_241), .A2(n_113), .A3(n_144), .B1(n_7), .B2(n_9), .B3(n_10), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_251), .B(n_224), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_256), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_270), .B(n_262), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_261), .B(n_256), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_270), .B(n_224), .Y(n_292) );
AND2x2_ASAP7_75t_SL g293 ( .A(n_265), .B(n_228), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_264), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_262), .B(n_211), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_264), .Y(n_296) );
AND3x1_ASAP7_75t_L g297 ( .A(n_276), .B(n_111), .C(n_6), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_266), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_266), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_277), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_265), .B(n_5), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_260), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_279), .B(n_211), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_260), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_267), .B(n_6), .Y(n_306) );
NOR4xp25_ASAP7_75t_L g307 ( .A(n_272), .B(n_9), .C(n_10), .D(n_11), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_267), .B(n_11), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_268), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_268), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_268), .Y(n_311) );
NAND3xp33_ASAP7_75t_L g312 ( .A(n_263), .B(n_116), .C(n_144), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_279), .B(n_116), .Y(n_313) );
NAND3xp33_ASAP7_75t_L g314 ( .A(n_274), .B(n_116), .C(n_139), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_288), .B(n_116), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_289), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_274), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_274), .Y(n_318) );
BUFx2_ASAP7_75t_SL g319 ( .A(n_274), .Y(n_319) );
OAI221xp5_ASAP7_75t_L g320 ( .A1(n_281), .A2(n_162), .B1(n_142), .B2(n_158), .C(n_147), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_271), .B(n_12), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_274), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_273), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_289), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_288), .B(n_253), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_273), .B(n_253), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_273), .B(n_12), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_265), .B(n_14), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_278), .B(n_15), .Y(n_329) );
NOR2x1p5_ASAP7_75t_L g330 ( .A(n_286), .B(n_194), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_297), .A2(n_275), .B1(n_287), .B2(n_282), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_314), .A2(n_282), .B(n_269), .Y(n_332) );
NAND3xp33_ASAP7_75t_L g333 ( .A(n_302), .B(n_274), .C(n_286), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_303), .B(n_280), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_306), .B(n_275), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_294), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_297), .A2(n_275), .B1(n_278), .B2(n_280), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_290), .B(n_278), .Y(n_338) );
OAI21xp33_ASAP7_75t_L g339 ( .A1(n_328), .A2(n_280), .B(n_283), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_294), .Y(n_340) );
OR2x6_ASAP7_75t_L g341 ( .A(n_319), .B(n_284), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_290), .B(n_16), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_321), .B(n_17), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_303), .B(n_17), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_321), .B(n_18), .Y(n_345) );
OAI322xp33_ASAP7_75t_L g346 ( .A1(n_308), .A2(n_285), .A3(n_162), .B1(n_20), .B2(n_21), .C1(n_18), .C2(n_19), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_296), .Y(n_347) );
XNOR2xp5_ASAP7_75t_L g348 ( .A(n_330), .B(n_20), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_305), .B(n_283), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_305), .B(n_142), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_296), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_298), .B(n_141), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_298), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_291), .B(n_158), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_299), .B(n_141), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_316), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_315), .B(n_285), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_295), .B(n_23), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_299), .B(n_141), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_324), .Y(n_360) );
AOI31xp33_ASAP7_75t_L g361 ( .A1(n_317), .A2(n_162), .A3(n_154), .B(n_172), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_293), .B(n_186), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_295), .B(n_24), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_300), .B(n_139), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_300), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_304), .B(n_27), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_301), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_304), .B(n_28), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_307), .A2(n_184), .B(n_185), .Y(n_369) );
INVxp67_ASAP7_75t_L g370 ( .A(n_319), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_315), .B(n_29), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_317), .B(n_33), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_327), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_313), .B(n_138), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_301), .B(n_139), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_309), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_293), .A2(n_165), .B1(n_161), .B2(n_147), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_293), .B(n_186), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_313), .B(n_138), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_335), .A2(n_330), .B1(n_292), .B2(n_313), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_336), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_340), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_337), .A2(n_314), .B(n_318), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_338), .B(n_325), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_347), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_356), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_342), .B(n_318), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_360), .B(n_313), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_357), .Y(n_389) );
INVx1_ASAP7_75t_SL g390 ( .A(n_348), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_351), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_334), .B(n_311), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_370), .B(n_322), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_334), .B(n_326), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_353), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_341), .B(n_322), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_365), .B(n_326), .Y(n_397) );
AOI21xp33_ASAP7_75t_L g398 ( .A1(n_343), .A2(n_329), .B(n_327), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_367), .B(n_311), .Y(n_399) );
NAND2xp33_ASAP7_75t_SL g400 ( .A(n_345), .B(n_322), .Y(n_400) );
NAND4xp25_ASAP7_75t_L g401 ( .A(n_344), .B(n_312), .C(n_329), .D(n_322), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_346), .B(n_312), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_373), .B(n_323), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_350), .B(n_310), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_364), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_358), .A2(n_310), .B1(n_309), .B2(n_320), .Y(n_406) );
NOR2xp33_ASAP7_75t_SL g407 ( .A(n_366), .B(n_310), .Y(n_407) );
NAND2x1_ASAP7_75t_L g408 ( .A(n_341), .B(n_191), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_375), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_371), .Y(n_410) );
XNOR2xp5_ASAP7_75t_L g411 ( .A(n_368), .B(n_165), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_352), .Y(n_412) );
AOI322xp5_ASAP7_75t_L g413 ( .A1(n_339), .A2(n_349), .A3(n_363), .B1(n_372), .B2(n_362), .C1(n_378), .C2(n_377), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_349), .A2(n_139), .B1(n_161), .B2(n_159), .Y(n_414) );
NOR3xp33_ASAP7_75t_L g415 ( .A(n_369), .B(n_161), .C(n_147), .Y(n_415) );
XNOR2x1_ASAP7_75t_L g416 ( .A(n_354), .B(n_34), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_341), .A2(n_147), .B1(n_159), .B2(n_192), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_355), .Y(n_418) );
NAND2xp33_ASAP7_75t_SL g419 ( .A(n_374), .B(n_191), .Y(n_419) );
XNOR2x1_ASAP7_75t_L g420 ( .A(n_379), .B(n_39), .Y(n_420) );
AOI211xp5_ASAP7_75t_L g421 ( .A1(n_332), .A2(n_188), .B(n_157), .C(n_186), .Y(n_421) );
OAI21xp33_ASAP7_75t_L g422 ( .A1(n_361), .A2(n_172), .B(n_189), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_355), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_359), .B(n_40), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_369), .A2(n_172), .B1(n_159), .B2(n_192), .C(n_189), .Y(n_425) );
OAI32xp33_ASAP7_75t_SL g426 ( .A1(n_333), .A2(n_44), .A3(n_45), .B1(n_48), .B2(n_52), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_338), .B(n_53), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_376), .Y(n_428) );
XNOR2x1_ASAP7_75t_L g429 ( .A(n_348), .B(n_54), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g430 ( .A1(n_337), .A2(n_188), .B1(n_186), .B2(n_159), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_336), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_356), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_334), .B(n_55), .Y(n_433) );
OAI21xp33_ASAP7_75t_L g434 ( .A1(n_331), .A2(n_188), .B(n_58), .Y(n_434) );
OAI211xp5_ASAP7_75t_L g435 ( .A1(n_331), .A2(n_68), .B(n_59), .C(n_60), .Y(n_435) );
AO22x2_ASAP7_75t_L g436 ( .A1(n_356), .A2(n_56), .B1(n_61), .B2(n_66), .Y(n_436) );
INVxp67_ASAP7_75t_L g437 ( .A(n_356), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_403), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_397), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_389), .A2(n_387), .B1(n_402), .B2(n_390), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_432), .B(n_396), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_434), .A2(n_410), .B1(n_380), .B2(n_401), .Y(n_443) );
AOI221xp5_ASAP7_75t_SL g444 ( .A1(n_437), .A2(n_386), .B1(n_383), .B2(n_432), .C(n_394), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_426), .A2(n_398), .B1(n_394), .B2(n_381), .C(n_382), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_411), .Y(n_446) );
AOI211xp5_ASAP7_75t_SL g447 ( .A1(n_435), .A2(n_398), .B(n_421), .C(n_425), .Y(n_447) );
NAND2xp33_ASAP7_75t_L g448 ( .A(n_419), .B(n_415), .Y(n_448) );
OAI211xp5_ASAP7_75t_SL g449 ( .A1(n_413), .A2(n_406), .B(n_417), .C(n_430), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_425), .A2(n_408), .B(n_433), .C(n_393), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_433), .B(n_429), .C(n_409), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_396), .A2(n_407), .B1(n_416), .B2(n_397), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_440), .Y(n_453) );
AOI322xp5_ASAP7_75t_L g454 ( .A1(n_444), .A2(n_384), .A3(n_431), .B1(n_395), .B2(n_385), .C1(n_391), .C2(n_423), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_448), .A2(n_420), .B(n_436), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_445), .A2(n_418), .B1(n_412), .B2(n_399), .C(n_404), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_449), .A2(n_427), .B(n_424), .C(n_422), .Y(n_457) );
AO22x2_ASAP7_75t_L g458 ( .A1(n_451), .A2(n_388), .B1(n_392), .B2(n_428), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_446), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_439), .B(n_405), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_453), .Y(n_461) );
NAND3xp33_ASAP7_75t_SL g462 ( .A(n_456), .B(n_452), .C(n_447), .Y(n_462) );
NOR4xp25_ASAP7_75t_L g463 ( .A(n_457), .B(n_450), .C(n_438), .D(n_442), .Y(n_463) );
NAND5xp2_ASAP7_75t_L g464 ( .A(n_455), .B(n_443), .C(n_441), .D(n_414), .E(n_424), .Y(n_464) );
OAI221xp5_ASAP7_75t_SL g465 ( .A1(n_463), .A2(n_454), .B1(n_458), .B2(n_459), .C(n_460), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_461), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_466), .Y(n_467) );
XNOR2x1_ASAP7_75t_L g468 ( .A(n_465), .B(n_464), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_467), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_469), .Y(n_470) );
INVxp67_ASAP7_75t_L g471 ( .A(n_470), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_471), .A2(n_468), .B(n_462), .Y(n_472) );
endmodule