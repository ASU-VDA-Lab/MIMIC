module fake_jpeg_22709_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_44),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_25),
.B1(n_27),
.B2(n_18),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_48),
.B1(n_53),
.B2(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_27),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_18),
.B1(n_25),
.B2(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_30),
.B1(n_25),
.B2(n_18),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_56),
.B(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_24),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_28),
.B1(n_20),
.B2(n_15),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_60),
.B1(n_59),
.B2(n_58),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_30),
.B1(n_20),
.B2(n_19),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_0),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_31),
.A2(n_30),
.B1(n_21),
.B2(n_15),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_32),
.A2(n_30),
.B1(n_26),
.B2(n_17),
.Y(n_57)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_68),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_34),
.C(n_32),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_52),
.C(n_50),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_69),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_51),
.B(n_53),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_77),
.B(n_3),
.Y(n_100)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_24),
.B1(n_34),
.B2(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_75),
.Y(n_81)
);

BUFx2_ASAP7_75t_SL g71 ( 
.A(n_45),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_74),
.Y(n_91)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_43),
.A2(n_60),
.B1(n_59),
.B2(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_55),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_54),
.B(n_47),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_50),
.Y(n_87)
);

BUFx4f_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_92),
.A2(n_99),
.B1(n_72),
.B2(n_73),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_100),
.Y(n_110)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_58),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_55),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_48),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_82),
.B(n_100),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_104),
.B(n_105),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_79),
.B(n_65),
.C(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_80),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_90),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_122),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_129),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_84),
.B1(n_89),
.B2(n_98),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_137),
.B1(n_92),
.B2(n_4),
.Y(n_152)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_89),
.C(n_82),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_136),
.C(n_108),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_112),
.B(n_106),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_84),
.B1(n_114),
.B2(n_116),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_107),
.C(n_111),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_R g139 ( 
.A1(n_120),
.A2(n_110),
.B(n_105),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_140),
.B1(n_150),
.B2(n_152),
.Y(n_159)
);

OAI22x1_ASAP7_75t_SL g140 ( 
.A1(n_133),
.A2(n_132),
.B1(n_122),
.B2(n_135),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_146),
.C(n_130),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_149),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_110),
.C(n_102),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_124),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_104),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_76),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_148),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_135),
.A2(n_113),
.B1(n_92),
.B2(n_55),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_153),
.Y(n_167)
);

XOR2x2_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_128),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_151),
.B(n_144),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_136),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_146),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_165),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_160),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_127),
.B1(n_134),
.B2(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_164),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_161),
.C(n_153),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_168),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_150),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_172),
.C(n_175),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_11),
.C(n_12),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_175),
.C(n_170),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_181),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_171),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_159),
.C(n_155),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_156),
.C(n_12),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_183),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_176),
.B(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_187),
.Y(n_195)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_166),
.Y(n_190)
);

XNOR2x1_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_9),
.Y(n_193)
);

OAI221xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_191),
.A2(n_193),
.B(n_194),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_8),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_192),
.B(n_9),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_184),
.A2(n_189),
.B(n_188),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_196),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_195),
.B(n_190),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_198),
.C(n_9),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_199),
.Y(n_203)
);


endmodule