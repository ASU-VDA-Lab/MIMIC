module fake_jpeg_26619_n_219 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_219);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx2_ASAP7_75t_SL g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_25),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_29),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_11),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_17),
.B1(n_10),
.B2(n_12),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_39),
.B1(n_13),
.B2(n_21),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_10),
.B1(n_17),
.B2(n_16),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_20),
.B1(n_14),
.B2(n_13),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_28),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_10),
.B1(n_12),
.B2(n_11),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_12),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_44),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_29),
.B(n_22),
.C(n_23),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_53),
.B1(n_36),
.B2(n_14),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_16),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_23),
.B1(n_25),
.B2(n_10),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_46),
.B1(n_39),
.B2(n_38),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_33),
.B1(n_36),
.B2(n_31),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_33),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_69),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_31),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_21),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_32),
.C(n_27),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_73),
.C(n_55),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_66),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_4),
.B(n_9),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_46),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_45),
.B1(n_43),
.B2(n_51),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_24),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_70),
.B(n_67),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_85),
.B1(n_70),
.B2(n_71),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

MAJx2_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_55),
.C(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_87),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_47),
.B1(n_41),
.B2(n_42),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_88),
.B(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_60),
.B(n_41),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_38),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_95),
.Y(n_97)
);

OAI32xp33_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_13),
.A3(n_14),
.B1(n_20),
.B2(n_21),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_30),
.C(n_11),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_38),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

OA21x2_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_68),
.B(n_66),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_24),
.B1(n_30),
.B2(n_18),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_102),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_72),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_83),
.B1(n_96),
.B2(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_64),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_107),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_119),
.B(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_73),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_108),
.B(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_73),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_113),
.B(n_114),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_56),
.B1(n_49),
.B2(n_75),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_115),
.B1(n_15),
.B2(n_1),
.Y(n_139)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_75),
.B1(n_74),
.B2(n_38),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_38),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_24),
.C(n_18),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_20),
.B(n_15),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_119),
.B(n_101),
.Y(n_149)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_130),
.Y(n_154)
);

AOI22x1_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_77),
.B1(n_85),
.B2(n_79),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_127),
.B1(n_133),
.B2(n_138),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_98),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_132),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_94),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_28),
.C(n_27),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_135),
.C(n_144),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_11),
.C(n_18),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_139),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_4),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_142),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_4),
.Y(n_144)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_150),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_156),
.Y(n_170)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_126),
.A2(n_103),
.B1(n_117),
.B2(n_109),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_134),
.B1(n_114),
.B2(n_116),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_128),
.C(n_129),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_155),
.C(n_156),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_118),
.C(n_113),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_108),
.C(n_100),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_100),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_148),
.A2(n_132),
.B1(n_124),
.B2(n_139),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_164),
.A2(n_150),
.B1(n_146),
.B2(n_153),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_175),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_135),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_174),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_147),
.C(n_160),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_173),
.C(n_155),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_144),
.C(n_141),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_163),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_145),
.B1(n_134),
.B2(n_2),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_145),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_134),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_187),
.Y(n_195)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_167),
.B(n_161),
.CI(n_157),
.CON(n_181),
.SN(n_181)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_183),
.B1(n_5),
.B2(n_7),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_157),
.C(n_161),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_173),
.C(n_177),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_158),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_162),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_172),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_176),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_191),
.C(n_178),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_196),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_180),
.B(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_193),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_4),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_0),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_198),
.Y(n_205)
);

NOR2x1_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_203),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_188),
.C(n_184),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_2),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_186),
.B(n_184),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_189),
.C(n_183),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_206),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_5),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_200),
.A2(n_5),
.A3(n_7),
.B1(n_2),
.B2(n_3),
.C1(n_8),
.C2(n_6),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_8),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_3),
.C(n_6),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_213),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_3),
.C(n_8),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_208),
.C(n_1),
.Y(n_215)
);

OAI21x1_ASAP7_75t_SL g216 ( 
.A1(n_215),
.A2(n_211),
.B(n_8),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_214),
.B1(n_0),
.B2(n_1),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_0),
.C(n_1),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_0),
.Y(n_219)
);


endmodule