module fake_jpeg_12435_n_537 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_537);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_537;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_14),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_6),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_60),
.B(n_65),
.Y(n_141)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_61),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_30),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_62),
.B(n_68),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_64),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_67),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_9),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_72),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_73),
.Y(n_150)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_76),
.Y(n_172)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_77),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_33),
.B(n_16),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_80),
.B(n_85),
.Y(n_154)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_82),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_41),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_83),
.B(n_100),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_41),
.A2(n_9),
.B1(n_14),
.B2(n_3),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_84),
.A2(n_98),
.B1(n_114),
.B2(n_112),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_40),
.B(n_24),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_86),
.Y(n_129)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_40),
.B(n_7),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_88),
.B(n_109),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_90),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_93),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_95),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

CKINVDCx6p67_ASAP7_75t_R g193 ( 
.A(n_97),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_98),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_37),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_105),
.Y(n_182)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_24),
.B(n_6),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_18),
.Y(n_110)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_10),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_111),
.B(n_13),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_20),
.Y(n_113)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_20),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_122),
.Y(n_126)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_46),
.Y(n_118)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_29),
.Y(n_119)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_18),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_27),
.Y(n_140)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_34),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_45),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_137),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_140),
.B(n_155),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_39),
.B1(n_22),
.B2(n_21),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_142),
.A2(n_151),
.B1(n_157),
.B2(n_171),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_95),
.A2(n_39),
.B1(n_22),
.B2(n_21),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_143),
.A2(n_144),
.B(n_167),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_83),
.A2(n_48),
.B1(n_43),
.B2(n_54),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_48),
.B1(n_52),
.B2(n_54),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_62),
.B(n_53),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_153),
.B(n_163),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_68),
.B(n_53),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_47),
.B1(n_38),
.B2(n_32),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_88),
.B(n_47),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_170),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_160),
.B(n_2),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_38),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_79),
.A2(n_32),
.B1(n_27),
.B2(n_35),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_70),
.B(n_5),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_73),
.A2(n_11),
.B1(n_13),
.B2(n_3),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_74),
.B(n_4),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_194),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_82),
.A2(n_15),
.B1(n_4),
.B2(n_11),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_181),
.A2(n_183),
.B1(n_197),
.B2(n_199),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_59),
.A2(n_0),
.B1(n_2),
.B2(n_12),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_84),
.A2(n_12),
.B(n_13),
.C(n_15),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_191),
.A2(n_193),
.B(n_147),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_69),
.A2(n_0),
.B1(n_2),
.B2(n_15),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_198),
.A2(n_202),
.B1(n_126),
.B2(n_160),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_91),
.A2(n_96),
.B1(n_107),
.B2(n_99),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_117),
.A2(n_0),
.B1(n_2),
.B2(n_93),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_203),
.Y(n_275)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_183),
.A2(n_76),
.B1(n_0),
.B2(n_2),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_206),
.A2(n_224),
.B1(n_239),
.B2(n_251),
.Y(n_298)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_138),
.Y(n_208)
);

INVx3_ASAP7_75t_SL g272 ( 
.A(n_208),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_150),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_209),
.B(n_218),
.Y(n_312)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_210),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_137),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_211),
.B(n_225),
.Y(n_276)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_212),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_214),
.Y(n_293)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_215),
.Y(n_294)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_216),
.Y(n_310)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_217),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_135),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_220),
.Y(n_270)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_221),
.Y(n_278)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_146),
.Y(n_222)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_222),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_223),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_197),
.A2(n_141),
.B1(n_143),
.B2(n_154),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_130),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_150),
.A2(n_124),
.B1(n_128),
.B2(n_201),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_158),
.Y(n_227)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_227),
.Y(n_285)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_125),
.Y(n_228)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_228),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_231),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_127),
.B(n_155),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_232),
.B(n_233),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_168),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_145),
.Y(n_234)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_234),
.Y(n_288)
);

OA22x2_ASAP7_75t_L g235 ( 
.A1(n_157),
.A2(n_202),
.B1(n_191),
.B2(n_196),
.Y(n_235)
);

OA22x2_ASAP7_75t_L g320 ( 
.A1(n_235),
.A2(n_217),
.B1(n_262),
.B2(n_264),
.Y(n_320)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_145),
.Y(n_237)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_237),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_144),
.A2(n_167),
.B1(n_149),
.B2(n_178),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_175),
.A2(n_184),
.B1(n_129),
.B2(n_134),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_240),
.A2(n_257),
.B1(n_262),
.B2(n_264),
.Y(n_289)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_138),
.Y(n_241)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_241),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_165),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_242),
.B(n_248),
.Y(n_302)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_129),
.Y(n_243)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_243),
.Y(n_314)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_244),
.Y(n_319)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_245),
.B(n_247),
.Y(n_296)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_133),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_136),
.B(n_161),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_134),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_249),
.Y(n_280)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_139),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_250),
.B(n_252),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_171),
.A2(n_192),
.B1(n_188),
.B2(n_190),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_182),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_229),
.B1(n_238),
.B2(n_204),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_137),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_254),
.B(n_255),
.Y(n_308)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_148),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_165),
.B(n_166),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_256),
.B(n_258),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_134),
.A2(n_174),
.B1(n_131),
.B2(n_177),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_126),
.B(n_131),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_259),
.A2(n_249),
.B(n_219),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_148),
.A2(n_152),
.B1(n_186),
.B2(n_190),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_260),
.A2(n_206),
.B1(n_241),
.B2(n_208),
.Y(n_299)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_152),
.Y(n_261)
);

NAND2xp33_ASAP7_75t_R g290 ( 
.A(n_261),
.B(n_263),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_147),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_177),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_180),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_231),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_180),
.B(n_172),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_267),
.Y(n_273)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_172),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_268),
.Y(n_297)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_164),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_228),
.Y(n_304)
);

AOI32xp33_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_207),
.A3(n_213),
.B1(n_224),
.B2(n_265),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_274),
.B(n_277),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_253),
.A2(n_229),
.B1(n_246),
.B2(n_235),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_279),
.A2(n_321),
.B1(n_307),
.B2(n_277),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_282),
.B(n_318),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_L g353 ( 
.A1(n_299),
.A2(n_315),
.B1(n_275),
.B2(n_281),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_304),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_235),
.A2(n_260),
.B1(n_258),
.B2(n_218),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_305),
.A2(n_317),
.B1(n_298),
.B2(n_299),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_L g307 ( 
.A1(n_235),
.A2(n_225),
.B(n_219),
.C(n_209),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_SL g338 ( 
.A1(n_307),
.A2(n_320),
.B(n_290),
.C(n_321),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_247),
.B(n_252),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_286),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_222),
.A2(n_255),
.B1(n_269),
.B2(n_210),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_203),
.A2(n_205),
.B1(n_234),
.B2(n_237),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_268),
.A2(n_230),
.B1(n_244),
.B2(n_214),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_295),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_322),
.B(n_323),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_301),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_316),
.Y(n_324)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_324),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_303),
.B(n_223),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_325),
.B(n_331),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_326),
.A2(n_337),
.B1(n_347),
.B2(n_353),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_282),
.B(n_279),
.C(n_318),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_328),
.B(n_336),
.Y(n_369)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_329),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_330),
.A2(n_333),
.B1(n_334),
.B2(n_349),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_332),
.B(n_294),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_298),
.A2(n_320),
.B1(n_305),
.B2(n_274),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_320),
.A2(n_273),
.B1(n_302),
.B2(n_312),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_273),
.C(n_312),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_320),
.A2(n_302),
.B1(n_300),
.B2(n_289),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_338),
.A2(n_343),
.B(n_294),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_276),
.C(n_285),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_341),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_308),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_344),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_285),
.B(n_314),
.C(n_278),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_278),
.B(n_270),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_342),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_300),
.A2(n_297),
.B1(n_306),
.B2(n_288),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_296),
.B(n_314),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_317),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_352),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_297),
.A2(n_272),
.B1(n_288),
.B2(n_306),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_319),
.A2(n_272),
.B1(n_271),
.B2(n_291),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_348),
.A2(n_358),
.B1(n_359),
.B2(n_354),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_286),
.A2(n_271),
.B1(n_272),
.B2(n_319),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_283),
.Y(n_350)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_350),
.Y(n_373)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_283),
.Y(n_351)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_351),
.Y(n_375)
);

AND2x6_ASAP7_75t_L g352 ( 
.A(n_280),
.B(n_291),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_354),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_292),
.B(n_284),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_355),
.B(n_357),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_316),
.A2(n_292),
.B1(n_311),
.B2(n_281),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_356),
.A2(n_351),
.B1(n_349),
.B2(n_361),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_284),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_359),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_287),
.B(n_310),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_360),
.B(n_361),
.Y(n_388)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_341),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_363),
.B(n_389),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_346),
.A2(n_293),
.B(n_287),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_364),
.A2(n_371),
.B(n_377),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_365),
.B(n_378),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_346),
.A2(n_328),
.B(n_332),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_374),
.A2(n_380),
.B(n_371),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_346),
.A2(n_330),
.B(n_335),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_337),
.A2(n_326),
.B1(n_336),
.B2(n_340),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_379),
.A2(n_374),
.B(n_380),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_334),
.B(n_333),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_382),
.A2(n_364),
.B(n_377),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_360),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_384),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_385),
.A2(n_362),
.B1(n_370),
.B2(n_390),
.Y(n_408)
);

MAJx2_ASAP7_75t_L g386 ( 
.A(n_339),
.B(n_327),
.C(n_329),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_393),
.C(n_338),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_344),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_327),
.A2(n_343),
.B1(n_338),
.B2(n_331),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_390),
.A2(n_338),
.B1(n_353),
.B2(n_352),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_357),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_395),
.A2(n_408),
.B1(n_368),
.B2(n_365),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_387),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_419),
.Y(n_426)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_375),
.Y(n_397)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_388),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_399),
.Y(n_436)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_375),
.Y(n_400)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_400),
.Y(n_430)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_388),
.Y(n_401)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_401),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_367),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_402),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_403),
.B(n_413),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_379),
.A2(n_338),
.B1(n_324),
.B2(n_356),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_404),
.A2(n_409),
.B1(n_412),
.B2(n_415),
.Y(n_424)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_373),
.Y(n_405)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_405),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_406),
.B(n_386),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_380),
.A2(n_394),
.B1(n_374),
.B2(n_370),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_373),
.Y(n_410)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_410),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_411),
.A2(n_414),
.B(n_393),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_394),
.A2(n_372),
.B1(n_362),
.B2(n_363),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_372),
.A2(n_384),
.B(n_376),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_389),
.A2(n_368),
.B1(n_376),
.B2(n_382),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_381),
.Y(n_417)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_381),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_392),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_387),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_369),
.B(n_365),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_378),
.C(n_386),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_367),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_421),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_402),
.B(n_383),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_423),
.B(n_442),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_425),
.A2(n_440),
.B(n_407),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_427),
.A2(n_403),
.B1(n_398),
.B2(n_401),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_404),
.A2(n_415),
.B1(n_409),
.B2(n_412),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_428),
.A2(n_408),
.B1(n_395),
.B2(n_416),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_369),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_434),
.C(n_444),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_439),
.B(n_420),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_SL g440 ( 
.A(n_403),
.B(n_391),
.C(n_392),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_422),
.Y(n_442)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_443),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_413),
.B(n_385),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_422),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_447),
.A2(n_421),
.B1(n_400),
.B2(n_397),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_449),
.A2(n_465),
.B1(n_466),
.B2(n_429),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_454),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_468),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_439),
.B(n_420),
.Y(n_454)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_455),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_435),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_457),
.Y(n_474)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_435),
.Y(n_457)
);

AOI21x1_ASAP7_75t_SL g458 ( 
.A1(n_425),
.A2(n_398),
.B(n_407),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_R g473 ( 
.A(n_458),
.B(n_467),
.C(n_443),
.Y(n_473)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_443),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_459),
.B(n_463),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_433),
.A2(n_406),
.B(n_411),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_428),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_461),
.A2(n_464),
.B1(n_431),
.B2(n_433),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_416),
.C(n_414),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_440),
.C(n_426),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_399),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_424),
.A2(n_395),
.B1(n_419),
.B2(n_396),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_427),
.A2(n_417),
.B1(n_418),
.B2(n_405),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_424),
.A2(n_410),
.B1(n_366),
.B2(n_391),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_437),
.B(n_366),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_444),
.B(n_434),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_437),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_441),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_475),
.Y(n_488)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_473),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_476),
.A2(n_483),
.B(n_467),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_468),
.B(n_446),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_481),
.C(n_454),
.Y(n_491)
);

FAx1_ASAP7_75t_SL g478 ( 
.A(n_462),
.B(n_446),
.CI(n_430),
.CON(n_478),
.SN(n_478)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_478),
.B(n_480),
.Y(n_498)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_479),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_451),
.B(n_429),
.C(n_430),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_445),
.C(n_438),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_469),
.A2(n_445),
.B(n_438),
.Y(n_483)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_484),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_461),
.A2(n_441),
.B1(n_464),
.B2(n_448),
.Y(n_486)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_486),
.Y(n_496)
);

OAI21xp33_ASAP7_75t_L g489 ( 
.A1(n_485),
.A2(n_463),
.B(n_458),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_489),
.Y(n_501)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_490),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_477),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_472),
.A2(n_452),
.B(n_465),
.Y(n_492)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_492),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_480),
.B(n_450),
.C(n_449),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_481),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_474),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_484),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_471),
.A2(n_467),
.B(n_453),
.Y(n_499)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_499),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_491),
.C(n_493),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_503),
.B(n_510),
.Y(n_511)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_489),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_504),
.B(n_505),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_494),
.A2(n_475),
.B1(n_473),
.B2(n_460),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_499),
.A2(n_486),
.B1(n_483),
.B2(n_478),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_509),
.Y(n_519)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_490),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_513),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_500),
.B(n_498),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_508),
.B(n_488),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_495),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_488),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_516),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_502),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_504),
.A2(n_487),
.B(n_492),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_518),
.A2(n_496),
.B(n_482),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_511),
.B(n_509),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_520),
.A2(n_523),
.B(n_526),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_517),
.A2(n_501),
.B(n_506),
.Y(n_523)
);

MAJx2_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_519),
.C(n_478),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_516),
.B(n_482),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_525),
.B(n_515),
.C(n_514),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_520),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_530),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_528),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_531),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_521),
.B(n_532),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_529),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_522),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_470),
.Y(n_537)
);


endmodule