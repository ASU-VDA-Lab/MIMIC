module fake_jpeg_10374_n_312 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_8),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_58),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_18),
.B1(n_22),
.B2(n_21),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_59),
.B1(n_61),
.B2(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_54),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_22),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_23),
.C(n_34),
.Y(n_88)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_21),
.B1(n_18),
.B2(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_25),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_21),
.B1(n_18),
.B2(n_35),
.Y(n_61)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_28),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_39),
.A2(n_34),
.B1(n_32),
.B2(n_25),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_70),
.B(n_71),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_72),
.B(n_73),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_15),
.B(n_16),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_81),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_79),
.A2(n_91),
.B1(n_101),
.B2(n_30),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_86),
.Y(n_110)
);

OR2x4_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_27),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_60),
.B(n_17),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_22),
.Y(n_86)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_25),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_11),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_45),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_26),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_98),
.C(n_31),
.Y(n_121)
);

BUFx4f_ASAP7_75t_SL g95 ( 
.A(n_65),
.Y(n_95)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

AOI32xp33_ASAP7_75t_L g98 ( 
.A1(n_47),
.A2(n_39),
.A3(n_40),
.B1(n_29),
.B2(n_33),
.Y(n_98)
);

CKINVDCx12_ASAP7_75t_R g99 ( 
.A(n_50),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_20),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_17),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_67),
.Y(n_103)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_12),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_109),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_74),
.A2(n_47),
.B1(n_62),
.B2(n_66),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_113),
.A2(n_120),
.B1(n_80),
.B2(n_102),
.Y(n_161)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_116),
.Y(n_138)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_58),
.B1(n_49),
.B2(n_67),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_119),
.B1(n_128),
.B2(n_80),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_48),
.B1(n_51),
.B2(n_32),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_130),
.Y(n_139)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_96),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_71),
.A2(n_29),
.B1(n_26),
.B2(n_33),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_132),
.B(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_135),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_88),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_123),
.C(n_112),
.Y(n_164)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_140),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_146),
.B1(n_147),
.B2(n_161),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_86),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_145),
.Y(n_171)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_107),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_97),
.B1(n_79),
.B2(n_77),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_90),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_151),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_69),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_94),
.B(n_75),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_159),
.B(n_28),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_154),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_90),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_156),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_69),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_157),
.A2(n_123),
.B(n_109),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_76),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_163),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_117),
.A2(n_87),
.B(n_103),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_112),
.B(n_40),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_150),
.B(n_140),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_70),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_186),
.C(n_189),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_192),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_178),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_24),
.B(n_106),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_174),
.A2(n_187),
.B1(n_142),
.B2(n_134),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_161),
.B1(n_148),
.B2(n_137),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_175),
.A2(n_93),
.B1(n_143),
.B2(n_114),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_133),
.A2(n_115),
.B(n_111),
.Y(n_178)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_106),
.A3(n_124),
.B1(n_95),
.B2(n_111),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_115),
.B(n_124),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_185),
.B1(n_193),
.B2(n_183),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_24),
.B(n_106),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_81),
.C(n_83),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_135),
.A2(n_93),
.B1(n_125),
.B2(n_92),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_191),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_95),
.C(n_116),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_193),
.B(n_158),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_116),
.C(n_114),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_147),
.C(n_138),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_11),
.B(n_16),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_7),
.C(n_14),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_197),
.B(n_201),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_159),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_210),
.C(n_215),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_170),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_202),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_R g203 ( 
.A(n_174),
.B(n_163),
.C(n_139),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_203),
.B(n_205),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_154),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_141),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_184),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_216),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_213),
.A2(n_218),
.B1(n_204),
.B2(n_183),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_SL g214 ( 
.A1(n_184),
.A2(n_163),
.B(n_153),
.C(n_162),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_185),
.B1(n_172),
.B2(n_182),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_139),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_139),
.C(n_138),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_186),
.C(n_181),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_220),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_141),
.Y(n_219)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_221),
.A2(n_179),
.B1(n_188),
.B2(n_167),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_222),
.B(n_210),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_189),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_233),
.C(n_200),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_226),
.A2(n_228),
.B1(n_232),
.B2(n_235),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_241),
.B1(n_242),
.B2(n_19),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_166),
.B1(n_169),
.B2(n_180),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_166),
.B1(n_191),
.B2(n_167),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_19),
.B(n_1),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_168),
.B1(n_182),
.B2(n_165),
.Y(n_235)
);

AOI322xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_176),
.A3(n_172),
.B1(n_171),
.B2(n_194),
.C1(n_165),
.C2(n_153),
.Y(n_238)
);

AOI21xp33_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_198),
.B(n_217),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_162),
.B1(n_122),
.B2(n_82),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_122),
.B1(n_82),
.B2(n_2),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_234),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_255),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_SL g247 ( 
.A(n_237),
.B(n_240),
.C(n_243),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_250),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_214),
.B(n_199),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_231),
.C(n_233),
.Y(n_264)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_214),
.B(n_200),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_251),
.B(n_254),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_259),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_229),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_253),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_235),
.A2(n_226),
.B(n_230),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_236),
.B(n_7),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_242),
.Y(n_275)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_260),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_223),
.B(n_6),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_227),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_239),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_273),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_260),
.B(n_224),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_275),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_231),
.C(n_225),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_250),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_282),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_256),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_283),
.C(n_284),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_263),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_278),
.B(n_266),
.Y(n_294)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_251),
.B(n_248),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_280),
.A2(n_259),
.B(n_279),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_253),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_270),
.A2(n_224),
.B1(n_257),
.B2(n_252),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_271),
.B1(n_268),
.B2(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_287),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_240),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_277),
.B(n_275),
.Y(n_288)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_295),
.B(n_0),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_264),
.C(n_6),
.Y(n_297)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_262),
.B(n_247),
.Y(n_292)
);

A2O1A1O1Ixp25_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_15),
.B(n_13),
.C(n_9),
.D(n_8),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_9),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_296),
.A2(n_293),
.B(n_291),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_298),
.C(n_302),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_301),
.A2(n_303),
.B(n_0),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_0),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_299),
.C(n_2),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_1),
.C(n_2),
.Y(n_309)
);

AOI321xp33_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_3),
.A3(n_4),
.B1(n_304),
.B2(n_247),
.C(n_271),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_310),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_308),
.Y(n_312)
);


endmodule