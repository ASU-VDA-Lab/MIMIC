module fake_jpeg_2106_n_396 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_27),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_53),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_54),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_59),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_84),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_61),
.Y(n_178)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_19),
.B(n_9),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_93),
.Y(n_122)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

CKINVDCx9p33_ASAP7_75t_R g75 ( 
.A(n_27),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g157 ( 
.A(n_75),
.Y(n_157)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_77),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_79),
.B(n_35),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_80),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_81),
.Y(n_173)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_17),
.B(n_9),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

BUFx2_ASAP7_75t_SL g166 ( 
.A(n_87),
.Y(n_166)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_33),
.B(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_99),
.Y(n_123)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_92),
.B(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_8),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_97),
.Y(n_180)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g99 ( 
.A(n_27),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_100),
.Y(n_164)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_104),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_105),
.Y(n_129)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_SL g170 ( 
.A(n_103),
.Y(n_170)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_107),
.Y(n_135)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_41),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_SL g112 ( 
.A1(n_109),
.A2(n_110),
.B(n_47),
.Y(n_112)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_112),
.B(n_130),
.C(n_104),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_38),
.B1(n_47),
.B2(n_46),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_113),
.A2(n_132),
.B1(n_69),
.B2(n_71),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_65),
.A2(n_41),
.B1(n_33),
.B2(n_35),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_127),
.A2(n_128),
.B1(n_143),
.B2(n_153),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_79),
.A2(n_98),
.B1(n_80),
.B2(n_81),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_28),
.B1(n_46),
.B2(n_45),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_55),
.A2(n_45),
.B1(n_38),
.B2(n_28),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_77),
.B(n_32),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_149),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_148),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_77),
.B(n_24),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_56),
.A2(n_51),
.B1(n_42),
.B2(n_26),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_62),
.B(n_24),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_162),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_106),
.B(n_37),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_156),
.B(n_108),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_54),
.A2(n_37),
.B1(n_32),
.B2(n_29),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_159),
.A2(n_161),
.B1(n_167),
.B2(n_171),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_78),
.A2(n_29),
.B1(n_42),
.B2(n_31),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_89),
.B(n_51),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_58),
.A2(n_31),
.B1(n_26),
.B2(n_3),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_110),
.B(n_10),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_175),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_54),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_66),
.B(n_7),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_174),
.B(n_137),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_101),
.B(n_11),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_86),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_176),
.A2(n_179),
.B1(n_181),
.B2(n_171),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_61),
.A2(n_1),
.B1(n_5),
.B2(n_12),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_57),
.A2(n_1),
.B1(n_5),
.B2(n_13),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_87),
.B(n_102),
.C(n_57),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_182),
.A2(n_184),
.B(n_185),
.C(n_230),
.Y(n_265)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_186),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_74),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_187),
.B(n_196),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_188),
.B(n_201),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_179),
.A2(n_90),
.B1(n_97),
.B2(n_100),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_189),
.A2(n_193),
.B1(n_230),
.B2(n_186),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g277 ( 
.A(n_190),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_191),
.B(n_194),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_L g193 ( 
.A1(n_114),
.A2(n_15),
.B1(n_127),
.B2(n_135),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_151),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_119),
.B(n_139),
.C(n_151),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_195),
.B(n_212),
.C(n_221),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_152),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_125),
.A2(n_166),
.B1(n_155),
.B2(n_164),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_199),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_123),
.B(n_115),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_203),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_126),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_204),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_205),
.B(n_206),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_131),
.B(n_153),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_207),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_129),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_208),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_111),
.B(n_118),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_209),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_117),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_210),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_146),
.B(n_141),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_213),
.B(n_218),
.Y(n_258)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_116),
.Y(n_214)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_167),
.A2(n_143),
.B1(n_159),
.B2(n_124),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_217),
.A2(n_238),
.B1(n_195),
.B2(n_210),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_113),
.B(n_121),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_133),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_219),
.A2(n_223),
.B1(n_225),
.B2(n_227),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_173),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_220),
.B(n_221),
.Y(n_275)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_145),
.A2(n_180),
.B1(n_163),
.B2(n_120),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_222),
.A2(n_229),
.B1(n_231),
.B2(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_160),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_224),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_133),
.A2(n_138),
.B1(n_160),
.B2(n_116),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_117),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_226),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_140),
.B(n_134),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_140),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_232),
.B1(n_234),
.B2(n_236),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_172),
.A2(n_181),
.B1(n_170),
.B2(n_136),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_134),
.A2(n_136),
.B1(n_178),
.B2(n_170),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_178),
.A2(n_75),
.B1(n_65),
.B2(n_53),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_177),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_233),
.A2(n_237),
.B(n_239),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_151),
.A2(n_75),
.B1(n_65),
.B2(n_99),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_141),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_123),
.B(n_115),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_161),
.A2(n_60),
.B1(n_75),
.B2(n_128),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_151),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_141),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_243),
.A2(n_260),
.B1(n_268),
.B2(n_278),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_192),
.A2(n_217),
.B1(n_189),
.B2(n_204),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_246),
.A2(n_273),
.B1(n_280),
.B2(n_282),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_194),
.A2(n_239),
.B(n_216),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_254),
.A2(n_256),
.B(n_281),
.Y(n_288)
);

OAI32xp33_ASAP7_75t_L g257 ( 
.A1(n_187),
.A2(n_206),
.A3(n_216),
.B1(n_202),
.B2(n_205),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_261),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_193),
.A2(n_215),
.B1(n_196),
.B2(n_220),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_265),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_266),
.A2(n_280),
.B1(n_245),
.B2(n_244),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_200),
.A2(n_183),
.B1(n_198),
.B2(n_226),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_272),
.B(n_276),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_228),
.A2(n_224),
.B1(n_197),
.B2(n_211),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_190),
.C(n_232),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_236),
.A2(n_214),
.B1(n_182),
.B2(n_234),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_207),
.A2(n_204),
.B1(n_192),
.B2(n_223),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_207),
.A2(n_204),
.B1(n_192),
.B2(n_223),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_246),
.A2(n_207),
.B1(n_244),
.B2(n_282),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_283),
.A2(n_286),
.B1(n_302),
.B2(n_299),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_281),
.B(n_248),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_284),
.B(n_289),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_268),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_290),
.Y(n_314)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_252),
.Y(n_287)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_288),
.A2(n_310),
.B(n_250),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_263),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_262),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_292),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

XOR2x1_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_260),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_308),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_256),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_297),
.B(n_298),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_272),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_253),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_300),
.B(n_305),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_241),
.B(n_242),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_266),
.A2(n_243),
.B1(n_269),
.B2(n_247),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_258),
.A2(n_274),
.B(n_269),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_304),
.A2(n_306),
.B(n_277),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_253),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_278),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_271),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_307),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_271),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_247),
.A2(n_265),
.B1(n_273),
.B2(n_251),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_309),
.A2(n_302),
.B1(n_295),
.B2(n_306),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_255),
.B(n_276),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_L g311 ( 
.A1(n_296),
.A2(n_264),
.B1(n_249),
.B2(n_255),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_311),
.A2(n_313),
.B1(n_309),
.B2(n_283),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_270),
.C(n_264),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_293),
.C(n_310),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_307),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_319),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_308),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_299),
.A2(n_249),
.B1(n_270),
.B2(n_277),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_320),
.A2(n_328),
.B1(n_283),
.B2(n_306),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_301),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_303),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_286),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_327),
.B(n_330),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_304),
.A2(n_295),
.B(n_289),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_304),
.A2(n_288),
.B(n_297),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_312),
.Y(n_331)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_331),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_339),
.C(n_341),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_334),
.A2(n_296),
.B1(n_328),
.B2(n_319),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_326),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_343),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_313),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_294),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_329),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_294),
.C(n_285),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_284),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_340),
.B(n_342),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_305),
.C(n_300),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_321),
.B(n_290),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_291),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_347),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_346),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_298),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_335),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_350),
.A2(n_358),
.B1(n_334),
.B2(n_318),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_353),
.C(n_339),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_330),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_SL g365 ( 
.A(n_355),
.B(n_337),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_341),
.B(n_317),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_356),
.B(n_359),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_335),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_350),
.A2(n_332),
.B(n_325),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_361),
.A2(n_365),
.B(n_353),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_360),
.A2(n_332),
.B(n_327),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_362),
.A2(n_369),
.B(n_370),
.Y(n_373)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_357),
.Y(n_364)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_364),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_368),
.C(n_351),
.Y(n_372)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_357),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_367),
.B(n_323),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_338),
.C(n_343),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_360),
.A2(n_346),
.B(n_315),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_370),
.A2(n_364),
.B1(n_363),
.B2(n_361),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_371),
.A2(n_378),
.B1(n_329),
.B2(n_355),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_377),
.Y(n_383)
);

XNOR2x1_ASAP7_75t_SL g379 ( 
.A(n_374),
.B(n_366),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_376),
.Y(n_380)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_368),
.Y(n_377)
);

A2O1A1Ixp33_ASAP7_75t_L g378 ( 
.A1(n_362),
.A2(n_345),
.B(n_354),
.C(n_322),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_382),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_381),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_352),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_373),
.A2(n_348),
.B1(n_336),
.B2(n_349),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_384),
.B(n_380),
.Y(n_387)
);

A2O1A1Ixp33_ASAP7_75t_L g390 ( 
.A1(n_387),
.A2(n_388),
.B(n_378),
.C(n_371),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_383),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_385),
.B(n_372),
.C(n_379),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_391),
.Y(n_393)
);

OAI21xp33_ASAP7_75t_L g392 ( 
.A1(n_390),
.A2(n_386),
.B(n_375),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_386),
.B(n_382),
.C(n_381),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_392),
.B(n_375),
.C(n_374),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_393),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_377),
.Y(n_396)
);


endmodule