module fake_jpeg_1767_n_192 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_192);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_29),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_61),
.Y(n_84)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_54),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_48),
.Y(n_88)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_69),
.B(n_51),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_66),
.C(n_54),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_90),
.B(n_62),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_64),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_51),
.B1(n_59),
.B2(n_53),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_98),
.B1(n_82),
.B2(n_77),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_73),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_77),
.B1(n_59),
.B2(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_50),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_101),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_55),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_55),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_114),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_96),
.B1(n_102),
.B2(n_85),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_46),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_46),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_25),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_22),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_120),
.B(n_122),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_63),
.C(n_49),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_53),
.B1(n_56),
.B2(n_94),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_124),
.B1(n_107),
.B2(n_40),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_127),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_82),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_49),
.B1(n_46),
.B2(n_73),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_73),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_133),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_49),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_137),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_120),
.C(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_140),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

AO22x1_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_56),
.B1(n_85),
.B2(n_63),
.Y(n_141)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_142),
.B(n_36),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_45),
.B(n_44),
.C(n_41),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_134),
.A2(n_38),
.B(n_37),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_146),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_0),
.B(n_2),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_152),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_2),
.B(n_3),
.Y(n_152)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_159),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_6),
.B(n_7),
.Y(n_160)
);

NOR5xp2_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_161),
.C(n_146),
.D(n_152),
.E(n_10),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_127),
.A2(n_32),
.B(n_21),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_136),
.A3(n_139),
.B1(n_142),
.B2(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_169),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_172),
.B1(n_147),
.B2(n_146),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_19),
.C(n_18),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_170),
.C(n_160),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_8),
.C(n_9),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_174),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_156),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_175),
.A2(n_177),
.B(n_163),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_156),
.C(n_148),
.Y(n_176)
);

OA21x2_ASAP7_75t_SL g182 ( 
.A1(n_176),
.A2(n_168),
.B(n_167),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_155),
.B1(n_154),
.B2(n_11),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_9),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_170),
.B(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_181),
.B(n_182),
.Y(n_184)
);

AOI211xp5_ASAP7_75t_SL g185 ( 
.A1(n_183),
.A2(n_173),
.B(n_179),
.C(n_174),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_180),
.C(n_11),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_186),
.A2(n_184),
.B1(n_12),
.B2(n_13),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_17),
.C(n_12),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_10),
.B(n_13),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_14),
.C(n_15),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_15),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_191),
.B(n_16),
.Y(n_192)
);


endmodule