module real_aes_8351_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g427 ( .A(n_0), .Y(n_427) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_1), .A2(n_132), .B(n_135), .C(n_215), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_2), .A2(n_161), .B(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g502 ( .A(n_3), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_4), .B(n_191), .Y(n_190) );
AOI21xp33_ASAP7_75t_L g485 ( .A1(n_5), .A2(n_161), .B(n_486), .Y(n_485) );
AND2x6_ASAP7_75t_L g132 ( .A(n_6), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g228 ( .A(n_7), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_8), .B(n_43), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_9), .A2(n_160), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_10), .B(n_144), .Y(n_217) );
INVx1_ASAP7_75t_L g490 ( .A(n_11), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_12), .B(n_185), .Y(n_525) );
OAI22xp5_ASAP7_75t_SL g444 ( .A1(n_13), .A2(n_445), .B1(n_446), .B2(n_452), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_13), .Y(n_452) );
INVx1_ASAP7_75t_L g124 ( .A(n_14), .Y(n_124) );
INVx1_ASAP7_75t_L g537 ( .A(n_15), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_16), .A2(n_80), .B1(n_450), .B2(n_451), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_16), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_17), .A2(n_169), .B(n_250), .C(n_252), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_18), .B(n_191), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_19), .B(n_468), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_20), .B(n_161), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_21), .B(n_175), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_22), .A2(n_185), .B(n_236), .C(n_238), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_23), .B(n_191), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_24), .B(n_144), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_25), .A2(n_171), .B(n_252), .C(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_26), .B(n_144), .Y(n_199) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_27), .Y(n_126) );
INVx1_ASAP7_75t_L g198 ( .A(n_28), .Y(n_198) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_29), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_30), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_31), .B(n_144), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_32), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g167 ( .A(n_33), .Y(n_167) );
INVx1_ASAP7_75t_L g480 ( .A(n_34), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_35), .A2(n_447), .B1(n_448), .B2(n_449), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_35), .Y(n_447) );
INVx2_ASAP7_75t_L g130 ( .A(n_36), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_37), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_38), .A2(n_185), .B(n_186), .C(n_188), .Y(n_184) );
INVxp67_ASAP7_75t_L g170 ( .A(n_39), .Y(n_170) );
CKINVDCx14_ASAP7_75t_R g183 ( .A(n_40), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_41), .A2(n_135), .B(n_197), .C(n_201), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_42), .A2(n_132), .B(n_135), .C(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g479 ( .A(n_44), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_45), .A2(n_146), .B(n_226), .C(n_227), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_46), .B(n_144), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_47), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_48), .Y(n_163) );
INVx1_ASAP7_75t_L g234 ( .A(n_49), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_50), .Y(n_481) );
AOI222xp33_ASAP7_75t_SL g442 ( .A1(n_51), .A2(n_443), .B1(n_444), .B2(n_453), .C1(n_740), .C2(n_743), .Y(n_442) );
OAI22xp5_ASAP7_75t_SL g415 ( .A1(n_52), .A2(n_61), .B1(n_416), .B2(n_417), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_52), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_53), .B(n_161), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_54), .A2(n_135), .B1(n_238), .B2(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_55), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_56), .Y(n_499) );
CKINVDCx14_ASAP7_75t_R g224 ( .A(n_57), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_58), .A2(n_188), .B(n_226), .C(n_489), .Y(n_488) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_59), .A2(n_104), .B1(n_432), .B2(n_441), .C1(n_745), .C2(n_750), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_59), .A2(n_106), .B1(n_107), .B2(n_420), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_59), .Y(n_420) );
INVx1_ASAP7_75t_L g487 ( .A(n_60), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_61), .Y(n_417) );
INVx1_ASAP7_75t_L g133 ( .A(n_62), .Y(n_133) );
INVx1_ASAP7_75t_L g123 ( .A(n_63), .Y(n_123) );
INVx1_ASAP7_75t_SL g187 ( .A(n_64), .Y(n_187) );
OAI22xp5_ASAP7_75t_SL g414 ( .A1(n_65), .A2(n_415), .B1(n_418), .B2(n_419), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_65), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_66), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_67), .B(n_191), .Y(n_240) );
INVx1_ASAP7_75t_L g139 ( .A(n_68), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_SL g467 ( .A1(n_69), .A2(n_188), .B(n_468), .C(n_469), .Y(n_467) );
INVxp67_ASAP7_75t_L g470 ( .A(n_70), .Y(n_470) );
INVx1_ASAP7_75t_L g440 ( .A(n_71), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_72), .A2(n_161), .B(n_223), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_73), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_74), .A2(n_161), .B(n_247), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_75), .Y(n_483) );
INVx1_ASAP7_75t_L g543 ( .A(n_76), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_77), .A2(n_160), .B(n_162), .Y(n_159) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_78), .Y(n_195) );
INVx1_ASAP7_75t_L g248 ( .A(n_79), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_80), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_81), .A2(n_132), .B(n_135), .C(n_545), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_82), .A2(n_161), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g251 ( .A(n_83), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_84), .B(n_168), .Y(n_514) );
INVx2_ASAP7_75t_L g121 ( .A(n_85), .Y(n_121) );
INVx1_ASAP7_75t_L g216 ( .A(n_86), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_87), .B(n_468), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_88), .A2(n_132), .B(n_135), .C(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g424 ( .A(n_89), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g454 ( .A(n_89), .B(n_426), .Y(n_454) );
INVx2_ASAP7_75t_L g739 ( .A(n_89), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g134 ( .A1(n_90), .A2(n_135), .B(n_138), .C(n_148), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_91), .B(n_153), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_92), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_93), .A2(n_132), .B(n_135), .C(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_94), .Y(n_529) );
INVx1_ASAP7_75t_L g466 ( .A(n_95), .Y(n_466) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_96), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_97), .B(n_168), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_98), .B(n_119), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_99), .B(n_119), .Y(n_538) );
INVx2_ASAP7_75t_L g237 ( .A(n_100), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_101), .B(n_440), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_102), .A2(n_161), .B(n_465), .Y(n_464) );
OAI21xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_421), .B(n_429), .Y(n_104) );
INVxp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
XOR2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_414), .Y(n_107) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_108), .A2(n_454), .B1(n_455), .B2(n_736), .Y(n_453) );
INVx2_ASAP7_75t_L g744 ( .A(n_108), .Y(n_744) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_348), .Y(n_108) );
NAND5xp2_ASAP7_75t_L g109 ( .A(n_110), .B(n_277), .C(n_307), .D(n_328), .E(n_334), .Y(n_109) );
AOI221xp5_ASAP7_75t_SL g110 ( .A1(n_111), .A2(n_207), .B1(n_241), .B2(n_243), .C(n_254), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_204), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_176), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_SL g328 ( .A1(n_115), .A2(n_192), .B(n_329), .C(n_332), .Y(n_328) );
AND2x2_ASAP7_75t_L g398 ( .A(n_115), .B(n_193), .Y(n_398) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_154), .Y(n_115) );
AND2x2_ASAP7_75t_L g256 ( .A(n_116), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g260 ( .A(n_116), .B(n_257), .Y(n_260) );
OR2x2_ASAP7_75t_L g286 ( .A(n_116), .B(n_193), .Y(n_286) );
AND2x2_ASAP7_75t_L g288 ( .A(n_116), .B(n_179), .Y(n_288) );
AND2x2_ASAP7_75t_L g306 ( .A(n_116), .B(n_178), .Y(n_306) );
INVx1_ASAP7_75t_L g339 ( .A(n_116), .Y(n_339) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g206 ( .A(n_117), .Y(n_206) );
AND2x2_ASAP7_75t_L g242 ( .A(n_117), .B(n_179), .Y(n_242) );
AND2x2_ASAP7_75t_L g395 ( .A(n_117), .B(n_193), .Y(n_395) );
AO21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_125), .B(n_150), .Y(n_117) );
INVx3_ASAP7_75t_L g191 ( .A(n_118), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_118), .B(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_118), .B(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_SL g516 ( .A(n_118), .B(n_517), .Y(n_516) );
INVx4_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_119), .Y(n_180) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_119), .A2(n_464), .B(n_471), .Y(n_463) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g157 ( .A(n_120), .Y(n_157) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_121), .B(n_122), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
OAI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B(n_134), .Y(n_125) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_127), .A2(n_153), .B(n_195), .C(n_196), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_127), .A2(n_213), .B(n_214), .Y(n_212) );
OAI22xp33_ASAP7_75t_L g476 ( .A1(n_127), .A2(n_149), .B1(n_477), .B2(n_481), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_127), .A2(n_499), .B(n_500), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_127), .A2(n_543), .B(n_544), .Y(n_542) );
NAND2x1p5_ASAP7_75t_L g127 ( .A(n_128), .B(n_132), .Y(n_127) );
AND2x4_ASAP7_75t_L g161 ( .A(n_128), .B(n_132), .Y(n_161) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
INVx1_ASAP7_75t_L g239 ( .A(n_130), .Y(n_239) );
INVx1_ASAP7_75t_L g137 ( .A(n_131), .Y(n_137) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_131), .Y(n_142) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
INVx3_ASAP7_75t_L g169 ( .A(n_131), .Y(n_169) );
INVx1_ASAP7_75t_L g468 ( .A(n_131), .Y(n_468) );
INVx4_ASAP7_75t_SL g149 ( .A(n_132), .Y(n_149) );
BUFx3_ASAP7_75t_L g201 ( .A(n_132), .Y(n_201) );
INVx5_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
AND2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx3_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_136), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_143), .C(n_145), .Y(n_138) );
O2A1O1Ixp5_ASAP7_75t_L g215 ( .A1(n_140), .A2(n_145), .B(n_216), .C(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OAI22xp5_ASAP7_75t_SL g478 ( .A1(n_141), .A2(n_142), .B1(n_479), .B2(n_480), .Y(n_478) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx4_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
INVx4_ASAP7_75t_L g185 ( .A(n_144), .Y(n_185) );
INVx2_ASAP7_75t_L g226 ( .A(n_144), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_145), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_145), .A2(n_546), .B(n_547), .Y(n_545) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g252 ( .A(n_147), .Y(n_252) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_SL g162 ( .A1(n_149), .A2(n_163), .B(n_164), .C(n_165), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_149), .A2(n_164), .B(n_183), .C(n_184), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_SL g223 ( .A1(n_149), .A2(n_164), .B(n_224), .C(n_225), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_SL g233 ( .A1(n_149), .A2(n_164), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_SL g247 ( .A1(n_149), .A2(n_164), .B(n_248), .C(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_149), .A2(n_164), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_149), .A2(n_164), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_149), .A2(n_164), .B(n_534), .C(n_535), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
INVx1_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_152), .A2(n_521), .B(n_528), .Y(n_520) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g211 ( .A(n_153), .Y(n_211) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_153), .A2(n_222), .B(n_229), .Y(n_221) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_153), .A2(n_532), .B(n_538), .Y(n_531) );
AND2x2_ASAP7_75t_L g276 ( .A(n_154), .B(n_177), .Y(n_276) );
OR2x2_ASAP7_75t_L g280 ( .A(n_154), .B(n_193), .Y(n_280) );
AND2x2_ASAP7_75t_L g305 ( .A(n_154), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g352 ( .A(n_154), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_154), .B(n_314), .Y(n_400) );
AO21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_158), .B(n_173), .Y(n_154) );
INVx1_ASAP7_75t_L g258 ( .A(n_155), .Y(n_258) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_155), .A2(n_542), .B(n_548), .Y(n_541) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_SL g510 ( .A1(n_156), .A2(n_511), .B(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_157), .A2(n_476), .B(n_482), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_157), .B(n_483), .Y(n_482) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_157), .A2(n_498), .B(n_505), .Y(n_497) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OA21x2_ASAP7_75t_L g257 ( .A1(n_159), .A2(n_174), .B(n_258), .Y(n_257) );
BUFx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_166), .B(n_172), .Y(n_165) );
OAI22xp33_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B1(n_170), .B2(n_171), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_168), .A2(n_198), .B(n_199), .C(n_200), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_168), .A2(n_502), .B(n_503), .C(n_504), .Y(n_501) );
INVx5_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_169), .B(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_169), .B(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_169), .B(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_171), .B(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_171), .B(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_171), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g200 ( .A(n_172), .Y(n_200) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OAI322xp33_ASAP7_75t_L g401 ( .A1(n_176), .A2(n_337), .A3(n_360), .B1(n_381), .B2(n_402), .C1(n_404), .C2(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_177), .B(n_257), .Y(n_404) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_192), .Y(n_177) );
AND2x2_ASAP7_75t_L g205 ( .A(n_178), .B(n_206), .Y(n_205) );
AND2x4_ASAP7_75t_L g273 ( .A(n_178), .B(n_193), .Y(n_273) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g314 ( .A(n_179), .B(n_193), .Y(n_314) );
AND2x2_ASAP7_75t_L g358 ( .A(n_179), .B(n_192), .Y(n_358) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_190), .Y(n_179) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_180), .A2(n_232), .B(n_240), .Y(n_231) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_180), .A2(n_246), .B(n_253), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_185), .B(n_187), .Y(n_186) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_189), .Y(n_526) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_191), .A2(n_485), .B(n_491), .Y(n_484) );
AND2x2_ASAP7_75t_L g241 ( .A(n_192), .B(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g259 ( .A(n_192), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_192), .B(n_288), .Y(n_412) );
INVx3_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g204 ( .A(n_193), .B(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_193), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g326 ( .A(n_193), .B(n_257), .Y(n_326) );
AND2x2_ASAP7_75t_L g353 ( .A(n_193), .B(n_288), .Y(n_353) );
OR2x2_ASAP7_75t_L g409 ( .A(n_193), .B(n_260), .Y(n_409) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_202), .Y(n_193) );
INVx1_ASAP7_75t_SL g295 ( .A(n_204), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_205), .B(n_326), .Y(n_327) );
AND2x2_ASAP7_75t_L g361 ( .A(n_205), .B(n_351), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_205), .B(n_284), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_205), .B(n_406), .Y(n_405) );
OAI31xp33_ASAP7_75t_L g379 ( .A1(n_207), .A2(n_241), .A3(n_380), .B(n_382), .Y(n_379) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_220), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_208), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g362 ( .A(n_208), .B(n_297), .Y(n_362) );
OR2x2_ASAP7_75t_L g369 ( .A(n_208), .B(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g381 ( .A(n_208), .B(n_270), .Y(n_381) );
CKINVDCx16_ASAP7_75t_R g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g315 ( .A(n_209), .B(n_316), .Y(n_315) );
BUFx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g243 ( .A(n_210), .B(n_244), .Y(n_243) );
INVx4_ASAP7_75t_L g264 ( .A(n_210), .Y(n_264) );
AND2x2_ASAP7_75t_L g301 ( .A(n_210), .B(n_245), .Y(n_301) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_218), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_211), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_211), .B(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_211), .B(n_420), .Y(n_548) );
AND2x2_ASAP7_75t_L g300 ( .A(n_220), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_SL g370 ( .A(n_220), .Y(n_370) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_230), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_221), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g270 ( .A(n_221), .B(n_231), .Y(n_270) );
INVx2_ASAP7_75t_L g290 ( .A(n_221), .Y(n_290) );
AND2x2_ASAP7_75t_L g304 ( .A(n_221), .B(n_231), .Y(n_304) );
AND2x2_ASAP7_75t_L g311 ( .A(n_221), .B(n_267), .Y(n_311) );
BUFx3_ASAP7_75t_L g321 ( .A(n_221), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_221), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g266 ( .A(n_230), .Y(n_266) );
AND2x2_ASAP7_75t_L g274 ( .A(n_230), .B(n_264), .Y(n_274) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g244 ( .A(n_231), .B(n_245), .Y(n_244) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_231), .Y(n_298) );
INVx2_ASAP7_75t_L g504 ( .A(n_238), .Y(n_504) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_SL g281 ( .A(n_242), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_242), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_242), .B(n_351), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_243), .B(n_321), .Y(n_374) );
INVx1_ASAP7_75t_SL g408 ( .A(n_243), .Y(n_408) );
INVx1_ASAP7_75t_SL g316 ( .A(n_244), .Y(n_316) );
INVx1_ASAP7_75t_SL g267 ( .A(n_245), .Y(n_267) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_245), .Y(n_278) );
OR2x2_ASAP7_75t_L g289 ( .A(n_245), .B(n_264), .Y(n_289) );
AND2x2_ASAP7_75t_L g303 ( .A(n_245), .B(n_264), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_245), .B(n_293), .Y(n_355) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_259), .B(n_261), .C(n_272), .Y(n_254) );
AOI31xp33_ASAP7_75t_L g371 ( .A1(n_255), .A2(n_372), .A3(n_373), .B(n_374), .Y(n_371) );
AND2x2_ASAP7_75t_L g344 ( .A(n_256), .B(n_273), .Y(n_344) );
BUFx3_ASAP7_75t_L g284 ( .A(n_257), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_257), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g320 ( .A(n_257), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_257), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g275 ( .A(n_260), .Y(n_275) );
OAI222xp33_ASAP7_75t_L g384 ( .A1(n_260), .A2(n_385), .B1(n_388), .B2(n_389), .C1(n_390), .C2(n_391), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_268), .Y(n_261) );
INVx1_ASAP7_75t_L g390 ( .A(n_262), .Y(n_390) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_264), .B(n_267), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_264), .B(n_290), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_264), .B(n_265), .Y(n_360) );
INVx1_ASAP7_75t_L g411 ( .A(n_264), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_265), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g413 ( .A(n_265), .Y(n_413) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g293 ( .A(n_266), .Y(n_293) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_267), .Y(n_336) );
AOI32xp33_ASAP7_75t_L g272 ( .A1(n_268), .A2(n_273), .A3(n_274), .B1(n_275), .B2(n_276), .Y(n_272) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_270), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g347 ( .A(n_270), .Y(n_347) );
OR2x2_ASAP7_75t_L g388 ( .A(n_270), .B(n_289), .Y(n_388) );
INVx1_ASAP7_75t_L g324 ( .A(n_271), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_273), .B(n_284), .Y(n_309) );
INVx3_ASAP7_75t_L g318 ( .A(n_273), .Y(n_318) );
AOI322xp5_ASAP7_75t_L g334 ( .A1(n_273), .A2(n_318), .A3(n_335), .B1(n_337), .B2(n_340), .C1(n_344), .C2(n_345), .Y(n_334) );
AND2x2_ASAP7_75t_L g310 ( .A(n_274), .B(n_311), .Y(n_310) );
INVxp67_ASAP7_75t_L g387 ( .A(n_274), .Y(n_387) );
A2O1A1O1Ixp25_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_279), .B(n_282), .C(n_290), .D(n_291), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_278), .B(n_321), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
OAI221xp5_ASAP7_75t_L g291 ( .A1(n_280), .A2(n_292), .B1(n_295), .B2(n_296), .C(n_299), .Y(n_291) );
INVx1_ASAP7_75t_SL g406 ( .A(n_280), .Y(n_406) );
AOI21xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_287), .B(n_289), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_284), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OAI221xp5_ASAP7_75t_SL g376 ( .A1(n_286), .A2(n_370), .B1(n_377), .B2(n_378), .C(n_379), .Y(n_376) );
OAI222xp33_ASAP7_75t_L g407 ( .A1(n_287), .A2(n_408), .B1(n_409), .B2(n_410), .C1(n_412), .C2(n_413), .Y(n_407) );
AND2x2_ASAP7_75t_L g365 ( .A(n_288), .B(n_351), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_288), .A2(n_303), .B(n_350), .Y(n_377) );
INVx1_ASAP7_75t_L g391 ( .A(n_288), .Y(n_391) );
INVx2_ASAP7_75t_SL g294 ( .A(n_289), .Y(n_294) );
AND2x2_ASAP7_75t_L g297 ( .A(n_290), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_SL g331 ( .A(n_293), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_293), .B(n_303), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_294), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_294), .B(n_304), .Y(n_333) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OAI21xp5_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_302), .B(n_305), .Y(n_299) );
INVx1_ASAP7_75t_SL g317 ( .A(n_301), .Y(n_317) );
AND2x2_ASAP7_75t_L g364 ( .A(n_301), .B(n_347), .Y(n_364) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x2_ASAP7_75t_L g403 ( .A(n_303), .B(n_321), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_304), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g389 ( .A(n_305), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_310), .B1(n_312), .B2(n_319), .C(n_322), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_315), .B1(n_317), .B2(n_318), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI22xp33_ASAP7_75t_L g322 ( .A1(n_316), .A2(n_323), .B1(n_325), .B2(n_327), .Y(n_322) );
OR2x2_ASAP7_75t_L g393 ( .A(n_317), .B(n_321), .Y(n_393) );
OR2x2_ASAP7_75t_L g396 ( .A(n_317), .B(n_331), .Y(n_396) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI221xp5_ASAP7_75t_L g392 ( .A1(n_338), .A2(n_393), .B1(n_394), .B2(n_396), .C(n_397), .Y(n_392) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND3xp33_ASAP7_75t_SL g348 ( .A(n_349), .B(n_363), .C(n_375), .Y(n_348) );
AOI222xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_354), .B1(n_356), .B2(n_359), .C1(n_361), .C2(n_362), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_351), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g373 ( .A(n_353), .Y(n_373) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_366), .B2(n_368), .C(n_371), .Y(n_363) );
INVx1_ASAP7_75t_L g378 ( .A(n_364), .Y(n_378) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI21xp33_ASAP7_75t_L g397 ( .A1(n_368), .A2(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NOR5xp2_ASAP7_75t_L g375 ( .A(n_376), .B(n_384), .C(n_392), .D(n_401), .E(n_407), .Y(n_375) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_415), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
BUFx2_ASAP7_75t_L g431 ( .A(n_424), .Y(n_431) );
INVx1_ASAP7_75t_SL g749 ( .A(n_424), .Y(n_749) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_425), .B(n_739), .Y(n_742) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g738 ( .A(n_426), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OA21x2_ASAP7_75t_L g751 ( .A1(n_431), .A2(n_437), .B(n_438), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_433), .Y(n_432) );
CKINVDCx6p67_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_438), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NOR2xp33_ASAP7_75t_SL g747 ( .A(n_437), .B(n_439), .Y(n_747) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_454), .A2(n_456), .B1(n_736), .B2(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_457), .B(n_673), .Y(n_456) );
NOR4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_603), .C(n_634), .D(n_653), .Y(n_457) );
NAND4xp25_ASAP7_75t_L g458 ( .A(n_459), .B(n_561), .C(n_576), .D(n_594), .Y(n_458) );
AOI222xp33_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_507), .B1(n_539), .B2(n_549), .C1(n_554), .C2(n_556), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_492), .Y(n_460) );
INVx1_ASAP7_75t_L g617 ( .A(n_461), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_472), .Y(n_461) );
AND2x2_ASAP7_75t_L g493 ( .A(n_462), .B(n_484), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_462), .B(n_496), .Y(n_646) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g553 ( .A(n_463), .B(n_474), .Y(n_553) );
AND2x2_ASAP7_75t_L g562 ( .A(n_463), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g588 ( .A(n_463), .Y(n_588) );
AND2x2_ASAP7_75t_L g609 ( .A(n_463), .B(n_474), .Y(n_609) );
BUFx2_ASAP7_75t_L g632 ( .A(n_463), .Y(n_632) );
AND2x2_ASAP7_75t_L g656 ( .A(n_463), .B(n_475), .Y(n_656) );
AND2x2_ASAP7_75t_L g720 ( .A(n_463), .B(n_484), .Y(n_720) );
AND2x2_ASAP7_75t_L g621 ( .A(n_472), .B(n_552), .Y(n_621) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_473), .B(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .Y(n_473) );
OR2x2_ASAP7_75t_L g581 ( .A(n_474), .B(n_497), .Y(n_581) );
AND2x2_ASAP7_75t_L g593 ( .A(n_474), .B(n_552), .Y(n_593) );
BUFx2_ASAP7_75t_L g725 ( .A(n_474), .Y(n_725) );
INVx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g495 ( .A(n_475), .B(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g575 ( .A(n_475), .B(n_497), .Y(n_575) );
AND2x2_ASAP7_75t_L g628 ( .A(n_475), .B(n_484), .Y(n_628) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_475), .Y(n_664) );
AND2x2_ASAP7_75t_L g551 ( .A(n_484), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_SL g563 ( .A(n_484), .Y(n_563) );
INVx2_ASAP7_75t_L g574 ( .A(n_484), .Y(n_574) );
BUFx2_ASAP7_75t_L g598 ( .A(n_484), .Y(n_598) );
AND2x2_ASAP7_75t_SL g655 ( .A(n_484), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
AOI332xp33_ASAP7_75t_L g576 ( .A1(n_493), .A2(n_577), .A3(n_581), .B1(n_582), .B2(n_586), .B3(n_589), .C1(n_590), .C2(n_592), .Y(n_576) );
NAND2x1_ASAP7_75t_L g661 ( .A(n_493), .B(n_552), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_493), .B(n_566), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_SL g594 ( .A1(n_494), .A2(n_595), .B(n_598), .C(n_599), .Y(n_594) );
AND2x2_ASAP7_75t_L g733 ( .A(n_494), .B(n_574), .Y(n_733) );
INVx3_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g630 ( .A(n_495), .B(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g635 ( .A(n_495), .B(n_632), .Y(n_635) );
INVx1_ASAP7_75t_L g566 ( .A(n_496), .Y(n_566) );
AND2x2_ASAP7_75t_L g669 ( .A(n_496), .B(n_628), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_496), .B(n_609), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_496), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_496), .B(n_587), .Y(n_695) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx3_ASAP7_75t_L g552 ( .A(n_497), .Y(n_552) );
OAI31xp33_ASAP7_75t_L g734 ( .A1(n_507), .A2(n_655), .A3(n_662), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_518), .Y(n_507) );
AND2x2_ASAP7_75t_L g539 ( .A(n_508), .B(n_540), .Y(n_539) );
NAND2x1_ASAP7_75t_SL g557 ( .A(n_508), .B(n_558), .Y(n_557) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_508), .Y(n_644) );
AND2x2_ASAP7_75t_L g649 ( .A(n_508), .B(n_560), .Y(n_649) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_509), .A2(n_562), .B(n_564), .C(n_567), .Y(n_561) );
OR2x2_ASAP7_75t_L g578 ( .A(n_509), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g591 ( .A(n_509), .Y(n_591) );
AND2x2_ASAP7_75t_L g597 ( .A(n_509), .B(n_541), .Y(n_597) );
INVx2_ASAP7_75t_L g615 ( .A(n_509), .Y(n_615) );
AND2x2_ASAP7_75t_L g626 ( .A(n_509), .B(n_580), .Y(n_626) );
AND2x2_ASAP7_75t_L g658 ( .A(n_509), .B(n_616), .Y(n_658) );
AND2x2_ASAP7_75t_L g662 ( .A(n_509), .B(n_585), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_509), .B(n_518), .Y(n_667) );
AND2x2_ASAP7_75t_L g701 ( .A(n_509), .B(n_702), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_509), .B(n_604), .Y(n_735) );
OR2x6_ASAP7_75t_L g509 ( .A(n_510), .B(n_516), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_518), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g643 ( .A(n_518), .Y(n_643) );
AND2x2_ASAP7_75t_L g705 ( .A(n_518), .B(n_626), .Y(n_705) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .Y(n_518) );
OR2x2_ASAP7_75t_L g559 ( .A(n_519), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g569 ( .A(n_519), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_519), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g677 ( .A(n_519), .Y(n_677) );
AND2x2_ASAP7_75t_L g694 ( .A(n_519), .B(n_541), .Y(n_694) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g585 ( .A(n_520), .B(n_530), .Y(n_585) );
AND2x2_ASAP7_75t_L g614 ( .A(n_520), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g625 ( .A(n_520), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_520), .B(n_580), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_526), .Y(n_523) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g540 ( .A(n_531), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g560 ( .A(n_531), .Y(n_560) );
AND2x2_ASAP7_75t_L g616 ( .A(n_531), .B(n_580), .Y(n_616) );
INVx1_ASAP7_75t_L g718 ( .A(n_539), .Y(n_718) );
INVx1_ASAP7_75t_L g722 ( .A(n_540), .Y(n_722) );
INVx2_ASAP7_75t_L g580 ( .A(n_541), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_551), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_551), .B(n_656), .Y(n_714) );
OR2x2_ASAP7_75t_L g555 ( .A(n_552), .B(n_553), .Y(n_555) );
INVx1_ASAP7_75t_SL g607 ( .A(n_552), .Y(n_607) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_558), .A2(n_611), .B1(n_613), .B2(n_617), .C(n_618), .Y(n_610) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g638 ( .A(n_559), .B(n_602), .Y(n_638) );
INVx2_ASAP7_75t_L g570 ( .A(n_560), .Y(n_570) );
INVx1_ASAP7_75t_L g596 ( .A(n_560), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_560), .B(n_580), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_560), .B(n_583), .Y(n_690) );
INVx1_ASAP7_75t_L g698 ( .A(n_560), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_562), .B(n_566), .Y(n_612) );
AND2x4_ASAP7_75t_L g587 ( .A(n_563), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g700 ( .A(n_566), .B(n_656), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_569), .B(n_601), .Y(n_600) );
INVxp67_ASAP7_75t_L g708 ( .A(n_570), .Y(n_708) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g608 ( .A(n_574), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g680 ( .A(n_574), .B(n_656), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_574), .B(n_593), .Y(n_686) );
AOI322xp5_ASAP7_75t_L g640 ( .A1(n_575), .A2(n_609), .A3(n_616), .B1(n_641), .B2(n_644), .C1(n_645), .C2(n_647), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_575), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g706 ( .A(n_578), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g652 ( .A(n_579), .Y(n_652) );
INVx2_ASAP7_75t_L g583 ( .A(n_580), .Y(n_583) );
INVx1_ASAP7_75t_L g642 ( .A(n_580), .Y(n_642) );
CKINVDCx16_ASAP7_75t_R g589 ( .A(n_581), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AND2x2_ASAP7_75t_L g678 ( .A(n_583), .B(n_591), .Y(n_678) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g590 ( .A(n_585), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g633 ( .A(n_585), .B(n_626), .Y(n_633) );
AND2x2_ASAP7_75t_L g637 ( .A(n_585), .B(n_597), .Y(n_637) );
OAI21xp33_ASAP7_75t_SL g647 ( .A1(n_586), .A2(n_648), .B(n_650), .Y(n_647) );
OAI22xp33_ASAP7_75t_L g717 ( .A1(n_586), .A2(n_718), .B1(n_719), .B2(n_721), .Y(n_717) );
INVx3_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g592 ( .A(n_587), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_587), .B(n_607), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_589), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g729 ( .A(n_596), .Y(n_729) );
INVx4_ASAP7_75t_L g602 ( .A(n_597), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_597), .B(n_624), .Y(n_672) );
INVx1_ASAP7_75t_SL g684 ( .A(n_598), .Y(n_684) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NOR2xp67_ASAP7_75t_L g697 ( .A(n_602), .B(n_698), .Y(n_697) );
OAI211xp5_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_605), .B(n_610), .C(n_627), .Y(n_603) );
OAI221xp5_ASAP7_75t_SL g723 ( .A1(n_605), .A2(n_643), .B1(n_722), .B2(n_724), .C(n_726), .Y(n_723) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_607), .B(n_720), .Y(n_719) );
OAI31xp33_ASAP7_75t_L g699 ( .A1(n_608), .A2(n_685), .A3(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g639 ( .A(n_609), .Y(n_639) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g689 ( .A(n_614), .Y(n_689) );
AND2x2_ASAP7_75t_L g702 ( .A(n_616), .B(n_625), .Y(n_702) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B(n_622), .Y(n_618) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_626), .B(n_729), .Y(n_728) );
OAI21xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B(n_633), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI221xp5_ASAP7_75t_SL g634 ( .A1(n_635), .A2(n_636), .B1(n_638), .B2(n_639), .C(n_640), .Y(n_634) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_635), .A2(n_704), .B(n_706), .C(n_709), .Y(n_703) );
CKINVDCx16_ASAP7_75t_R g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_638), .B(n_688), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx1_ASAP7_75t_L g665 ( .A(n_646), .Y(n_665) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g651 ( .A(n_649), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g693 ( .A(n_649), .B(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI211xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_657), .B(n_659), .C(n_668), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI221xp5_ASAP7_75t_L g730 ( .A1(n_657), .A2(n_667), .B1(n_731), .B2(n_732), .C(n_734), .Y(n_730) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_662), .B1(n_663), .B2(n_666), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OAI21xp5_ASAP7_75t_SL g668 ( .A1(n_669), .A2(n_670), .B(n_671), .Y(n_668) );
INVx1_ASAP7_75t_SL g731 ( .A(n_670), .Y(n_731) );
INVxp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NOR4xp25_ASAP7_75t_L g673 ( .A(n_674), .B(n_703), .C(n_723), .D(n_730), .Y(n_673) );
OAI211xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_679), .B(n_681), .C(n_699), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVxp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_685), .B(n_687), .C(n_691), .Y(n_681) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g710 ( .A(n_688), .Y(n_710) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
OR2x2_ASAP7_75t_L g721 ( .A(n_689), .B(n_722), .Y(n_721) );
OAI21xp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_695), .B(n_696), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B1(n_713), .B2(n_715), .C(n_717), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_720), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
NAND2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
endmodule