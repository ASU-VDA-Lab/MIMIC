module fake_jpeg_23561_n_137 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_SL g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_30),
.B(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_35),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_22),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_55),
.Y(n_71)
);

CKINVDCx12_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_52),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_26),
.B1(n_18),
.B2(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_48),
.B1(n_53),
.B2(n_16),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_26),
.B1(n_18),
.B2(n_24),
.Y(n_48)
);

AND2x6_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_2),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_56),
.C(n_10),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_15),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_2),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_31),
.B1(n_22),
.B2(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_22),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_16),
.C(n_8),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_34),
.A2(n_29),
.B1(n_27),
.B2(n_30),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_17),
.B2(n_23),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_34),
.A2(n_29),
.B1(n_27),
.B2(n_22),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_66),
.B1(n_51),
.B2(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_68),
.Y(n_91)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_20),
.B1(n_14),
.B2(n_13),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_35),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_20),
.B(n_14),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_12),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_12),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_76),
.Y(n_78)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_76),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_46),
.C(n_48),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_90),
.C(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_90),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_49),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_72),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_75),
.B(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_41),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_94),
.C(n_86),
.Y(n_110)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_95),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_61),
.C(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_103),
.B1(n_89),
.B2(n_79),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_74),
.C(n_72),
.Y(n_98)
);

BUFx12f_ASAP7_75t_SL g108 ( 
.A(n_98),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_102),
.B1(n_87),
.B2(n_77),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_41),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_88),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_104),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_109),
.A2(n_111),
.B1(n_93),
.B2(n_94),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_84),
.C(n_11),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_83),
.B1(n_84),
.B2(n_63),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_113),
.B(n_114),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_99),
.B(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_116),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_10),
.C(n_4),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_124),
.B(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_112),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_110),
.C(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_126),
.B(n_127),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_129),
.A2(n_5),
.B1(n_7),
.B2(n_128),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_3),
.B(n_4),
.Y(n_130)
);

OAI21x1_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_3),
.B(n_4),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_129),
.C(n_7),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_132),
.C(n_7),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_136),
.B(n_135),
.CI(n_131),
.CON(n_137),
.SN(n_137)
);


endmodule