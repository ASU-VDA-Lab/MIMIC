module fake_jpeg_12782_n_45 (n_3, n_2, n_1, n_0, n_4, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_1),
.B(n_0),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_19),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx3_ASAP7_75t_SL g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_SL g20 ( 
.A1(n_9),
.A2(n_6),
.B(n_14),
.C(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_13),
.A2(n_0),
.B(n_5),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_5),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_7),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_12),
.B1(n_8),
.B2(n_11),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_32),
.B(n_23),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_21),
.B(n_20),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_31),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_17),
.B(n_10),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_30),
.C(n_18),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_38),
.B1(n_27),
.B2(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_37),
.C(n_30),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_42),
.B(n_27),
.Y(n_45)
);


endmodule