module fake_jpeg_678_n_359 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_359);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_359;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_51),
.B(n_54),
.Y(n_111)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_52),
.Y(n_130)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_6),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_59),
.Y(n_103)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_57),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_18),
.B(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_61),
.B(n_64),
.Y(n_112)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_19),
.Y(n_65)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_21),
.B(n_4),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_84),
.Y(n_115)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_42),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_SL g131 ( 
.A1(n_72),
.A2(n_37),
.B(n_36),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_80),
.Y(n_121)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_77),
.Y(n_135)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_22),
.B(n_4),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g123 ( 
.A(n_82),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_26),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_26),
.B(n_4),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_90),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

BUFx2_ASAP7_75t_SL g116 ( 
.A(n_89),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_27),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_93),
.Y(n_114)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_3),
.C(n_7),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_96),
.Y(n_137)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_27),
.B(n_3),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_28),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_100),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_28),
.B(n_7),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_31),
.B(n_8),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_101),
.B(n_1),
.Y(n_159)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_102),
.B(n_0),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_23),
.B1(n_39),
.B2(n_30),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_104),
.B(n_138),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_69),
.A2(n_45),
.B1(n_25),
.B2(n_37),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_118),
.A2(n_120),
.B1(n_122),
.B2(n_127),
.Y(n_163)
);

OR2x2_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_97),
.Y(n_119)
);

OR2x2_ASAP7_75t_SL g203 ( 
.A(n_119),
.B(n_131),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_31),
.B1(n_46),
.B2(n_41),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_41),
.B1(n_46),
.B2(n_38),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_34),
.B1(n_30),
.B2(n_43),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_50),
.A2(n_35),
.B1(n_43),
.B2(n_39),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_128),
.A2(n_140),
.B1(n_141),
.B2(n_150),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_76),
.A2(n_45),
.B1(n_25),
.B2(n_38),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_55),
.A2(n_45),
.B1(n_25),
.B2(n_35),
.Y(n_141)
);

BUFx12f_ASAP7_75t_SL g142 ( 
.A(n_86),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g200 ( 
.A(n_142),
.B(n_159),
.C(n_116),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_58),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_149),
.B(n_83),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_68),
.A2(n_34),
.B1(n_23),
.B2(n_36),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_74),
.A2(n_49),
.B1(n_8),
.B2(n_10),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_2),
.B1(n_49),
.B2(n_89),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_95),
.A2(n_8),
.B1(n_10),
.B2(n_49),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_156),
.A2(n_160),
.B1(n_65),
.B2(n_53),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_52),
.A2(n_2),
.B1(n_49),
.B2(n_67),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_161),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_165),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_114),
.A2(n_73),
.B1(n_92),
.B2(n_71),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_166),
.A2(n_193),
.B1(n_132),
.B2(n_130),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_167),
.A2(n_175),
.B1(n_176),
.B2(n_192),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_79),
.C(n_88),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_150),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_172),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_111),
.B(n_78),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_177),
.Y(n_212)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_174),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_147),
.A2(n_81),
.B1(n_77),
.B2(n_62),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_114),
.A2(n_57),
.B1(n_91),
.B2(n_63),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_178),
.B(n_182),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_115),
.B(n_2),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_180),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_144),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_185),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_123),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_183),
.A2(n_135),
.B1(n_155),
.B2(n_132),
.Y(n_216)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_112),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_187),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_189),
.Y(n_234)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_191),
.Y(n_210)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_125),
.A2(n_86),
.B1(n_99),
.B2(n_2),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_148),
.B1(n_136),
.B2(n_141),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_133),
.B(n_137),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_194),
.B(n_195),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_121),
.B(n_103),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_125),
.B(n_105),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_124),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_200),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_145),
.B(n_108),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_202),
.Y(n_215)
);

INVx6_ASAP7_75t_SL g202 ( 
.A(n_142),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_205),
.B(n_213),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_118),
.B1(n_140),
.B2(n_158),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_208),
.B(n_224),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_203),
.A2(n_158),
.B(n_107),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_223),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_151),
.B(n_130),
.C(n_129),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_197),
.A2(n_106),
.B1(n_129),
.B2(n_117),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_190),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_168),
.A2(n_117),
.B(n_106),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_213),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_186),
.A2(n_193),
.B1(n_202),
.B2(n_163),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_235),
.B1(n_191),
.B2(n_184),
.Y(n_242)
);

AND2x6_ASAP7_75t_L g232 ( 
.A(n_180),
.B(n_166),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_174),
.Y(n_238)
);

AOI22x1_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_185),
.B1(n_171),
.B2(n_199),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_179),
.C(n_161),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_248),
.C(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_254),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_164),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_239),
.B(n_240),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_181),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_258),
.B1(n_260),
.B2(n_224),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_219),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_243),
.B(n_244),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_209),
.B(n_188),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_204),
.B(n_177),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_247),
.B(n_257),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_170),
.C(n_165),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_250),
.B(n_251),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_209),
.B(n_162),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_234),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_255),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_207),
.B(n_177),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_259),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_207),
.B(n_211),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_212),
.B(n_215),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_254),
.A2(n_232),
.B1(n_223),
.B2(n_211),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_262),
.B(n_263),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_214),
.B(n_227),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_268),
.A2(n_270),
.B(n_281),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_246),
.B(n_242),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_246),
.A2(n_252),
.B1(n_259),
.B2(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_272),
.A2(n_275),
.B1(n_278),
.B2(n_249),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_252),
.A2(n_215),
.B1(n_214),
.B2(n_220),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_252),
.A2(n_218),
.B1(n_220),
.B2(n_216),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_210),
.B(n_226),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_210),
.C(n_234),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_253),
.C(n_248),
.Y(n_292)
);

AO22x1_ASAP7_75t_L g283 ( 
.A1(n_241),
.A2(n_228),
.B1(n_229),
.B2(n_222),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_228),
.B(n_236),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_265),
.Y(n_285)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_264),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_295),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_270),
.A2(n_255),
.B1(n_237),
.B2(n_250),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_288),
.A2(n_272),
.B1(n_262),
.B2(n_266),
.Y(n_312)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_289),
.A2(n_291),
.B(n_299),
.Y(n_308)
);

BUFx12f_ASAP7_75t_SL g290 ( 
.A(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_290),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_275),
.A2(n_244),
.B1(n_251),
.B2(n_245),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_294),
.C(n_267),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_269),
.B(n_243),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_293),
.B(n_300),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_269),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_298),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_277),
.B(n_218),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_281),
.B(n_271),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_309),
.B(n_311),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_316),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_294),
.B(n_282),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_315),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_273),
.C(n_271),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_273),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_268),
.B(n_263),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_284),
.Y(n_322)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_318),
.A2(n_319),
.B1(n_326),
.B2(n_327),
.Y(n_333)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_306),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_303),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_320),
.B(n_323),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_308),
.Y(n_337)
);

AO221x1_ASAP7_75t_L g323 ( 
.A1(n_312),
.A2(n_290),
.B1(n_285),
.B2(n_287),
.C(n_293),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_307),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_325),
.B(n_314),
.Y(n_335)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_305),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_304),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_315),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_331),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_318),
.A2(n_319),
.B1(n_301),
.B2(n_289),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_309),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_335),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_322),
.A2(n_301),
.B1(n_317),
.B2(n_310),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_334),
.A2(n_295),
.B1(n_286),
.B2(n_291),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_327),
.B(n_313),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_336),
.B(n_337),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_328),
.C(n_321),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_339),
.C(n_311),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_313),
.C(n_316),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_341),
.A2(n_334),
.B1(n_331),
.B2(n_333),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_340),
.A2(n_330),
.B(n_337),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_344),
.B(n_347),
.C(n_348),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_342),
.A2(n_308),
.B(n_326),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_345),
.A2(n_300),
.B(n_297),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_346),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_302),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_348),
.B(n_338),
.C(n_299),
.Y(n_350)
);

AOI31xp33_ASAP7_75t_L g353 ( 
.A1(n_350),
.A2(n_352),
.A3(n_296),
.B(n_279),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_353),
.B(n_354),
.Y(n_356)
);

AOI322xp5_ASAP7_75t_L g354 ( 
.A1(n_351),
.A2(n_278),
.A3(n_279),
.B1(n_222),
.B2(n_225),
.C1(n_206),
.C2(n_229),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_353),
.B(n_349),
.C(n_225),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_355),
.B(n_206),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_357),
.B(n_356),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_217),
.Y(n_359)
);


endmodule