module fake_ariane_1878_n_5359 (n_913, n_589, n_1174, n_691, n_423, n_603, n_373, n_1250, n_1169, n_789, n_850, n_610, n_245, n_96, n_319, n_49, n_690, n_416, n_1109, n_525, n_187, n_1238, n_817, n_924, n_781, n_189, n_717, n_72, n_952, n_864, n_1096, n_57, n_117, n_524, n_1214, n_634, n_1246, n_1138, n_214, n_764, n_462, n_1196, n_1181, n_32, n_410, n_1187, n_1131, n_1225, n_737, n_137, n_232, n_52, n_568, n_1088, n_77, n_766, n_377, n_520, n_870, n_279, n_945, n_958, n_813, n_419, n_146, n_270, n_338, n_995, n_285, n_1184, n_202, n_500, n_665, n_754, n_903, n_871, n_1073, n_239, n_402, n_1277, n_54, n_829, n_1062, n_339, n_738, n_672, n_740, n_1283, n_167, n_1018, n_69, n_259, n_953, n_143, n_1224, n_625, n_557, n_1107, n_989, n_242, n_645, n_331, n_559, n_267, n_495, n_350, n_381, n_795, n_721, n_1084, n_1276, n_200, n_1284, n_1241, n_821, n_561, n_770, n_507, n_486, n_901, n_569, n_1145, n_971, n_787, n_31, n_1195, n_518, n_1207, n_222, n_786, n_868, n_884, n_1034, n_1085, n_277, n_432, n_293, n_823, n_620, n_93, n_1074, n_859, n_108, n_587, n_693, n_863, n_303, n_1254, n_929, n_206, n_352, n_899, n_611, n_238, n_365, n_1013, n_136, n_334, n_192, n_661, n_300, n_533, n_104, n_438, n_16, n_440, n_273, n_1230, n_612, n_333, n_376, n_512, n_579, n_844, n_1012, n_1267, n_149, n_1213, n_237, n_780, n_1021, n_491, n_1142, n_1140, n_705, n_570, n_260, n_942, n_7, n_461, n_1121, n_209, n_490, n_17, n_225, n_1006, n_575, n_546, n_503, n_1112, n_700, n_1159, n_772, n_1216, n_1245, n_676, n_42, n_680, n_287, n_302, n_380, n_94, n_4, n_249, n_1108, n_355, n_212, n_65, n_123, n_444, n_851, n_1274, n_257, n_652, n_475, n_135, n_947, n_930, n_1260, n_1179, n_468, n_102, n_182, n_696, n_482, n_798, n_577, n_407, n_27, n_916, n_912, n_460, n_366, n_762, n_1253, n_555, n_804, n_966, n_992, n_955, n_1182, n_794, n_78, n_514, n_418, n_513, n_288, n_179, n_1292, n_1178, n_1026, n_306, n_92, n_203, n_436, n_150, n_324, n_669, n_931, n_619, n_337, n_437, n_111, n_21, n_274, n_967, n_1083, n_746, n_292, n_1079, n_615, n_1139, n_76, n_517, n_0, n_824, n_428, n_159, n_892, n_959, n_30, n_1101, n_563, n_144, n_990, n_867, n_1226, n_944, n_749, n_815, n_542, n_470, n_1240, n_1087, n_632, n_477, n_650, n_425, n_1155, n_1071, n_712, n_976, n_909, n_767, n_964, n_382, n_489, n_80, n_251, n_974, n_506, n_799, n_1147, n_397, n_471, n_351, n_965, n_155, n_934, n_1220, n_356, n_698, n_124, n_307, n_1209, n_1020, n_646, n_34, n_404, n_172, n_1058, n_347, n_1042, n_183, n_1234, n_479, n_299, n_836, n_1279, n_564, n_133, n_66, n_205, n_1029, n_1247, n_760, n_522, n_20, n_367, n_1111, n_970, n_713, n_1255, n_598, n_345, n_1237, n_927, n_261, n_1095, n_370, n_706, n_286, n_776, n_424, n_85, n_130, n_466, n_1263, n_346, n_348, n_552, n_670, n_379, n_138, n_162, n_264, n_441, n_1032, n_1217, n_637, n_73, n_327, n_1259, n_1177, n_1231, n_980, n_905, n_207, n_720, n_926, n_41, n_194, n_1163, n_186, n_145, n_59, n_1173, n_1068, n_1198, n_487, n_90, n_855, n_158, n_808, n_553, n_814, n_578, n_1287, n_405, n_120, n_320, n_1134, n_647, n_481, n_600, n_1053, n_529, n_502, n_218, n_247, n_1105, n_547, n_439, n_604, n_677, n_478, n_703, n_1061, n_326, n_681, n_227, n_874, n_1278, n_707, n_11, n_129, n_126, n_983, n_590, n_699, n_727, n_301, n_545, n_1015, n_1162, n_536, n_325, n_688, n_636, n_427, n_1098, n_442, n_777, n_1080, n_920, n_1086, n_1092, n_986, n_1104, n_729, n_887, n_1122, n_1205, n_163, n_1132, n_390, n_1156, n_501, n_314, n_1120, n_1202, n_627, n_1188, n_233, n_957, n_388, n_1242, n_1218, n_221, n_321, n_86, n_861, n_877, n_1119, n_616, n_1055, n_1189, n_1089, n_281, n_262, n_735, n_297, n_1005, n_527, n_46, n_84, n_845, n_888, n_178, n_551, n_417, n_70, n_343, n_1222, n_582, n_755, n_1097, n_1219, n_710, n_534, n_1239, n_278, n_560, n_890, n_842, n_148, n_451, n_745, n_61, n_742, n_1081, n_1266, n_769, n_13, n_476, n_832, n_55, n_535, n_744, n_982, n_915, n_215, n_1075, n_454, n_298, n_1227, n_655, n_403, n_1007, n_657, n_837, n_812, n_606, n_951, n_862, n_659, n_509, n_666, n_430, n_1206, n_722, n_1171, n_1030, n_785, n_999, n_456, n_852, n_704, n_1060, n_1044, n_521, n_873, n_1243, n_342, n_358, n_608, n_1037, n_317, n_134, n_1257, n_1078, n_266, n_157, n_1161, n_811, n_624, n_791, n_876, n_618, n_1191, n_736, n_1025, n_1215, n_241, n_687, n_797, n_480, n_211, n_642, n_97, n_408, n_595, n_602, n_592, n_854, n_393, n_474, n_805, n_295, n_190, n_1072, n_695, n_64, n_180, n_730, n_386, n_1281, n_516, n_1137, n_1258, n_197, n_640, n_463, n_943, n_1118, n_678, n_651, n_1293, n_961, n_469, n_1046, n_726, n_1123, n_878, n_771, n_752, n_71, n_985, n_421, n_906, n_1180, n_283, n_806, n_649, n_374, n_643, n_226, n_682, n_36, n_819, n_586, n_686, n_605, n_1154, n_584, n_1130, n_349, n_756, n_1016, n_1149, n_979, n_2, n_897, n_949, n_515, n_807, n_891, n_885, n_198, n_1208, n_396, n_802, n_23, n_1151, n_554, n_960, n_1256, n_87, n_714, n_790, n_354, n_140, n_725, n_151, n_28, n_1009, n_230, n_1133, n_154, n_883, n_142, n_473, n_801, n_1286, n_818, n_779, n_594, n_35, n_1052, n_272, n_833, n_879, n_1117, n_38, n_422, n_1269, n_597, n_75, n_1047, n_95, n_1050, n_566, n_152, n_169, n_106, n_1201, n_1288, n_173, n_858, n_1185, n_335, n_1035, n_1143, n_344, n_426, n_433, n_398, n_62, n_210, n_1090, n_166, n_253, n_928, n_1153, n_271, n_465, n_825, n_1103, n_732, n_1192, n_128, n_224, n_82, n_894, n_420, n_1291, n_562, n_748, n_510, n_1045, n_256, n_1160, n_1023, n_988, n_330, n_914, n_400, n_689, n_1116, n_282, n_328, n_368, n_467, n_644, n_1197, n_276, n_497, n_1165, n_168, n_81, n_538, n_576, n_843, n_511, n_455, n_429, n_588, n_638, n_1128, n_1048, n_775, n_667, n_1049, n_14, n_869, n_141, n_846, n_305, n_312, n_56, n_60, n_728, n_413, n_715, n_889, n_1066, n_935, n_685, n_911, n_361, n_89, n_623, n_1065, n_453, n_74, n_810, n_19, n_40, n_1290, n_181, n_617, n_543, n_236, n_601, n_683, n_565, n_628, n_743, n_1194, n_907, n_660, n_464, n_962, n_941, n_1210, n_847, n_747, n_1135, n_918, n_107, n_639, n_452, n_673, n_1038, n_414, n_571, n_6, n_284, n_593, n_1164, n_37, n_58, n_609, n_1193, n_613, n_1022, n_1033, n_409, n_171, n_519, n_384, n_1166, n_1056, n_526, n_1040, n_674, n_1158, n_316, n_125, n_820, n_43, n_872, n_254, n_1157, n_234, n_848, n_280, n_629, n_161, n_532, n_763, n_99, n_540, n_216, n_692, n_5, n_984, n_223, n_750, n_834, n_800, n_395, n_621, n_213, n_67, n_1014, n_724, n_493, n_114, n_1100, n_585, n_875, n_827, n_697, n_622, n_296, n_880, n_793, n_1175, n_132, n_751, n_1027, n_1070, n_739, n_1028, n_1221, n_530, n_792, n_1262, n_580, n_494, n_434, n_975, n_229, n_394, n_923, n_1124, n_932, n_1183, n_981, n_1110, n_243, n_185, n_1204, n_994, n_973, n_268, n_972, n_164, n_184, n_856, n_1248, n_1176, n_1054, n_508, n_118, n_121, n_353, n_1057, n_191, n_978, n_1011, n_828, n_322, n_558, n_116, n_39, n_653, n_783, n_556, n_1127, n_170, n_160, n_119, n_1008, n_332, n_581, n_294, n_1024, n_830, n_176, n_987, n_936, n_541, n_499, n_788, n_12, n_908, n_1036, n_341, n_1270, n_109, n_1167, n_1272, n_549, n_591, n_969, n_919, n_50, n_318, n_103, n_244, n_679, n_220, n_663, n_443, n_528, n_1200, n_387, n_406, n_826, n_139, n_391, n_940, n_1077, n_607, n_956, n_445, n_765, n_122, n_1268, n_385, n_917, n_1271, n_372, n_15, n_631, n_399, n_1170, n_1261, n_702, n_857, n_898, n_363, n_968, n_1067, n_1235, n_1064, n_633, n_900, n_1282, n_1093, n_1285, n_193, n_733, n_761, n_731, n_336, n_315, n_311, n_8, n_668, n_758, n_1106, n_47, n_153, n_18, n_648, n_784, n_269, n_816, n_835, n_446, n_1076, n_753, n_701, n_1003, n_1125, n_309, n_115, n_401, n_485, n_504, n_483, n_435, n_1141, n_291, n_822, n_1094, n_840, n_1099, n_839, n_79, n_3, n_759, n_567, n_91, n_240, n_369, n_44, n_1172, n_614, n_1212, n_831, n_778, n_48, n_188, n_323, n_550, n_997, n_635, n_694, n_1113, n_248, n_1152, n_921, n_1236, n_228, n_1265, n_671, n_1, n_1148, n_654, n_1275, n_488, n_904, n_505, n_88, n_498, n_1059, n_684, n_1039, n_539, n_1150, n_977, n_449, n_392, n_1289, n_459, n_1136, n_458, n_1190, n_1144, n_383, n_838, n_175, n_950, n_1017, n_711, n_734, n_723, n_658, n_630, n_53, n_362, n_310, n_709, n_24, n_809, n_235, n_881, n_1019, n_662, n_641, n_910, n_290, n_741, n_939, n_371, n_199, n_217, n_1114, n_708, n_308, n_1223, n_201, n_572, n_1199, n_865, n_10, n_1273, n_1041, n_993, n_948, n_922, n_1004, n_448, n_860, n_1043, n_255, n_450, n_896, n_902, n_1031, n_853, n_716, n_196, n_774, n_933, n_596, n_954, n_1168, n_219, n_231, n_656, n_492, n_574, n_252, n_664, n_1229, n_68, n_415, n_63, n_1280, n_544, n_1186, n_599, n_768, n_1091, n_537, n_1063, n_25, n_991, n_83, n_389, n_1126, n_195, n_938, n_895, n_110, n_304, n_583, n_1000, n_313, n_626, n_378, n_98, n_946, n_757, n_375, n_113, n_33, n_1146, n_1203, n_998, n_472, n_937, n_265, n_208, n_156, n_174, n_275, n_100, n_147, n_204, n_1232, n_996, n_1211, n_963, n_1264, n_51, n_1082, n_496, n_866, n_26, n_246, n_925, n_1001, n_1115, n_1002, n_105, n_1051, n_719, n_131, n_263, n_1102, n_360, n_1129, n_1252, n_250, n_773, n_165, n_1010, n_882, n_1249, n_101, n_803, n_329, n_718, n_340, n_289, n_9, n_112, n_45, n_548, n_523, n_457, n_177, n_782, n_364, n_258, n_431, n_1228, n_1244, n_411, n_484, n_849, n_22, n_29, n_357, n_412, n_1251, n_447, n_1233, n_893, n_841, n_886, n_1069, n_359, n_573, n_796, n_127, n_531, n_675, n_5359);

input n_913;
input n_589;
input n_1174;
input n_691;
input n_423;
input n_603;
input n_373;
input n_1250;
input n_1169;
input n_789;
input n_850;
input n_610;
input n_245;
input n_96;
input n_319;
input n_49;
input n_690;
input n_416;
input n_1109;
input n_525;
input n_187;
input n_1238;
input n_817;
input n_924;
input n_781;
input n_189;
input n_717;
input n_72;
input n_952;
input n_864;
input n_1096;
input n_57;
input n_117;
input n_524;
input n_1214;
input n_634;
input n_1246;
input n_1138;
input n_214;
input n_764;
input n_462;
input n_1196;
input n_1181;
input n_32;
input n_410;
input n_1187;
input n_1131;
input n_1225;
input n_737;
input n_137;
input n_232;
input n_52;
input n_568;
input n_1088;
input n_77;
input n_766;
input n_377;
input n_520;
input n_870;
input n_279;
input n_945;
input n_958;
input n_813;
input n_419;
input n_146;
input n_270;
input n_338;
input n_995;
input n_285;
input n_1184;
input n_202;
input n_500;
input n_665;
input n_754;
input n_903;
input n_871;
input n_1073;
input n_239;
input n_402;
input n_1277;
input n_54;
input n_829;
input n_1062;
input n_339;
input n_738;
input n_672;
input n_740;
input n_1283;
input n_167;
input n_1018;
input n_69;
input n_259;
input n_953;
input n_143;
input n_1224;
input n_625;
input n_557;
input n_1107;
input n_989;
input n_242;
input n_645;
input n_331;
input n_559;
input n_267;
input n_495;
input n_350;
input n_381;
input n_795;
input n_721;
input n_1084;
input n_1276;
input n_200;
input n_1284;
input n_1241;
input n_821;
input n_561;
input n_770;
input n_507;
input n_486;
input n_901;
input n_569;
input n_1145;
input n_971;
input n_787;
input n_31;
input n_1195;
input n_518;
input n_1207;
input n_222;
input n_786;
input n_868;
input n_884;
input n_1034;
input n_1085;
input n_277;
input n_432;
input n_293;
input n_823;
input n_620;
input n_93;
input n_1074;
input n_859;
input n_108;
input n_587;
input n_693;
input n_863;
input n_303;
input n_1254;
input n_929;
input n_206;
input n_352;
input n_899;
input n_611;
input n_238;
input n_365;
input n_1013;
input n_136;
input n_334;
input n_192;
input n_661;
input n_300;
input n_533;
input n_104;
input n_438;
input n_16;
input n_440;
input n_273;
input n_1230;
input n_612;
input n_333;
input n_376;
input n_512;
input n_579;
input n_844;
input n_1012;
input n_1267;
input n_149;
input n_1213;
input n_237;
input n_780;
input n_1021;
input n_491;
input n_1142;
input n_1140;
input n_705;
input n_570;
input n_260;
input n_942;
input n_7;
input n_461;
input n_1121;
input n_209;
input n_490;
input n_17;
input n_225;
input n_1006;
input n_575;
input n_546;
input n_503;
input n_1112;
input n_700;
input n_1159;
input n_772;
input n_1216;
input n_1245;
input n_676;
input n_42;
input n_680;
input n_287;
input n_302;
input n_380;
input n_94;
input n_4;
input n_249;
input n_1108;
input n_355;
input n_212;
input n_65;
input n_123;
input n_444;
input n_851;
input n_1274;
input n_257;
input n_652;
input n_475;
input n_135;
input n_947;
input n_930;
input n_1260;
input n_1179;
input n_468;
input n_102;
input n_182;
input n_696;
input n_482;
input n_798;
input n_577;
input n_407;
input n_27;
input n_916;
input n_912;
input n_460;
input n_366;
input n_762;
input n_1253;
input n_555;
input n_804;
input n_966;
input n_992;
input n_955;
input n_1182;
input n_794;
input n_78;
input n_514;
input n_418;
input n_513;
input n_288;
input n_179;
input n_1292;
input n_1178;
input n_1026;
input n_306;
input n_92;
input n_203;
input n_436;
input n_150;
input n_324;
input n_669;
input n_931;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_967;
input n_1083;
input n_746;
input n_292;
input n_1079;
input n_615;
input n_1139;
input n_76;
input n_517;
input n_0;
input n_824;
input n_428;
input n_159;
input n_892;
input n_959;
input n_30;
input n_1101;
input n_563;
input n_144;
input n_990;
input n_867;
input n_1226;
input n_944;
input n_749;
input n_815;
input n_542;
input n_470;
input n_1240;
input n_1087;
input n_632;
input n_477;
input n_650;
input n_425;
input n_1155;
input n_1071;
input n_712;
input n_976;
input n_909;
input n_767;
input n_964;
input n_382;
input n_489;
input n_80;
input n_251;
input n_974;
input n_506;
input n_799;
input n_1147;
input n_397;
input n_471;
input n_351;
input n_965;
input n_155;
input n_934;
input n_1220;
input n_356;
input n_698;
input n_124;
input n_307;
input n_1209;
input n_1020;
input n_646;
input n_34;
input n_404;
input n_172;
input n_1058;
input n_347;
input n_1042;
input n_183;
input n_1234;
input n_479;
input n_299;
input n_836;
input n_1279;
input n_564;
input n_133;
input n_66;
input n_205;
input n_1029;
input n_1247;
input n_760;
input n_522;
input n_20;
input n_367;
input n_1111;
input n_970;
input n_713;
input n_1255;
input n_598;
input n_345;
input n_1237;
input n_927;
input n_261;
input n_1095;
input n_370;
input n_706;
input n_286;
input n_776;
input n_424;
input n_85;
input n_130;
input n_466;
input n_1263;
input n_346;
input n_348;
input n_552;
input n_670;
input n_379;
input n_138;
input n_162;
input n_264;
input n_441;
input n_1032;
input n_1217;
input n_637;
input n_73;
input n_327;
input n_1259;
input n_1177;
input n_1231;
input n_980;
input n_905;
input n_207;
input n_720;
input n_926;
input n_41;
input n_194;
input n_1163;
input n_186;
input n_145;
input n_59;
input n_1173;
input n_1068;
input n_1198;
input n_487;
input n_90;
input n_855;
input n_158;
input n_808;
input n_553;
input n_814;
input n_578;
input n_1287;
input n_405;
input n_120;
input n_320;
input n_1134;
input n_647;
input n_481;
input n_600;
input n_1053;
input n_529;
input n_502;
input n_218;
input n_247;
input n_1105;
input n_547;
input n_439;
input n_604;
input n_677;
input n_478;
input n_703;
input n_1061;
input n_326;
input n_681;
input n_227;
input n_874;
input n_1278;
input n_707;
input n_11;
input n_129;
input n_126;
input n_983;
input n_590;
input n_699;
input n_727;
input n_301;
input n_545;
input n_1015;
input n_1162;
input n_536;
input n_325;
input n_688;
input n_636;
input n_427;
input n_1098;
input n_442;
input n_777;
input n_1080;
input n_920;
input n_1086;
input n_1092;
input n_986;
input n_1104;
input n_729;
input n_887;
input n_1122;
input n_1205;
input n_163;
input n_1132;
input n_390;
input n_1156;
input n_501;
input n_314;
input n_1120;
input n_1202;
input n_627;
input n_1188;
input n_233;
input n_957;
input n_388;
input n_1242;
input n_1218;
input n_221;
input n_321;
input n_86;
input n_861;
input n_877;
input n_1119;
input n_616;
input n_1055;
input n_1189;
input n_1089;
input n_281;
input n_262;
input n_735;
input n_297;
input n_1005;
input n_527;
input n_46;
input n_84;
input n_845;
input n_888;
input n_178;
input n_551;
input n_417;
input n_70;
input n_343;
input n_1222;
input n_582;
input n_755;
input n_1097;
input n_1219;
input n_710;
input n_534;
input n_1239;
input n_278;
input n_560;
input n_890;
input n_842;
input n_148;
input n_451;
input n_745;
input n_61;
input n_742;
input n_1081;
input n_1266;
input n_769;
input n_13;
input n_476;
input n_832;
input n_55;
input n_535;
input n_744;
input n_982;
input n_915;
input n_215;
input n_1075;
input n_454;
input n_298;
input n_1227;
input n_655;
input n_403;
input n_1007;
input n_657;
input n_837;
input n_812;
input n_606;
input n_951;
input n_862;
input n_659;
input n_509;
input n_666;
input n_430;
input n_1206;
input n_722;
input n_1171;
input n_1030;
input n_785;
input n_999;
input n_456;
input n_852;
input n_704;
input n_1060;
input n_1044;
input n_521;
input n_873;
input n_1243;
input n_342;
input n_358;
input n_608;
input n_1037;
input n_317;
input n_134;
input n_1257;
input n_1078;
input n_266;
input n_157;
input n_1161;
input n_811;
input n_624;
input n_791;
input n_876;
input n_618;
input n_1191;
input n_736;
input n_1025;
input n_1215;
input n_241;
input n_687;
input n_797;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_602;
input n_592;
input n_854;
input n_393;
input n_474;
input n_805;
input n_295;
input n_190;
input n_1072;
input n_695;
input n_64;
input n_180;
input n_730;
input n_386;
input n_1281;
input n_516;
input n_1137;
input n_1258;
input n_197;
input n_640;
input n_463;
input n_943;
input n_1118;
input n_678;
input n_651;
input n_1293;
input n_961;
input n_469;
input n_1046;
input n_726;
input n_1123;
input n_878;
input n_771;
input n_752;
input n_71;
input n_985;
input n_421;
input n_906;
input n_1180;
input n_283;
input n_806;
input n_649;
input n_374;
input n_643;
input n_226;
input n_682;
input n_36;
input n_819;
input n_586;
input n_686;
input n_605;
input n_1154;
input n_584;
input n_1130;
input n_349;
input n_756;
input n_1016;
input n_1149;
input n_979;
input n_2;
input n_897;
input n_949;
input n_515;
input n_807;
input n_891;
input n_885;
input n_198;
input n_1208;
input n_396;
input n_802;
input n_23;
input n_1151;
input n_554;
input n_960;
input n_1256;
input n_87;
input n_714;
input n_790;
input n_354;
input n_140;
input n_725;
input n_151;
input n_28;
input n_1009;
input n_230;
input n_1133;
input n_154;
input n_883;
input n_142;
input n_473;
input n_801;
input n_1286;
input n_818;
input n_779;
input n_594;
input n_35;
input n_1052;
input n_272;
input n_833;
input n_879;
input n_1117;
input n_38;
input n_422;
input n_1269;
input n_597;
input n_75;
input n_1047;
input n_95;
input n_1050;
input n_566;
input n_152;
input n_169;
input n_106;
input n_1201;
input n_1288;
input n_173;
input n_858;
input n_1185;
input n_335;
input n_1035;
input n_1143;
input n_344;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_1090;
input n_166;
input n_253;
input n_928;
input n_1153;
input n_271;
input n_465;
input n_825;
input n_1103;
input n_732;
input n_1192;
input n_128;
input n_224;
input n_82;
input n_894;
input n_420;
input n_1291;
input n_562;
input n_748;
input n_510;
input n_1045;
input n_256;
input n_1160;
input n_1023;
input n_988;
input n_330;
input n_914;
input n_400;
input n_689;
input n_1116;
input n_282;
input n_328;
input n_368;
input n_467;
input n_644;
input n_1197;
input n_276;
input n_497;
input n_1165;
input n_168;
input n_81;
input n_538;
input n_576;
input n_843;
input n_511;
input n_455;
input n_429;
input n_588;
input n_638;
input n_1128;
input n_1048;
input n_775;
input n_667;
input n_1049;
input n_14;
input n_869;
input n_141;
input n_846;
input n_305;
input n_312;
input n_56;
input n_60;
input n_728;
input n_413;
input n_715;
input n_889;
input n_1066;
input n_935;
input n_685;
input n_911;
input n_361;
input n_89;
input n_623;
input n_1065;
input n_453;
input n_74;
input n_810;
input n_19;
input n_40;
input n_1290;
input n_181;
input n_617;
input n_543;
input n_236;
input n_601;
input n_683;
input n_565;
input n_628;
input n_743;
input n_1194;
input n_907;
input n_660;
input n_464;
input n_962;
input n_941;
input n_1210;
input n_847;
input n_747;
input n_1135;
input n_918;
input n_107;
input n_639;
input n_452;
input n_673;
input n_1038;
input n_414;
input n_571;
input n_6;
input n_284;
input n_593;
input n_1164;
input n_37;
input n_58;
input n_609;
input n_1193;
input n_613;
input n_1022;
input n_1033;
input n_409;
input n_171;
input n_519;
input n_384;
input n_1166;
input n_1056;
input n_526;
input n_1040;
input n_674;
input n_1158;
input n_316;
input n_125;
input n_820;
input n_43;
input n_872;
input n_254;
input n_1157;
input n_234;
input n_848;
input n_280;
input n_629;
input n_161;
input n_532;
input n_763;
input n_99;
input n_540;
input n_216;
input n_692;
input n_5;
input n_984;
input n_223;
input n_750;
input n_834;
input n_800;
input n_395;
input n_621;
input n_213;
input n_67;
input n_1014;
input n_724;
input n_493;
input n_114;
input n_1100;
input n_585;
input n_875;
input n_827;
input n_697;
input n_622;
input n_296;
input n_880;
input n_793;
input n_1175;
input n_132;
input n_751;
input n_1027;
input n_1070;
input n_739;
input n_1028;
input n_1221;
input n_530;
input n_792;
input n_1262;
input n_580;
input n_494;
input n_434;
input n_975;
input n_229;
input n_394;
input n_923;
input n_1124;
input n_932;
input n_1183;
input n_981;
input n_1110;
input n_243;
input n_185;
input n_1204;
input n_994;
input n_973;
input n_268;
input n_972;
input n_164;
input n_184;
input n_856;
input n_1248;
input n_1176;
input n_1054;
input n_508;
input n_118;
input n_121;
input n_353;
input n_1057;
input n_191;
input n_978;
input n_1011;
input n_828;
input n_322;
input n_558;
input n_116;
input n_39;
input n_653;
input n_783;
input n_556;
input n_1127;
input n_170;
input n_160;
input n_119;
input n_1008;
input n_332;
input n_581;
input n_294;
input n_1024;
input n_830;
input n_176;
input n_987;
input n_936;
input n_541;
input n_499;
input n_788;
input n_12;
input n_908;
input n_1036;
input n_341;
input n_1270;
input n_109;
input n_1167;
input n_1272;
input n_549;
input n_591;
input n_969;
input n_919;
input n_50;
input n_318;
input n_103;
input n_244;
input n_679;
input n_220;
input n_663;
input n_443;
input n_528;
input n_1200;
input n_387;
input n_406;
input n_826;
input n_139;
input n_391;
input n_940;
input n_1077;
input n_607;
input n_956;
input n_445;
input n_765;
input n_122;
input n_1268;
input n_385;
input n_917;
input n_1271;
input n_372;
input n_15;
input n_631;
input n_399;
input n_1170;
input n_1261;
input n_702;
input n_857;
input n_898;
input n_363;
input n_968;
input n_1067;
input n_1235;
input n_1064;
input n_633;
input n_900;
input n_1282;
input n_1093;
input n_1285;
input n_193;
input n_733;
input n_761;
input n_731;
input n_336;
input n_315;
input n_311;
input n_8;
input n_668;
input n_758;
input n_1106;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_816;
input n_835;
input n_446;
input n_1076;
input n_753;
input n_701;
input n_1003;
input n_1125;
input n_309;
input n_115;
input n_401;
input n_485;
input n_504;
input n_483;
input n_435;
input n_1141;
input n_291;
input n_822;
input n_1094;
input n_840;
input n_1099;
input n_839;
input n_79;
input n_3;
input n_759;
input n_567;
input n_91;
input n_240;
input n_369;
input n_44;
input n_1172;
input n_614;
input n_1212;
input n_831;
input n_778;
input n_48;
input n_188;
input n_323;
input n_550;
input n_997;
input n_635;
input n_694;
input n_1113;
input n_248;
input n_1152;
input n_921;
input n_1236;
input n_228;
input n_1265;
input n_671;
input n_1;
input n_1148;
input n_654;
input n_1275;
input n_488;
input n_904;
input n_505;
input n_88;
input n_498;
input n_1059;
input n_684;
input n_1039;
input n_539;
input n_1150;
input n_977;
input n_449;
input n_392;
input n_1289;
input n_459;
input n_1136;
input n_458;
input n_1190;
input n_1144;
input n_383;
input n_838;
input n_175;
input n_950;
input n_1017;
input n_711;
input n_734;
input n_723;
input n_658;
input n_630;
input n_53;
input n_362;
input n_310;
input n_709;
input n_24;
input n_809;
input n_235;
input n_881;
input n_1019;
input n_662;
input n_641;
input n_910;
input n_290;
input n_741;
input n_939;
input n_371;
input n_199;
input n_217;
input n_1114;
input n_708;
input n_308;
input n_1223;
input n_201;
input n_572;
input n_1199;
input n_865;
input n_10;
input n_1273;
input n_1041;
input n_993;
input n_948;
input n_922;
input n_1004;
input n_448;
input n_860;
input n_1043;
input n_255;
input n_450;
input n_896;
input n_902;
input n_1031;
input n_853;
input n_716;
input n_196;
input n_774;
input n_933;
input n_596;
input n_954;
input n_1168;
input n_219;
input n_231;
input n_656;
input n_492;
input n_574;
input n_252;
input n_664;
input n_1229;
input n_68;
input n_415;
input n_63;
input n_1280;
input n_544;
input n_1186;
input n_599;
input n_768;
input n_1091;
input n_537;
input n_1063;
input n_25;
input n_991;
input n_83;
input n_389;
input n_1126;
input n_195;
input n_938;
input n_895;
input n_110;
input n_304;
input n_583;
input n_1000;
input n_313;
input n_626;
input n_378;
input n_98;
input n_946;
input n_757;
input n_375;
input n_113;
input n_33;
input n_1146;
input n_1203;
input n_998;
input n_472;
input n_937;
input n_265;
input n_208;
input n_156;
input n_174;
input n_275;
input n_100;
input n_147;
input n_204;
input n_1232;
input n_996;
input n_1211;
input n_963;
input n_1264;
input n_51;
input n_1082;
input n_496;
input n_866;
input n_26;
input n_246;
input n_925;
input n_1001;
input n_1115;
input n_1002;
input n_105;
input n_1051;
input n_719;
input n_131;
input n_263;
input n_1102;
input n_360;
input n_1129;
input n_1252;
input n_250;
input n_773;
input n_165;
input n_1010;
input n_882;
input n_1249;
input n_101;
input n_803;
input n_329;
input n_718;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_548;
input n_523;
input n_457;
input n_177;
input n_782;
input n_364;
input n_258;
input n_431;
input n_1228;
input n_1244;
input n_411;
input n_484;
input n_849;
input n_22;
input n_29;
input n_357;
input n_412;
input n_1251;
input n_447;
input n_1233;
input n_893;
input n_841;
input n_886;
input n_1069;
input n_359;
input n_573;
input n_796;
input n_127;
input n_531;
input n_675;

output n_5359;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_2182;
wire n_2680;
wire n_3264;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_2729;
wire n_4302;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_5302;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_2646;
wire n_2653;
wire n_4610;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_2482;
wire n_1682;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_4260;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_2322;
wire n_2663;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_1428;
wire n_4741;
wire n_4143;
wire n_4273;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_4567;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_3015;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_3482;
wire n_1900;
wire n_4268;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_5247;
wire n_4476;
wire n_2956;
wire n_5210;
wire n_2382;
wire n_5292;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_3458;
wire n_3511;
wire n_2077;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_3549;
wire n_3914;
wire n_1692;
wire n_2611;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5056;
wire n_2015;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_2257;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5179;
wire n_2435;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_3814;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_2019;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2649;
wire n_1568;
wire n_2919;
wire n_3108;
wire n_2632;
wire n_4314;
wire n_2980;
wire n_1728;
wire n_4315;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_2697;
wire n_1817;
wire n_3704;
wire n_4296;
wire n_2677;
wire n_2483;
wire n_5088;
wire n_1592;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_5149;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_5089;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_5296;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1349;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_4292;
wire n_2118;
wire n_1490;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_3025;
wire n_3051;
wire n_2802;
wire n_2125;
wire n_4974;
wire n_5123;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1498;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_2707;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_3713;
wire n_1863;
wire n_4798;
wire n_1500;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_3944;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_2448;
wire n_2211;
wire n_5318;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_2958;
wire n_1714;
wire n_4429;
wire n_3340;
wire n_5053;
wire n_3486;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_2520;
wire n_3864;
wire n_4694;
wire n_4664;
wire n_3450;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_1406;
wire n_5073;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_2991;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_4822;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_3740;
wire n_2417;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_3726;
wire n_4419;
wire n_3560;
wire n_3345;
wire n_3421;
wire n_1448;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_4966;
wire n_2250;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_3886;
wire n_2619;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_2613;
wire n_1517;
wire n_2647;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_1671;
wire n_5027;
wire n_2343;
wire n_3380;
wire n_2826;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_4631;
wire n_1504;
wire n_2110;
wire n_3822;
wire n_4355;
wire n_3818;
wire n_3587;
wire n_2608;
wire n_1948;
wire n_4155;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_4685;
wire n_3927;
wire n_2068;
wire n_3595;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_3396;
wire n_4093;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_2963;
wire n_2561;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_5125;
wire n_4922;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_3630;
wire n_1612;
wire n_1910;
wire n_2189;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_2931;
wire n_3433;
wire n_3597;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_3786;
wire n_2828;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_3645;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_5011;
wire n_1554;
wire n_3279;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_1679;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_4053;
wire n_3963;
wire n_3091;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_1775;
wire n_4083;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_3225;
wire n_3621;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_3633;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_2009;
wire n_4339;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_3457;
wire n_2324;
wire n_5283;
wire n_3454;
wire n_2139;
wire n_2521;
wire n_2740;
wire n_1991;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_5040;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_3628;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_3872;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_3555;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_4574;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_4663;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_3707;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_5304;
wire n_1581;
wire n_3058;
wire n_2047;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_5355;
wire n_3592;
wire n_5321;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_1368;
wire n_4120;
wire n_2880;
wire n_1313;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_1339;
wire n_5116;
wire n_3771;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_2830;
wire n_4622;
wire n_4757;
wire n_1871;
wire n_4016;
wire n_3334;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_4591;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_2259;
wire n_5337;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_4493;
wire n_1808;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_3181;
wire n_1916;
wire n_4602;
wire n_1713;
wire n_2818;
wire n_1436;
wire n_4900;
wire n_3578;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_1566;
wire n_2837;
wire n_2446;
wire n_4116;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_4439;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_2248;
wire n_4660;
wire n_3081;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_2844;
wire n_1979;
wire n_4814;
wire n_2221;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_2634;
wire n_2746;
wire n_5098;
wire n_5145;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_1528;
wire n_3315;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_5213;
wire n_3474;
wire n_2458;
wire n_3150;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1652;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_2061;
wire n_2685;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_4995;
wire n_4498;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_4850;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_3391;
wire n_4786;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_3240;
wire n_5066;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_5130;
wire n_4175;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_1399;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_3257;
wire n_3730;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_4003;
wire n_1832;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5159;
wire n_4022;
wire n_2495;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_3031;
wire n_2335;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_5287;
wire n_4719;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_2296;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_2059;
wire n_4713;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_4916;
wire n_4323;
wire n_1899;
wire n_3508;
wire n_4129;
wire n_3599;
wire n_4480;
wire n_3734;
wire n_3401;
wire n_3542;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_2218;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_2754;
wire n_4580;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_3995;
wire n_3908;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_2266;
wire n_4324;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_3671;
wire n_2366;
wire n_1753;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_3791;
wire n_2008;
wire n_4989;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_1332;
wire n_1747;
wire n_3990;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5256;
wire n_4779;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_1400;
wire n_3735;
wire n_1513;
wire n_1527;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1954;
wire n_3964;
wire n_3302;
wire n_2486;
wire n_1897;
wire n_2137;
wire n_3685;
wire n_4977;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_2912;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_3411;
wire n_5222;
wire n_3463;
wire n_2785;
wire n_4938;
wire n_2574;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1697;
wire n_2730;
wire n_5129;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_1561;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5161;
wire n_1557;
wire n_4744;
wire n_4706;
wire n_2022;
wire n_3879;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_4990;
wire n_2986;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_3317;
wire n_4835;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_4372;
wire n_4097;
wire n_4162;
wire n_5293;
wire n_4790;
wire n_4173;
wire n_5309;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_3973;
wire n_4799;
wire n_4534;
wire n_4960;
wire n_3738;
wire n_1380;
wire n_2020;
wire n_2310;
wire n_3600;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_3967;
wire n_4370;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_2234;
wire n_1341;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_2592;
wire n_3490;
wire n_5043;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_1968;
wire n_5020;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_4333;
wire n_5339;
wire n_2007;
wire n_3363;
wire n_1803;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_3481;
wire n_5101;
wire n_2236;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_2406;
wire n_4477;
wire n_4110;
wire n_5182;
wire n_4217;
wire n_5277;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_3873;
wire n_4649;
wire n_2428;
wire n_1360;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_4999;
wire n_4592;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_2385;
wire n_1980;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_3114;
wire n_2092;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_1458;
wire n_3047;
wire n_3163;
wire n_1550;
wire n_1358;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_3687;
wire n_2787;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_5193;
wire n_4933;
wire n_4144;
wire n_2375;
wire n_3278;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_4726;
wire n_5143;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_5273;
wire n_2469;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_3068;
wire n_1629;
wire n_1510;
wire n_3002;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_3132;
wire n_5002;
wire n_3681;
wire n_3970;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_4579;
wire n_4776;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_4165;
wire n_2056;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1941;
wire n_3637;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_2917;
wire n_3194;
wire n_2432;
wire n_2085;
wire n_5033;
wire n_1686;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_1410;
wire n_2297;
wire n_4203;
wire n_1325;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_3674;
wire n_1638;
wire n_1571;
wire n_5349;
wire n_3763;
wire n_3499;
wire n_1821;
wire n_3947;
wire n_3910;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_3088;
wire n_1724;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_3075;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_2304;
wire n_2514;
wire n_1299;
wire n_3430;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_4971;
wire n_2095;
wire n_2738;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_2423;
wire n_2208;
wire n_1421;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_2866;
wire n_3153;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_1383;
wire n_4259;
wire n_2030;
wire n_4299;
wire n_2407;
wire n_2243;
wire n_5288;
wire n_2694;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_5294;
wire n_2731;
wire n_3703;
wire n_5265;
wire n_2123;
wire n_2238;
wire n_4802;
wire n_4793;
wire n_3435;
wire n_2380;
wire n_4897;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_3220;
wire n_4581;
wire n_4625;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_5316;
wire n_2735;
wire n_4214;
wire n_1888;
wire n_5290;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_5048;
wire n_2233;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_4032;
wire n_2571;
wire n_4929;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_3634;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_4815;
wire n_4665;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_1461;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_4174;
wire n_5131;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_3119;
wire n_4740;
wire n_4394;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_2628;
wire n_1491;
wire n_3219;
wire n_5333;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_3479;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_2755;
wire n_5109;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_2220;
wire n_4433;
wire n_2829;
wire n_1914;
wire n_2253;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_3936;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_2473;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_3078;
wire n_3971;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_4751;
wire n_4242;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_4952;
wire n_4426;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_2112;
wire n_2640;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_4506;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_4039;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_3983;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_2338;
wire n_5261;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_2660;
wire n_1859;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1711;
wire n_4387;
wire n_3186;
wire n_2508;
wire n_2594;
wire n_5298;
wire n_3417;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_4328;
wire n_1854;
wire n_5191;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_4940;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_2280;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_3586;
wire n_4160;
wire n_1668;
wire n_4137;
wire n_4545;
wire n_4758;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_4535;
wire n_4385;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_4766;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1733;
wire n_4651;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_1352;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_2907;
wire n_2353;
wire n_1429;
wire n_2528;
wire n_1778;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_3718;
wire n_3390;
wire n_2298;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_3976;
wire n_2813;
wire n_2546;
wire n_3381;
wire n_3736;
wire n_4466;
wire n_1659;
wire n_3955;
wire n_5322;
wire n_1864;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_4377;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5270;
wire n_3468;
wire n_1877;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_2497;
wire n_4561;
wire n_3291;
wire n_1541;
wire n_1472;
wire n_2578;
wire n_2475;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5351;
wire n_5267;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_3358;
wire n_2533;
wire n_2003;
wire n_1307;
wire n_4682;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_3289;
wire n_1955;
wire n_1440;
wire n_1370;
wire n_5005;
wire n_1549;
wire n_5207;
wire n_2658;
wire n_3620;
wire n_4601;
wire n_4518;
wire n_2767;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_4711;
wire n_2749;
wire n_4413;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_3723;
wire n_4135;
wire n_5223;
wire n_3880;
wire n_3904;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_3532;
wire n_5154;
wire n_2609;
wire n_1767;
wire n_4138;
wire n_3131;
wire n_1973;
wire n_1444;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_4270;
wire n_4620;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_4406;
wire n_2180;
wire n_4271;
wire n_2809;
wire n_1645;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_2465;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_1834;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_4858;
wire n_1445;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_1663;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_3897;
wire n_1735;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_2186;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_3838;
wire n_4059;
wire n_5194;
wire n_2734;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_3273;
wire n_2918;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3001;
wire n_5260;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_2422;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_1393;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_3032;
wire n_4886;
wire n_5172;
wire n_1477;
wire n_1982;
wire n_5311;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_2982;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_4693;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_4487;
wire n_2674;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_3112;
wire n_2562;
wire n_1779;
wire n_2051;
wire n_3196;
wire n_2673;
wire n_4678;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2179;
wire n_3779;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_1891;
wire n_5348;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_1725;
wire n_2318;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_3045;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_4047;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_2135;
wire n_4475;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_1503;
wire n_5295;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_3383;
wire n_1835;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_2323;
wire n_4549;
wire n_1746;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_1988;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_2078;
wire n_4809;
wire n_4012;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_5042;
wire n_4768;
wire n_1889;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_2727;
wire n_5234;
wire n_1416;
wire n_1599;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_5253;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_5019;
wire n_1819;
wire n_3095;
wire n_3698;
wire n_4513;
wire n_1442;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2499;
wire n_2549;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_4264;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_4170;
wire n_2462;
wire n_2155;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_4267;
wire n_2083;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_2378;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_1483;
wire n_1363;
wire n_3467;
wire n_3179;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_3699;
wire n_2120;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_5335;
wire n_2801;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_3246;
wire n_3299;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_3276;
wire n_3682;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_2932;
wire n_2027;
wire n_3118;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_1467;
wire n_5209;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_5099;
wire n_3286;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_3009;
wire n_5219;
wire n_3951;
wire n_3035;
wire n_4261;
wire n_1823;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_1666;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_3224;
wire n_1969;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_1572;
wire n_4463;
wire n_5357;
wire n_3648;
wire n_1975;
wire n_1388;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_1532;
wire n_5181;
wire n_3208;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_2916;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_3650;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_5017;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_2091;
wire n_4312;
wire n_3789;
wire n_1658;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2725;
wire n_2667;
wire n_3746;
wire n_4537;
wire n_3694;
wire n_3893;
wire n_4847;
wire n_2307;
wire n_3702;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_2945;
wire n_1971;
wire n_3543;
wire n_1324;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_2698;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_5142;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_4595;
wire n_2352;
wire n_5201;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_4054;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_4732;
wire n_2203;
wire n_2076;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_4139;
wire n_4769;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_3509;
wire n_1403;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_3790;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_2174;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_1687;
wire n_4703;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_5228;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_4720;
wire n_2889;
wire n_2141;
wire n_1758;
wire n_3470;
wire n_5221;
wire n_1407;
wire n_2865;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_3677;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_4131;
wire n_4215;
wire n_2488;
wire n_1509;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_2169;
wire n_5133;
wire n_5305;
wire n_2175;
wire n_1625;
wire n_4578;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_2724;
wire n_2258;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_5343;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_2111;
wire n_3743;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_4472;
wire n_2699;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_2710;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_4371;
wire n_1902;
wire n_2784;
wire n_3898;
wire n_4749;
wire n_1845;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_4238;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_3094;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_5034;
wire n_3312;
wire n_2451;
wire n_2913;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_1764;
wire n_4807;
wire n_5115;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_4095;
wire n_1310;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1699;
wire n_5226;
wire n_2081;
wire n_1474;
wire n_1631;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_4516;
wire n_5235;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_1870;
wire n_4467;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_5258;

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1281),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1155),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_518),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_328),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1189),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1108),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_537),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1277),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_41),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1175),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_779),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1182),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_788),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1251),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_749),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_119),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_473),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_228),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1036),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_139),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1003),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_322),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_347),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_534),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_529),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_616),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_89),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1234),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_425),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_330),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1141),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1232),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_830),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_676),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_910),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1008),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_494),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1040),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_903),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_5),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1023),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1026),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_876),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_65),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1148),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_638),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_271),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1136),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_297),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1212),
.Y(n_1343)
);

BUFx8_ASAP7_75t_SL g1344 ( 
.A(n_111),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_390),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_106),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_569),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1285),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_295),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1016),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_219),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_995),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1138),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1071),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_798),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1134),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1255),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_751),
.Y(n_1358)
);

BUFx2_ASAP7_75t_SL g1359 ( 
.A(n_601),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_459),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1072),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_388),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1181),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_486),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_661),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1120),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_796),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_602),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_490),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_934),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_963),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_187),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_593),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_254),
.Y(n_1374)
);

CKINVDCx16_ASAP7_75t_R g1375 ( 
.A(n_1172),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_966),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1262),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1188),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_680),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1200),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1208),
.Y(n_1381)
);

INVxp67_ASAP7_75t_L g1382 ( 
.A(n_525),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_190),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1142),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1242),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_332),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_977),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_301),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1192),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_835),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_64),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_471),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_514),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_557),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_978),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1149),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1279),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_276),
.Y(n_1398)
);

CKINVDCx14_ASAP7_75t_R g1399 ( 
.A(n_559),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_924),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_839),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1275),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_26),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_446),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_205),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_946),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1055),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_721),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_404),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_337),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_547),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_463),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1197),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_998),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_419),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_475),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1258),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1007),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1177),
.Y(n_1419)
);

INVxp33_ASAP7_75t_L g1420 ( 
.A(n_895),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_657),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_56),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_933),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_807),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_753),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_218),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1203),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1057),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_979),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1083),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_570),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_277),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_988),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_191),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_879),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1270),
.Y(n_1436)
);

CKINVDCx16_ASAP7_75t_R g1437 ( 
.A(n_603),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_542),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_468),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_893),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_929),
.Y(n_1441)
);

BUFx10_ASAP7_75t_L g1442 ( 
.A(n_736),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1226),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1286),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_577),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_337),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_506),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_702),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_324),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1089),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1154),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_615),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_991),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1191),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1027),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_363),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_499),
.Y(n_1457)
);

BUFx5_ASAP7_75t_L g1458 ( 
.A(n_1107),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1207),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_401),
.Y(n_1460)
);

BUFx10_ASAP7_75t_L g1461 ( 
.A(n_184),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_539),
.Y(n_1462)
);

CKINVDCx20_ASAP7_75t_R g1463 ( 
.A(n_200),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_83),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_615),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_658),
.Y(n_1466)
);

CKINVDCx16_ASAP7_75t_R g1467 ( 
.A(n_529),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_782),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_299),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_712),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_423),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1021),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_781),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_943),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_293),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_623),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_254),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_457),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1044),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_49),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1159),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1152),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1199),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1113),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1000),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_747),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_780),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_222),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1040),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1095),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_333),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1160),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_7),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_958),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_862),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_223),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_614),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_954),
.Y(n_1498)
);

BUFx10_ASAP7_75t_L g1499 ( 
.A(n_843),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_639),
.Y(n_1500)
);

BUFx5_ASAP7_75t_L g1501 ( 
.A(n_798),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1263),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_395),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_483),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_920),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_801),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_635),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_180),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_780),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_207),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_648),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1259),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_391),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_766),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1187),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_61),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_764),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1150),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1171),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_678),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_938),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_319),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_824),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_298),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_723),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1110),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_812),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1291),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_872),
.Y(n_1529)
);

CKINVDCx20_ASAP7_75t_R g1530 ( 
.A(n_576),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_877),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_742),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1224),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1049),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1086),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1166),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_613),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_692),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_870),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_391),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_41),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_819),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_1024),
.Y(n_1543)
);

CKINVDCx16_ASAP7_75t_R g1544 ( 
.A(n_1041),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_140),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_302),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1228),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_107),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_538),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_897),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1237),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1126),
.Y(n_1552)
);

CKINVDCx16_ASAP7_75t_R g1553 ( 
.A(n_1202),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1018),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_518),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_779),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_993),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_247),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_567),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_646),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_630),
.Y(n_1561)
);

CKINVDCx16_ASAP7_75t_R g1562 ( 
.A(n_990),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_491),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1065),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_838),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_130),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1183),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_790),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_1139),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_885),
.Y(n_1570)
);

CKINVDCx16_ASAP7_75t_R g1571 ( 
.A(n_366),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_612),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_822),
.Y(n_1573)
);

BUFx5_ASAP7_75t_L g1574 ( 
.A(n_956),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1075),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1243),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1011),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_999),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_31),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_502),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_104),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1017),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_20),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_190),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_44),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_749),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_834),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_96),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1067),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_432),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_10),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_884),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_200),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_378),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_655),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1215),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1218),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_683),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_515),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_673),
.Y(n_1600)
);

CKINVDCx16_ASAP7_75t_R g1601 ( 
.A(n_1050),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1022),
.Y(n_1602)
);

CKINVDCx20_ASAP7_75t_R g1603 ( 
.A(n_542),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_1090),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_449),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_533),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_941),
.Y(n_1607)
);

BUFx10_ASAP7_75t_L g1608 ( 
.A(n_1000),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1289),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1161),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_677),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1168),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_2),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1216),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_329),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_568),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_246),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1165),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_922),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1238),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_608),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_669),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1250),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_787),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1204),
.Y(n_1625)
);

BUFx10_ASAP7_75t_L g1626 ( 
.A(n_688),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_502),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_666),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_651),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_913),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_704),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_330),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_130),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1211),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_412),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_36),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1180),
.Y(n_1637)
);

CKINVDCx20_ASAP7_75t_R g1638 ( 
.A(n_674),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_876),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_799),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_225),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_348),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_314),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_393),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_411),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_813),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_793),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1047),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_84),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_271),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1283),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1293),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_622),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_590),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_952),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_544),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_903),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1213),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_221),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_700),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1143),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1145),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1131),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1151),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_761),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_968),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1194),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_277),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1146),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1190),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1210),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_340),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1062),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_975),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_90),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1111),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_50),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_805),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_462),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_392),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_197),
.Y(n_1681)
);

BUFx10_ASAP7_75t_L g1682 ( 
.A(n_1006),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1016),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_918),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_87),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1214),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1153),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_933),
.Y(n_1688)
);

BUFx10_ASAP7_75t_L g1689 ( 
.A(n_1260),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1132),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_543),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_981),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1278),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1292),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_39),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1029),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_65),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1267),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_643),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1003),
.Y(n_1700)
);

CKINVDCx20_ASAP7_75t_R g1701 ( 
.A(n_1287),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_499),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_812),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_697),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_156),
.Y(n_1705)
);

BUFx3_ASAP7_75t_L g1706 ( 
.A(n_754),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_517),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_913),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_593),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1070),
.Y(n_1710)
);

BUFx10_ASAP7_75t_L g1711 ( 
.A(n_215),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_985),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_328),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_311),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_603),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_485),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_909),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_1249),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_244),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_957),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1222),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_247),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1014),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_1239),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_747),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1282),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_459),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1060),
.Y(n_1728)
);

INVxp33_ASAP7_75t_R g1729 ( 
.A(n_7),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_830),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_727),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_114),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_338),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1245),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_160),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_196),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_655),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_255),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_775),
.Y(n_1739)
);

CKINVDCx20_ASAP7_75t_R g1740 ( 
.A(n_554),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_577),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_678),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_74),
.Y(n_1743)
);

CKINVDCx16_ASAP7_75t_R g1744 ( 
.A(n_974),
.Y(n_1744)
);

BUFx10_ASAP7_75t_L g1745 ( 
.A(n_380),
.Y(n_1745)
);

BUFx10_ASAP7_75t_L g1746 ( 
.A(n_832),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_755),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_146),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1193),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_146),
.Y(n_1750)
);

CKINVDCx20_ASAP7_75t_R g1751 ( 
.A(n_580),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_475),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1137),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_217),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1186),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1020),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_860),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_984),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_867),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1082),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_549),
.Y(n_1761)
);

CKINVDCx20_ASAP7_75t_R g1762 ( 
.A(n_667),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_243),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_914),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1158),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_917),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1264),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_828),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_894),
.Y(n_1769)
);

CKINVDCx20_ASAP7_75t_R g1770 ( 
.A(n_1004),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_701),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_163),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_992),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1119),
.Y(n_1774)
);

CKINVDCx16_ASAP7_75t_R g1775 ( 
.A(n_989),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1042),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1125),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_859),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_60),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_184),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1219),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_706),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1196),
.Y(n_1783)
);

CKINVDCx20_ASAP7_75t_R g1784 ( 
.A(n_1028),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_127),
.Y(n_1785)
);

CKINVDCx20_ASAP7_75t_R g1786 ( 
.A(n_731),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_301),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_95),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1209),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_51),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_467),
.Y(n_1791)
);

CKINVDCx20_ASAP7_75t_R g1792 ( 
.A(n_265),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_266),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1034),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_909),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_820),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_137),
.Y(n_1797)
);

BUFx5_ASAP7_75t_L g1798 ( 
.A(n_201),
.Y(n_1798)
);

BUFx6f_ASAP7_75t_L g1799 ( 
.A(n_522),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1116),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_225),
.Y(n_1801)
);

BUFx5_ASAP7_75t_L g1802 ( 
.A(n_1217),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_164),
.Y(n_1803)
);

BUFx5_ASAP7_75t_L g1804 ( 
.A(n_583),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1227),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_626),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_848),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_714),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1122),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1109),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_246),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_952),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_10),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1244),
.Y(n_1814)
);

CKINVDCx20_ASAP7_75t_R g1815 ( 
.A(n_590),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_306),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_994),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_631),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_720),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_196),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_866),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_701),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_490),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1272),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1015),
.Y(n_1825)
);

CKINVDCx20_ASAP7_75t_R g1826 ( 
.A(n_321),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_720),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1129),
.Y(n_1828)
);

INVx1_ASAP7_75t_SL g1829 ( 
.A(n_387),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_928),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1254),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_1167),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_585),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1093),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_538),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_163),
.Y(n_1836)
);

CKINVDCx16_ASAP7_75t_R g1837 ( 
.A(n_1290),
.Y(n_1837)
);

CKINVDCx20_ASAP7_75t_R g1838 ( 
.A(n_787),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_176),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_407),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_412),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_253),
.Y(n_1842)
);

INVx1_ASAP7_75t_SL g1843 ( 
.A(n_1276),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_455),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_963),
.Y(n_1845)
);

BUFx10_ASAP7_75t_L g1846 ( 
.A(n_397),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1079),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_672),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1030),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_18),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_188),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_596),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_386),
.Y(n_1853)
);

CKINVDCx14_ASAP7_75t_R g1854 ( 
.A(n_657),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_336),
.Y(n_1855)
);

BUFx6f_ASAP7_75t_L g1856 ( 
.A(n_528),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_249),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1084),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_644),
.Y(n_1859)
);

BUFx2_ASAP7_75t_L g1860 ( 
.A(n_84),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_1038),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1229),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_861),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1174),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1284),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_976),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1002),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_956),
.Y(n_1868)
);

BUFx10_ASAP7_75t_L g1869 ( 
.A(n_30),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_889),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_92),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_809),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_696),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_837),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_800),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_1230),
.Y(n_1876)
);

BUFx6f_ASAP7_75t_L g1877 ( 
.A(n_1198),
.Y(n_1877)
);

BUFx8_ASAP7_75t_SL g1878 ( 
.A(n_878),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_432),
.Y(n_1879)
);

CKINVDCx20_ASAP7_75t_R g1880 ( 
.A(n_980),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1005),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1098),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_934),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_639),
.Y(n_1884)
);

BUFx10_ASAP7_75t_L g1885 ( 
.A(n_1162),
.Y(n_1885)
);

BUFx2_ASAP7_75t_L g1886 ( 
.A(n_1030),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_806),
.Y(n_1887)
);

CKINVDCx20_ASAP7_75t_R g1888 ( 
.A(n_1164),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_346),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_145),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1256),
.Y(n_1891)
);

INVx2_ASAP7_75t_SL g1892 ( 
.A(n_553),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1010),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_551),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_690),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_915),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1274),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_372),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_49),
.Y(n_1899)
);

CKINVDCx16_ASAP7_75t_R g1900 ( 
.A(n_245),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_318),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_907),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1114),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_693),
.Y(n_1904)
);

CKINVDCx16_ASAP7_75t_R g1905 ( 
.A(n_1248),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1179),
.Y(n_1906)
);

BUFx3_ASAP7_75t_L g1907 ( 
.A(n_37),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_345),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1280),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_842),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_758),
.Y(n_1911)
);

INVxp67_ASAP7_75t_L g1912 ( 
.A(n_1176),
.Y(n_1912)
);

INVx1_ASAP7_75t_SL g1913 ( 
.A(n_471),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_338),
.Y(n_1914)
);

INVx1_ASAP7_75t_SL g1915 ( 
.A(n_1169),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_559),
.Y(n_1916)
);

BUFx2_ASAP7_75t_L g1917 ( 
.A(n_555),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_722),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1268),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_1257),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_883),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1013),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_527),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_946),
.Y(n_1924)
);

CKINVDCx20_ASAP7_75t_R g1925 ( 
.A(n_183),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_667),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_759),
.Y(n_1927)
);

INVx1_ASAP7_75t_SL g1928 ( 
.A(n_755),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_664),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_526),
.Y(n_1930)
);

CKINVDCx20_ASAP7_75t_R g1931 ( 
.A(n_4),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_1025),
.Y(n_1932)
);

BUFx10_ASAP7_75t_L g1933 ( 
.A(n_487),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_644),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1144),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_982),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1265),
.Y(n_1937)
);

CKINVDCx20_ASAP7_75t_R g1938 ( 
.A(n_1043),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1261),
.Y(n_1939)
);

INVx2_ASAP7_75t_SL g1940 ( 
.A(n_1233),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1157),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1221),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_275),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_669),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_519),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1039),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1147),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_631),
.Y(n_1948)
);

INVx2_ASAP7_75t_SL g1949 ( 
.A(n_279),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1271),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_996),
.Y(n_1951)
);

CKINVDCx16_ASAP7_75t_R g1952 ( 
.A(n_1269),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_570),
.Y(n_1953)
);

BUFx3_ASAP7_75t_L g1954 ( 
.A(n_1102),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1247),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_861),
.Y(n_1956)
);

BUFx3_ASAP7_75t_L g1957 ( 
.A(n_1246),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1045),
.Y(n_1958)
);

CKINVDCx20_ASAP7_75t_R g1959 ( 
.A(n_323),
.Y(n_1959)
);

BUFx8_ASAP7_75t_SL g1960 ( 
.A(n_870),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_878),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_357),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_61),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_2),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_733),
.Y(n_1965)
);

BUFx3_ASAP7_75t_L g1966 ( 
.A(n_623),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_726),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_365),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_282),
.Y(n_1969)
);

BUFx3_ASAP7_75t_L g1970 ( 
.A(n_726),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1032),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_735),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_192),
.Y(n_1973)
);

CKINVDCx20_ASAP7_75t_R g1974 ( 
.A(n_1178),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_182),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_573),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_897),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_786),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_728),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1163),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_356),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_765),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_380),
.Y(n_1983)
);

CKINVDCx16_ASAP7_75t_R g1984 ( 
.A(n_723),
.Y(n_1984)
);

CKINVDCx20_ASAP7_75t_R g1985 ( 
.A(n_1019),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1273),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_598),
.Y(n_1987)
);

BUFx10_ASAP7_75t_L g1988 ( 
.A(n_44),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_284),
.Y(n_1989)
);

BUFx3_ASAP7_75t_L g1990 ( 
.A(n_318),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_766),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_857),
.Y(n_1992)
);

BUFx6f_ASAP7_75t_L g1993 ( 
.A(n_1184),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_74),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1156),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1173),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_267),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1009),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_1185),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_983),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1266),
.Y(n_2001)
);

BUFx5_ASAP7_75t_L g2002 ( 
.A(n_856),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_582),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_527),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1105),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_469),
.Y(n_2006)
);

INVx1_ASAP7_75t_SL g2007 ( 
.A(n_369),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_126),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1223),
.Y(n_2009)
);

CKINVDCx20_ASAP7_75t_R g2010 ( 
.A(n_456),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_1225),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_511),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_27),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1231),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_352),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_310),
.Y(n_2016)
);

BUFx3_ASAP7_75t_L g2017 ( 
.A(n_107),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1206),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_842),
.Y(n_2019)
);

INVx1_ASAP7_75t_SL g2020 ( 
.A(n_999),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_637),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_463),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_226),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_97),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_530),
.Y(n_2025)
);

BUFx6f_ASAP7_75t_L g2026 ( 
.A(n_966),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_930),
.Y(n_2027)
);

BUFx3_ASAP7_75t_L g2028 ( 
.A(n_1018),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1205),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1241),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_304),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_968),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_576),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_997),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_544),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_1140),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_403),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1170),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_256),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_139),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_441),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1252),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1236),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_62),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_520),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_953),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_918),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1240),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1201),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_548),
.Y(n_2050)
);

CKINVDCx20_ASAP7_75t_R g2051 ( 
.A(n_430),
.Y(n_2051)
);

INVx2_ASAP7_75t_SL g2052 ( 
.A(n_959),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1033),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1031),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1061),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_892),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_47),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_951),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_874),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_1288),
.Y(n_2060)
);

CKINVDCx16_ASAP7_75t_R g2061 ( 
.A(n_987),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1001),
.Y(n_2062)
);

CKINVDCx20_ASAP7_75t_R g2063 ( 
.A(n_97),
.Y(n_2063)
);

CKINVDCx14_ASAP7_75t_R g2064 ( 
.A(n_242),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1077),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_732),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_222),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1253),
.Y(n_2068)
);

BUFx10_ASAP7_75t_L g2069 ( 
.A(n_1037),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_630),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_807),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_75),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1100),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1135),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1035),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_1012),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_287),
.Y(n_2077)
);

CKINVDCx20_ASAP7_75t_R g2078 ( 
.A(n_1235),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_1017),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_169),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_201),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_1195),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_388),
.Y(n_2083)
);

CKINVDCx20_ASAP7_75t_R g2084 ( 
.A(n_40),
.Y(n_2084)
);

INVx2_ASAP7_75t_SL g2085 ( 
.A(n_343),
.Y(n_2085)
);

CKINVDCx5p33_ASAP7_75t_R g2086 ( 
.A(n_448),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_400),
.Y(n_2087)
);

BUFx10_ASAP7_75t_L g2088 ( 
.A(n_6),
.Y(n_2088)
);

BUFx3_ASAP7_75t_L g2089 ( 
.A(n_986),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_1220),
.Y(n_2090)
);

CKINVDCx5p33_ASAP7_75t_R g2091 ( 
.A(n_485),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_803),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_784),
.Y(n_2093)
);

CKINVDCx5p33_ASAP7_75t_R g2094 ( 
.A(n_947),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1501),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1501),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1501),
.Y(n_2097)
);

INVxp67_ASAP7_75t_SL g2098 ( 
.A(n_1497),
.Y(n_2098)
);

HB1xp67_ASAP7_75t_L g2099 ( 
.A(n_1566),
.Y(n_2099)
);

INVxp67_ASAP7_75t_SL g2100 ( 
.A(n_1497),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1501),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1501),
.Y(n_2102)
);

INVxp67_ASAP7_75t_L g2103 ( 
.A(n_1368),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1574),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1574),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1574),
.Y(n_2106)
);

BUFx3_ASAP7_75t_L g2107 ( 
.A(n_1689),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1574),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1574),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1798),
.Y(n_2110)
);

INVxp33_ASAP7_75t_L g2111 ( 
.A(n_2044),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1798),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1798),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1798),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1798),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1804),
.Y(n_2116)
);

CKINVDCx16_ASAP7_75t_R g2117 ( 
.A(n_1399),
.Y(n_2117)
);

INVxp67_ASAP7_75t_SL g2118 ( 
.A(n_1497),
.Y(n_2118)
);

INVxp33_ASAP7_75t_L g2119 ( 
.A(n_1344),
.Y(n_2119)
);

CKINVDCx16_ASAP7_75t_R g2120 ( 
.A(n_1854),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1804),
.Y(n_2121)
);

INVxp67_ASAP7_75t_SL g2122 ( 
.A(n_1506),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1804),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1804),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1804),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2002),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2002),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2002),
.Y(n_2128)
);

BUFx3_ASAP7_75t_L g2129 ( 
.A(n_1689),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2002),
.Y(n_2130)
);

INVxp33_ASAP7_75t_SL g2131 ( 
.A(n_1616),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2002),
.Y(n_2132)
);

CKINVDCx16_ASAP7_75t_R g2133 ( 
.A(n_2064),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1302),
.Y(n_2134)
);

CKINVDCx14_ASAP7_75t_R g2135 ( 
.A(n_1885),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1310),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1320),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1327),
.Y(n_2138)
);

BUFx10_ASAP7_75t_L g2139 ( 
.A(n_1668),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1329),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1330),
.Y(n_2141)
);

INVxp67_ASAP7_75t_SL g2142 ( 
.A(n_1506),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1332),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1333),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1336),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1337),
.Y(n_2146)
);

INVxp67_ASAP7_75t_SL g2147 ( 
.A(n_1506),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1340),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1350),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_1878),
.Y(n_2150)
);

NOR2xp33_ASAP7_75t_L g2151 ( 
.A(n_1420),
.B(n_1),
.Y(n_2151)
);

INVxp67_ASAP7_75t_L g2152 ( 
.A(n_1720),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1360),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1364),
.Y(n_2154)
);

CKINVDCx14_ASAP7_75t_R g2155 ( 
.A(n_1885),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1371),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_1960),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1372),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1374),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1376),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1379),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1388),
.Y(n_2162)
);

BUFx6f_ASAP7_75t_L g2163 ( 
.A(n_1590),
.Y(n_2163)
);

BUFx6f_ASAP7_75t_L g2164 ( 
.A(n_1590),
.Y(n_2164)
);

CKINVDCx16_ASAP7_75t_R g2165 ( 
.A(n_1437),
.Y(n_2165)
);

INVxp33_ASAP7_75t_SL g2166 ( 
.A(n_1860),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1393),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1395),
.Y(n_2168)
);

BUFx3_ASAP7_75t_L g2169 ( 
.A(n_1492),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1400),
.Y(n_2170)
);

BUFx5_ASAP7_75t_L g2171 ( 
.A(n_1298),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1411),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1412),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1426),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1435),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1590),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1592),
.Y(n_2177)
);

CKINVDCx20_ASAP7_75t_R g2178 ( 
.A(n_1341),
.Y(n_2178)
);

INVxp33_ASAP7_75t_SL g2179 ( 
.A(n_1886),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1438),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1445),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1448),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1453),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_1467),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1465),
.Y(n_2185)
);

CKINVDCx16_ASAP7_75t_R g2186 ( 
.A(n_1544),
.Y(n_2186)
);

BUFx2_ASAP7_75t_SL g2187 ( 
.A(n_1484),
.Y(n_2187)
);

INVxp67_ASAP7_75t_L g2188 ( 
.A(n_1917),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1592),
.Y(n_2189)
);

CKINVDCx20_ASAP7_75t_R g2190 ( 
.A(n_1569),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1468),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_1562),
.Y(n_2192)
);

CKINVDCx20_ASAP7_75t_R g2193 ( 
.A(n_1604),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1472),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1475),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1477),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1478),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1592),
.Y(n_2198)
);

CKINVDCx5p33_ASAP7_75t_R g2199 ( 
.A(n_1571),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1487),
.Y(n_2200)
);

INVxp33_ASAP7_75t_SL g2201 ( 
.A(n_1359),
.Y(n_2201)
);

CKINVDCx14_ASAP7_75t_R g2202 ( 
.A(n_1701),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1639),
.Y(n_2203)
);

INVxp33_ASAP7_75t_L g2204 ( 
.A(n_1308),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1489),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_1639),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1494),
.Y(n_2207)
);

INVxp67_ASAP7_75t_SL g2208 ( 
.A(n_1639),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1504),
.Y(n_2209)
);

BUFx6f_ASAP7_75t_L g2210 ( 
.A(n_1695),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1507),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1508),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1695),
.Y(n_2213)
);

CKINVDCx16_ASAP7_75t_R g2214 ( 
.A(n_1744),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1513),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1517),
.Y(n_2216)
);

INVxp33_ASAP7_75t_SL g2217 ( 
.A(n_1296),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_1775),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1524),
.Y(n_2219)
);

INVxp33_ASAP7_75t_SL g2220 ( 
.A(n_1300),
.Y(n_2220)
);

INVxp33_ASAP7_75t_SL g2221 ( 
.A(n_1304),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1532),
.Y(n_2222)
);

INVxp67_ASAP7_75t_SL g2223 ( 
.A(n_1695),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1554),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1555),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1799),
.Y(n_2226)
);

INVxp33_ASAP7_75t_SL g2227 ( 
.A(n_1306),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1559),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1561),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1573),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1799),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1799),
.Y(n_2232)
);

INVxp33_ASAP7_75t_SL g2233 ( 
.A(n_1309),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1856),
.Y(n_2234)
);

INVxp67_ASAP7_75t_L g2235 ( 
.A(n_1326),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1584),
.Y(n_2236)
);

INVxp33_ASAP7_75t_SL g2237 ( 
.A(n_1311),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1591),
.Y(n_2238)
);

INVxp67_ASAP7_75t_SL g2239 ( 
.A(n_1856),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1593),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1595),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_1856),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1602),
.Y(n_2243)
);

INVx2_ASAP7_75t_SL g2244 ( 
.A(n_1442),
.Y(n_2244)
);

INVxp33_ASAP7_75t_L g2245 ( 
.A(n_1346),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1621),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1627),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1629),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_1900),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1631),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1632),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1635),
.Y(n_2252)
);

INVxp33_ASAP7_75t_SL g2253 ( 
.A(n_1312),
.Y(n_2253)
);

CKINVDCx14_ASAP7_75t_R g2254 ( 
.A(n_1721),
.Y(n_2254)
);

CKINVDCx16_ASAP7_75t_R g2255 ( 
.A(n_1984),
.Y(n_2255)
);

BUFx6f_ASAP7_75t_L g2256 ( 
.A(n_1976),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1636),
.Y(n_2257)
);

CKINVDCx16_ASAP7_75t_R g2258 ( 
.A(n_2061),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1640),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2098),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2163),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2100),
.Y(n_2262)
);

CKINVDCx20_ASAP7_75t_R g2263 ( 
.A(n_2178),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2118),
.Y(n_2264)
);

BUFx6f_ASAP7_75t_L g2265 ( 
.A(n_2163),
.Y(n_2265)
);

INVx5_ASAP7_75t_L g2266 ( 
.A(n_2165),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_2107),
.B(n_1375),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2122),
.Y(n_2268)
);

INVx3_ASAP7_75t_L g2269 ( 
.A(n_2169),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_2164),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_2184),
.Y(n_2271)
);

OA21x2_ASAP7_75t_L g2272 ( 
.A1(n_2095),
.A2(n_1348),
.B(n_1324),
.Y(n_2272)
);

OA21x2_ASAP7_75t_L g2273 ( 
.A1(n_2096),
.A2(n_2101),
.B(n_2097),
.Y(n_2273)
);

OA21x2_ASAP7_75t_L g2274 ( 
.A1(n_2102),
.A2(n_1363),
.B(n_1356),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2142),
.Y(n_2275)
);

BUFx6f_ASAP7_75t_L g2276 ( 
.A(n_2164),
.Y(n_2276)
);

AND2x4_ASAP7_75t_L g2277 ( 
.A(n_2129),
.B(n_1334),
.Y(n_2277)
);

CKINVDCx5p33_ASAP7_75t_R g2278 ( 
.A(n_2202),
.Y(n_2278)
);

OAI22x1_ASAP7_75t_R g2279 ( 
.A1(n_2150),
.A2(n_1342),
.B1(n_1365),
.B2(n_1328),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2147),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2208),
.Y(n_2281)
);

OAI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_2103),
.A2(n_2152),
.B1(n_2188),
.B2(n_2166),
.Y(n_2282)
);

BUFx6f_ASAP7_75t_L g2283 ( 
.A(n_2206),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2223),
.B(n_1553),
.Y(n_2284)
);

BUFx6f_ASAP7_75t_L g2285 ( 
.A(n_2206),
.Y(n_2285)
);

OAI22xp5_ASAP7_75t_SL g2286 ( 
.A1(n_2190),
.A2(n_1440),
.B1(n_1463),
.B2(n_1432),
.Y(n_2286)
);

BUFx12f_ASAP7_75t_L g2287 ( 
.A(n_2157),
.Y(n_2287)
);

CKINVDCx16_ASAP7_75t_R g2288 ( 
.A(n_2117),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2239),
.Y(n_2289)
);

BUFx8_ASAP7_75t_L g2290 ( 
.A(n_2244),
.Y(n_2290)
);

INVx2_ASAP7_75t_SL g2291 ( 
.A(n_2139),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2210),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2104),
.Y(n_2293)
);

CKINVDCx5p33_ASAP7_75t_R g2294 ( 
.A(n_2254),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2171),
.B(n_1601),
.Y(n_2295)
);

OA21x2_ASAP7_75t_L g2296 ( 
.A1(n_2105),
.A2(n_1417),
.B(n_1385),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2171),
.B(n_1837),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2106),
.Y(n_2298)
);

BUFx6f_ASAP7_75t_L g2299 ( 
.A(n_2210),
.Y(n_2299)
);

INVx5_ASAP7_75t_L g2300 ( 
.A(n_2186),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2108),
.Y(n_2301)
);

BUFx6f_ASAP7_75t_L g2302 ( 
.A(n_2226),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2226),
.Y(n_2303)
);

OAI21x1_ASAP7_75t_L g2304 ( 
.A1(n_2114),
.A2(n_2110),
.B(n_2109),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_2187),
.Y(n_2305)
);

INVx2_ASAP7_75t_SL g2306 ( 
.A(n_2192),
.Y(n_2306)
);

BUFx8_ASAP7_75t_SL g2307 ( 
.A(n_2193),
.Y(n_2307)
);

BUFx6f_ASAP7_75t_L g2308 ( 
.A(n_2242),
.Y(n_2308)
);

INVx5_ASAP7_75t_L g2309 ( 
.A(n_2242),
.Y(n_2309)
);

OAI22x1_ASAP7_75t_L g2310 ( 
.A1(n_2099),
.A2(n_1729),
.B1(n_2218),
.B2(n_2199),
.Y(n_2310)
);

INVx4_ASAP7_75t_L g2311 ( 
.A(n_2120),
.Y(n_2311)
);

CKINVDCx5p33_ASAP7_75t_R g2312 ( 
.A(n_2135),
.Y(n_2312)
);

INVx3_ASAP7_75t_L g2313 ( 
.A(n_2256),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2256),
.Y(n_2314)
);

INVx3_ASAP7_75t_L g2315 ( 
.A(n_2176),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2177),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2189),
.Y(n_2317)
);

BUFx3_ASAP7_75t_L g2318 ( 
.A(n_2112),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2198),
.Y(n_2319)
);

INVx3_ASAP7_75t_L g2320 ( 
.A(n_2203),
.Y(n_2320)
);

BUFx8_ASAP7_75t_SL g2321 ( 
.A(n_2249),
.Y(n_2321)
);

BUFx6f_ASAP7_75t_L g2322 ( 
.A(n_2213),
.Y(n_2322)
);

BUFx8_ASAP7_75t_SL g2323 ( 
.A(n_2134),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2171),
.B(n_1905),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2155),
.B(n_1952),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2231),
.Y(n_2326)
);

CKINVDCx20_ASAP7_75t_R g2327 ( 
.A(n_2133),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_L g2328 ( 
.A(n_2217),
.B(n_2220),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2113),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2115),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_L g2331 ( 
.A(n_2221),
.B(n_1912),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_2232),
.Y(n_2332)
);

INVx4_ASAP7_75t_L g2333 ( 
.A(n_2171),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2116),
.Y(n_2334)
);

AND2x4_ASAP7_75t_L g2335 ( 
.A(n_2235),
.B(n_1392),
.Y(n_2335)
);

CKINVDCx5p33_ASAP7_75t_R g2336 ( 
.A(n_2227),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_2234),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2121),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_2233),
.B(n_1430),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2123),
.Y(n_2340)
);

BUFx6f_ASAP7_75t_L g2341 ( 
.A(n_2136),
.Y(n_2341)
);

INVx3_ASAP7_75t_L g2342 ( 
.A(n_2137),
.Y(n_2342)
);

BUFx6f_ASAP7_75t_L g2343 ( 
.A(n_2138),
.Y(n_2343)
);

INVx5_ASAP7_75t_L g2344 ( 
.A(n_2214),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2124),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2204),
.B(n_1442),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2125),
.Y(n_2347)
);

BUFx12f_ASAP7_75t_L g2348 ( 
.A(n_2119),
.Y(n_2348)
);

AND2x6_ASAP7_75t_L g2349 ( 
.A(n_2140),
.B(n_2141),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2126),
.Y(n_2350)
);

BUFx6f_ASAP7_75t_L g2351 ( 
.A(n_2143),
.Y(n_2351)
);

INVx5_ASAP7_75t_L g2352 ( 
.A(n_2255),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2127),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2128),
.Y(n_2354)
);

INVx2_ASAP7_75t_SL g2355 ( 
.A(n_2258),
.Y(n_2355)
);

INVx3_ASAP7_75t_L g2356 ( 
.A(n_2144),
.Y(n_2356)
);

BUFx6f_ASAP7_75t_L g2357 ( 
.A(n_2145),
.Y(n_2357)
);

INVx3_ASAP7_75t_L g2358 ( 
.A(n_2146),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_2148),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_2149),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_L g2361 ( 
.A(n_2237),
.B(n_2253),
.Y(n_2361)
);

BUFx8_ASAP7_75t_SL g2362 ( 
.A(n_2259),
.Y(n_2362)
);

AND2x4_ASAP7_75t_L g2363 ( 
.A(n_2153),
.B(n_1462),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2130),
.Y(n_2364)
);

INVx5_ASAP7_75t_L g2365 ( 
.A(n_2201),
.Y(n_2365)
);

BUFx3_ASAP7_75t_L g2366 ( 
.A(n_2132),
.Y(n_2366)
);

BUFx8_ASAP7_75t_SL g2367 ( 
.A(n_2154),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_2156),
.Y(n_2368)
);

AOI22xp5_ASAP7_75t_L g2369 ( 
.A1(n_2131),
.A2(n_1543),
.B1(n_1556),
.B2(n_1530),
.Y(n_2369)
);

INVx5_ASAP7_75t_L g2370 ( 
.A(n_2179),
.Y(n_2370)
);

HB1xp67_ASAP7_75t_L g2371 ( 
.A(n_2111),
.Y(n_2371)
);

BUFx6f_ASAP7_75t_L g2372 ( 
.A(n_2158),
.Y(n_2372)
);

OA21x2_ASAP7_75t_L g2373 ( 
.A1(n_2159),
.A2(n_1444),
.B(n_1443),
.Y(n_2373)
);

OAI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2151),
.A2(n_1638),
.B1(n_1643),
.B2(n_1603),
.Y(n_2374)
);

INVx6_ASAP7_75t_L g2375 ( 
.A(n_2245),
.Y(n_2375)
);

INVx5_ASAP7_75t_L g2376 ( 
.A(n_2160),
.Y(n_2376)
);

HB1xp67_ASAP7_75t_L g2377 ( 
.A(n_2161),
.Y(n_2377)
);

BUFx6f_ASAP7_75t_L g2378 ( 
.A(n_2162),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2167),
.Y(n_2379)
);

INVx3_ASAP7_75t_L g2380 ( 
.A(n_2168),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_2170),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_2172),
.B(n_1471),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2173),
.B(n_1461),
.Y(n_2383)
);

AOI22x1_ASAP7_75t_SL g2384 ( 
.A1(n_2174),
.A2(n_1719),
.B1(n_1731),
.B2(n_1656),
.Y(n_2384)
);

BUFx12f_ASAP7_75t_L g2385 ( 
.A(n_2175),
.Y(n_2385)
);

AND2x4_ASAP7_75t_L g2386 ( 
.A(n_2180),
.B(n_1480),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2181),
.Y(n_2387)
);

BUFx6f_ASAP7_75t_L g2388 ( 
.A(n_2182),
.Y(n_2388)
);

BUFx6f_ASAP7_75t_L g2389 ( 
.A(n_2183),
.Y(n_2389)
);

OAI22xp5_ASAP7_75t_L g2390 ( 
.A1(n_2185),
.A2(n_1751),
.B1(n_1762),
.B2(n_1740),
.Y(n_2390)
);

BUFx6f_ASAP7_75t_L g2391 ( 
.A(n_2191),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_2194),
.B(n_2195),
.Y(n_2392)
);

BUFx3_ASAP7_75t_L g2393 ( 
.A(n_2196),
.Y(n_2393)
);

OAI22x1_ASAP7_75t_SL g2394 ( 
.A1(n_2197),
.A2(n_1771),
.B1(n_1784),
.B2(n_1770),
.Y(n_2394)
);

AOI22x1_ASAP7_75t_SL g2395 ( 
.A1(n_2200),
.A2(n_1792),
.B1(n_1815),
.B2(n_1786),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2205),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2207),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2209),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2211),
.B(n_1461),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2212),
.Y(n_2400)
);

OAI21x1_ASAP7_75t_L g2401 ( 
.A1(n_2257),
.A2(n_1481),
.B(n_1451),
.Y(n_2401)
);

AND2x6_ASAP7_75t_L g2402 ( 
.A(n_2215),
.B(n_1516),
.Y(n_2402)
);

INVx5_ASAP7_75t_L g2403 ( 
.A(n_2216),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2219),
.Y(n_2404)
);

BUFx6f_ASAP7_75t_L g2405 ( 
.A(n_2222),
.Y(n_2405)
);

BUFx6f_ASAP7_75t_L g2406 ( 
.A(n_2224),
.Y(n_2406)
);

CKINVDCx20_ASAP7_75t_R g2407 ( 
.A(n_2225),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2228),
.Y(n_2408)
);

BUFx6f_ASAP7_75t_L g2409 ( 
.A(n_2229),
.Y(n_2409)
);

BUFx6f_ASAP7_75t_L g2410 ( 
.A(n_2230),
.Y(n_2410)
);

BUFx6f_ASAP7_75t_L g2411 ( 
.A(n_2236),
.Y(n_2411)
);

INVx4_ASAP7_75t_L g2412 ( 
.A(n_2238),
.Y(n_2412)
);

AOI22xp5_ASAP7_75t_L g2413 ( 
.A1(n_2240),
.A2(n_1838),
.B1(n_1880),
.B2(n_1826),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2241),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_2252),
.B(n_1502),
.Y(n_2415)
);

BUFx3_ASAP7_75t_L g2416 ( 
.A(n_2243),
.Y(n_2416)
);

BUFx12f_ASAP7_75t_L g2417 ( 
.A(n_2246),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2247),
.Y(n_2418)
);

BUFx3_ASAP7_75t_L g2419 ( 
.A(n_2248),
.Y(n_2419)
);

BUFx2_ASAP7_75t_L g2420 ( 
.A(n_2250),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2251),
.Y(n_2421)
);

BUFx8_ASAP7_75t_SL g2422 ( 
.A(n_2178),
.Y(n_2422)
);

BUFx6f_ASAP7_75t_L g2423 ( 
.A(n_2163),
.Y(n_2423)
);

AND2x6_ASAP7_75t_L g2424 ( 
.A(n_2107),
.B(n_1568),
.Y(n_2424)
);

AND2x4_ASAP7_75t_L g2425 ( 
.A(n_2107),
.B(n_1577),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2098),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2098),
.Y(n_2427)
);

INVx3_ASAP7_75t_L g2428 ( 
.A(n_2169),
.Y(n_2428)
);

BUFx12f_ASAP7_75t_L g2429 ( 
.A(n_2150),
.Y(n_2429)
);

INVxp67_ASAP7_75t_SL g2430 ( 
.A(n_2235),
.Y(n_2430)
);

BUFx6f_ASAP7_75t_L g2431 ( 
.A(n_2163),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2163),
.Y(n_2432)
);

NOR2x1_ASAP7_75t_L g2433 ( 
.A(n_2107),
.B(n_1954),
.Y(n_2433)
);

OA21x2_ASAP7_75t_L g2434 ( 
.A1(n_2095),
.A2(n_1528),
.B(n_1512),
.Y(n_2434)
);

INVx2_ASAP7_75t_SL g2435 ( 
.A(n_2107),
.Y(n_2435)
);

INVxp67_ASAP7_75t_L g2436 ( 
.A(n_2107),
.Y(n_2436)
);

BUFx6f_ASAP7_75t_L g2437 ( 
.A(n_2163),
.Y(n_2437)
);

INVxp33_ASAP7_75t_SL g2438 ( 
.A(n_2187),
.Y(n_2438)
);

BUFx8_ASAP7_75t_SL g2439 ( 
.A(n_2178),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2135),
.B(n_1499),
.Y(n_2440)
);

BUFx3_ASAP7_75t_L g2441 ( 
.A(n_2169),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2169),
.B(n_1533),
.Y(n_2442)
);

INVx3_ASAP7_75t_L g2443 ( 
.A(n_2169),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2169),
.B(n_1535),
.Y(n_2444)
);

BUFx6f_ASAP7_75t_L g2445 ( 
.A(n_2163),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2163),
.Y(n_2446)
);

INVx5_ASAP7_75t_L g2447 ( 
.A(n_2165),
.Y(n_2447)
);

AND2x4_ASAP7_75t_L g2448 ( 
.A(n_2107),
.B(n_1606),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2163),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2098),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2163),
.Y(n_2451)
);

BUFx6f_ASAP7_75t_L g2452 ( 
.A(n_2163),
.Y(n_2452)
);

BUFx6f_ASAP7_75t_L g2453 ( 
.A(n_2163),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2163),
.Y(n_2454)
);

CKINVDCx5p33_ASAP7_75t_R g2455 ( 
.A(n_2202),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2169),
.B(n_1551),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2169),
.B(n_1564),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2169),
.B(n_1567),
.Y(n_2458)
);

BUFx2_ASAP7_75t_L g2459 ( 
.A(n_2184),
.Y(n_2459)
);

BUFx2_ASAP7_75t_L g2460 ( 
.A(n_2184),
.Y(n_2460)
);

BUFx6f_ASAP7_75t_L g2461 ( 
.A(n_2163),
.Y(n_2461)
);

AND2x2_ASAP7_75t_L g2462 ( 
.A(n_2135),
.B(n_1499),
.Y(n_2462)
);

CKINVDCx5p33_ASAP7_75t_R g2463 ( 
.A(n_2202),
.Y(n_2463)
);

INVx5_ASAP7_75t_L g2464 ( 
.A(n_2165),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2163),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2169),
.B(n_1597),
.Y(n_2466)
);

INVx2_ASAP7_75t_SL g2467 ( 
.A(n_2107),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2135),
.B(n_1608),
.Y(n_2468)
);

HB1xp67_ASAP7_75t_L g2469 ( 
.A(n_2184),
.Y(n_2469)
);

INVx2_ASAP7_75t_SL g2470 ( 
.A(n_2107),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_2107),
.B(n_1622),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_SL g2472 ( 
.A(n_2117),
.B(n_1940),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2163),
.Y(n_2473)
);

INVx3_ASAP7_75t_L g2474 ( 
.A(n_2169),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2098),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2098),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2098),
.Y(n_2477)
);

BUFx3_ASAP7_75t_L g2478 ( 
.A(n_2169),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2169),
.B(n_1634),
.Y(n_2479)
);

HB1xp67_ASAP7_75t_L g2480 ( 
.A(n_2184),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_L g2481 ( 
.A(n_2107),
.B(n_1669),
.Y(n_2481)
);

AND2x4_ASAP7_75t_L g2482 ( 
.A(n_2107),
.B(n_1706),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2163),
.Y(n_2483)
);

OAI22x1_ASAP7_75t_R g2484 ( 
.A1(n_2150),
.A2(n_1931),
.B1(n_1938),
.B2(n_1925),
.Y(n_2484)
);

BUFx6f_ASAP7_75t_L g2485 ( 
.A(n_2163),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2098),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2135),
.B(n_1608),
.Y(n_2487)
);

AND2x4_ASAP7_75t_L g2488 ( 
.A(n_2107),
.B(n_1758),
.Y(n_2488)
);

BUFx6f_ASAP7_75t_L g2489 ( 
.A(n_2163),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2098),
.Y(n_2490)
);

BUFx6f_ASAP7_75t_L g2491 ( 
.A(n_2163),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2098),
.Y(n_2492)
);

BUFx3_ASAP7_75t_L g2493 ( 
.A(n_2169),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2098),
.Y(n_2494)
);

OAI21x1_ASAP7_75t_L g2495 ( 
.A1(n_2114),
.A2(n_1694),
.B(n_1670),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2163),
.Y(n_2496)
);

HB1xp67_ASAP7_75t_L g2497 ( 
.A(n_2184),
.Y(n_2497)
);

BUFx8_ASAP7_75t_L g2498 ( 
.A(n_2107),
.Y(n_2498)
);

BUFx12f_ASAP7_75t_L g2499 ( 
.A(n_2150),
.Y(n_2499)
);

BUFx6f_ASAP7_75t_L g2500 ( 
.A(n_2163),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_2163),
.Y(n_2501)
);

BUFx8_ASAP7_75t_L g2502 ( 
.A(n_2107),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_2202),
.Y(n_2503)
);

BUFx6f_ASAP7_75t_L g2504 ( 
.A(n_2163),
.Y(n_2504)
);

OAI22xp5_ASAP7_75t_L g2505 ( 
.A1(n_2103),
.A2(n_1985),
.B1(n_2010),
.B2(n_1959),
.Y(n_2505)
);

BUFx8_ASAP7_75t_SL g2506 ( 
.A(n_2178),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2169),
.Y(n_2507)
);

BUFx6f_ASAP7_75t_L g2508 ( 
.A(n_2163),
.Y(n_2508)
);

BUFx3_ASAP7_75t_L g2509 ( 
.A(n_2169),
.Y(n_2509)
);

INVx3_ASAP7_75t_L g2510 ( 
.A(n_2169),
.Y(n_2510)
);

NOR2xp33_ASAP7_75t_L g2511 ( 
.A(n_2107),
.B(n_1765),
.Y(n_2511)
);

INVx3_ASAP7_75t_L g2512 ( 
.A(n_2169),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2163),
.Y(n_2513)
);

BUFx12f_ASAP7_75t_L g2514 ( 
.A(n_2150),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2107),
.B(n_1781),
.Y(n_2515)
);

AOI22x1_ASAP7_75t_SL g2516 ( 
.A1(n_2178),
.A2(n_2063),
.B1(n_2084),
.B2(n_2051),
.Y(n_2516)
);

BUFx3_ASAP7_75t_L g2517 ( 
.A(n_2169),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2169),
.B(n_1783),
.Y(n_2518)
);

BUFx6f_ASAP7_75t_L g2519 ( 
.A(n_2163),
.Y(n_2519)
);

BUFx2_ASAP7_75t_L g2520 ( 
.A(n_2184),
.Y(n_2520)
);

BUFx6f_ASAP7_75t_L g2521 ( 
.A(n_2163),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2163),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2169),
.B(n_1789),
.Y(n_2523)
);

INVx3_ASAP7_75t_L g2524 ( 
.A(n_2169),
.Y(n_2524)
);

HB1xp67_ASAP7_75t_L g2525 ( 
.A(n_2184),
.Y(n_2525)
);

OAI21x1_ASAP7_75t_L g2526 ( 
.A1(n_2114),
.A2(n_1864),
.B(n_1831),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2169),
.B(n_1865),
.Y(n_2527)
);

BUFx6f_ASAP7_75t_L g2528 ( 
.A(n_2163),
.Y(n_2528)
);

INVx3_ASAP7_75t_L g2529 ( 
.A(n_2169),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2135),
.B(n_1626),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2163),
.Y(n_2531)
);

BUFx6f_ASAP7_75t_L g2532 ( 
.A(n_2163),
.Y(n_2532)
);

INVx5_ASAP7_75t_L g2533 ( 
.A(n_2165),
.Y(n_2533)
);

INVx5_ASAP7_75t_L g2534 ( 
.A(n_2165),
.Y(n_2534)
);

CKINVDCx5p33_ASAP7_75t_R g2535 ( 
.A(n_2202),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2098),
.Y(n_2536)
);

AND2x4_ASAP7_75t_L g2537 ( 
.A(n_2107),
.B(n_1791),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_L g2538 ( 
.A(n_2163),
.Y(n_2538)
);

INVx2_ASAP7_75t_SL g2539 ( 
.A(n_2107),
.Y(n_2539)
);

INVx3_ASAP7_75t_L g2540 ( 
.A(n_2169),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2098),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_SL g2542 ( 
.A(n_2117),
.B(n_1888),
.Y(n_2542)
);

BUFx2_ASAP7_75t_L g2543 ( 
.A(n_2184),
.Y(n_2543)
);

BUFx2_ASAP7_75t_L g2544 ( 
.A(n_2184),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2098),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2135),
.B(n_1626),
.Y(n_2546)
);

INVx5_ASAP7_75t_L g2547 ( 
.A(n_2165),
.Y(n_2547)
);

HB1xp67_ASAP7_75t_L g2548 ( 
.A(n_2184),
.Y(n_2548)
);

BUFx2_ASAP7_75t_L g2549 ( 
.A(n_2184),
.Y(n_2549)
);

AOI22xp5_ASAP7_75t_L g2550 ( 
.A1(n_2131),
.A2(n_2078),
.B1(n_1974),
.B2(n_1315),
.Y(n_2550)
);

BUFx12f_ASAP7_75t_L g2551 ( 
.A(n_2150),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2135),
.B(n_1682),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2098),
.Y(n_2553)
);

AND2x4_ASAP7_75t_L g2554 ( 
.A(n_2107),
.B(n_1825),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2184),
.Y(n_2555)
);

BUFx3_ASAP7_75t_L g2556 ( 
.A(n_2169),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2098),
.Y(n_2557)
);

OA21x2_ASAP7_75t_L g2558 ( 
.A1(n_2095),
.A2(n_1939),
.B(n_1906),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_2202),
.Y(n_2559)
);

OAI21x1_ASAP7_75t_L g2560 ( 
.A1(n_2114),
.A2(n_1950),
.B(n_1941),
.Y(n_2560)
);

OA21x2_ASAP7_75t_L g2561 ( 
.A1(n_2095),
.A2(n_2009),
.B(n_1980),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2135),
.B(n_1682),
.Y(n_2562)
);

INVx4_ASAP7_75t_L g2563 ( 
.A(n_2107),
.Y(n_2563)
);

INVx3_ASAP7_75t_L g2564 ( 
.A(n_2169),
.Y(n_2564)
);

INVx4_ASAP7_75t_L g2565 ( 
.A(n_2107),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2098),
.Y(n_2566)
);

INVx4_ASAP7_75t_L g2567 ( 
.A(n_2107),
.Y(n_2567)
);

BUFx6f_ASAP7_75t_L g2568 ( 
.A(n_2163),
.Y(n_2568)
);

AND2x4_ASAP7_75t_L g2569 ( 
.A(n_2107),
.B(n_1895),
.Y(n_2569)
);

BUFx12f_ASAP7_75t_L g2570 ( 
.A(n_2150),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2163),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2163),
.Y(n_2572)
);

INVx5_ASAP7_75t_L g2573 ( 
.A(n_2139),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2135),
.B(n_1711),
.Y(n_2574)
);

BUFx12f_ASAP7_75t_L g2575 ( 
.A(n_2150),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2098),
.Y(n_2576)
);

OAI22x1_ASAP7_75t_L g2577 ( 
.A1(n_2103),
.A2(n_1369),
.B1(n_1431),
.B2(n_1297),
.Y(n_2577)
);

OA21x2_ASAP7_75t_L g2578 ( 
.A1(n_2095),
.A2(n_2042),
.B(n_2029),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2163),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2135),
.B(n_1711),
.Y(n_2580)
);

BUFx6f_ASAP7_75t_L g2581 ( 
.A(n_2163),
.Y(n_2581)
);

HB1xp67_ASAP7_75t_L g2582 ( 
.A(n_2184),
.Y(n_2582)
);

BUFx12f_ASAP7_75t_L g2583 ( 
.A(n_2150),
.Y(n_2583)
);

BUFx12f_ASAP7_75t_L g2584 ( 
.A(n_2150),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2169),
.B(n_2048),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2135),
.B(n_1745),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2322),
.Y(n_2587)
);

BUFx6f_ASAP7_75t_L g2588 ( 
.A(n_2375),
.Y(n_2588)
);

OA21x2_ASAP7_75t_L g2589 ( 
.A1(n_2401),
.A2(n_2074),
.B(n_2049),
.Y(n_2589)
);

XOR2xp5_ASAP7_75t_L g2590 ( 
.A(n_2263),
.B(n_1313),
.Y(n_2590)
);

OA21x2_ASAP7_75t_L g2591 ( 
.A1(n_2495),
.A2(n_1515),
.B(n_1454),
.Y(n_2591)
);

NOR2xp67_ASAP7_75t_L g2592 ( 
.A(n_2312),
.B(n_1294),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2332),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2379),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_2307),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_2422),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2439),
.Y(n_2597)
);

XNOR2xp5_ASAP7_75t_L g2598 ( 
.A(n_2550),
.B(n_1460),
.Y(n_2598)
);

OAI21x1_ASAP7_75t_L g2599 ( 
.A1(n_2304),
.A2(n_2018),
.B(n_1398),
.Y(n_2599)
);

INVx3_ASAP7_75t_L g2600 ( 
.A(n_2269),
.Y(n_2600)
);

CKINVDCx20_ASAP7_75t_R g2601 ( 
.A(n_2506),
.Y(n_2601)
);

INVx1_ASAP7_75t_SL g2602 ( 
.A(n_2371),
.Y(n_2602)
);

AND2x4_ASAP7_75t_L g2603 ( 
.A(n_2266),
.B(n_1907),
.Y(n_2603)
);

OAI22xp5_ASAP7_75t_SL g2604 ( 
.A1(n_2286),
.A2(n_1493),
.B1(n_1560),
.B2(n_1476),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2346),
.B(n_1745),
.Y(n_2605)
);

AND2x4_ASAP7_75t_L g2606 ( 
.A(n_2300),
.B(n_1966),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2387),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_2321),
.Y(n_2608)
);

AND3x1_ASAP7_75t_L g2609 ( 
.A(n_2339),
.B(n_1649),
.C(n_1644),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2337),
.Y(n_2610)
);

NAND2xp33_ASAP7_75t_R g2611 ( 
.A(n_2271),
.B(n_1314),
.Y(n_2611)
);

CKINVDCx20_ASAP7_75t_R g2612 ( 
.A(n_2327),
.Y(n_2612)
);

CKINVDCx5p33_ASAP7_75t_R g2613 ( 
.A(n_2287),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2295),
.B(n_1325),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2396),
.Y(n_2615)
);

BUFx6f_ASAP7_75t_L g2616 ( 
.A(n_2441),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2397),
.Y(n_2617)
);

BUFx6f_ASAP7_75t_L g2618 ( 
.A(n_2478),
.Y(n_2618)
);

INVx3_ASAP7_75t_L g2619 ( 
.A(n_2428),
.Y(n_2619)
);

BUFx3_ASAP7_75t_L g2620 ( 
.A(n_2493),
.Y(n_2620)
);

CKINVDCx20_ASAP7_75t_R g2621 ( 
.A(n_2288),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2316),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2398),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2400),
.Y(n_2624)
);

BUFx6f_ASAP7_75t_L g2625 ( 
.A(n_2509),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2325),
.B(n_1746),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2317),
.Y(n_2627)
);

CKINVDCx5p33_ASAP7_75t_R g2628 ( 
.A(n_2429),
.Y(n_2628)
);

AND2x2_ASAP7_75t_L g2629 ( 
.A(n_2440),
.B(n_1746),
.Y(n_2629)
);

CKINVDCx5p33_ASAP7_75t_R g2630 ( 
.A(n_2499),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2404),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_2514),
.Y(n_2632)
);

CKINVDCx20_ASAP7_75t_R g2633 ( 
.A(n_2336),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2418),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_R g2635 ( 
.A(n_2278),
.B(n_1295),
.Y(n_2635)
);

CKINVDCx5p33_ASAP7_75t_R g2636 ( 
.A(n_2551),
.Y(n_2636)
);

OAI22xp5_ASAP7_75t_SL g2637 ( 
.A1(n_2369),
.A2(n_2505),
.B1(n_2374),
.B2(n_2413),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2421),
.Y(n_2638)
);

OA21x2_ASAP7_75t_L g2639 ( 
.A1(n_2526),
.A2(n_1301),
.B(n_1299),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2319),
.Y(n_2640)
);

AND2x4_ASAP7_75t_L g2641 ( 
.A(n_2344),
.B(n_1970),
.Y(n_2641)
);

CKINVDCx5p33_ASAP7_75t_R g2642 ( 
.A(n_2570),
.Y(n_2642)
);

CKINVDCx5p33_ASAP7_75t_R g2643 ( 
.A(n_2575),
.Y(n_2643)
);

AND2x6_ASAP7_75t_L g2644 ( 
.A(n_2586),
.B(n_1357),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2297),
.B(n_1377),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2326),
.Y(n_2646)
);

NOR2xp33_ASAP7_75t_L g2647 ( 
.A(n_2324),
.B(n_1380),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2341),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2343),
.Y(n_2649)
);

AND2x2_ASAP7_75t_L g2650 ( 
.A(n_2462),
.B(n_1846),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2351),
.Y(n_2651)
);

OA21x2_ASAP7_75t_L g2652 ( 
.A1(n_2560),
.A2(n_1305),
.B(n_1303),
.Y(n_2652)
);

BUFx2_ASAP7_75t_L g2653 ( 
.A(n_2459),
.Y(n_2653)
);

HB1xp67_ASAP7_75t_L g2654 ( 
.A(n_2355),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2357),
.Y(n_2655)
);

AND2x6_ASAP7_75t_L g2656 ( 
.A(n_2468),
.B(n_1357),
.Y(n_2656)
);

CKINVDCx5p33_ASAP7_75t_R g2657 ( 
.A(n_2583),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2360),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2315),
.Y(n_2659)
);

CKINVDCx5p33_ASAP7_75t_R g2660 ( 
.A(n_2584),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2331),
.B(n_1402),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2368),
.Y(n_2662)
);

CKINVDCx20_ASAP7_75t_R g2663 ( 
.A(n_2294),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2372),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2320),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_SL g2666 ( 
.A(n_2267),
.B(n_1316),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2378),
.Y(n_2667)
);

CKINVDCx5p33_ASAP7_75t_R g2668 ( 
.A(n_2305),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2381),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2487),
.B(n_1846),
.Y(n_2670)
);

INVx3_ASAP7_75t_L g2671 ( 
.A(n_2443),
.Y(n_2671)
);

AND2x2_ASAP7_75t_SL g2672 ( 
.A(n_2542),
.B(n_1391),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2388),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2338),
.Y(n_2674)
);

INVx1_ASAP7_75t_SL g2675 ( 
.A(n_2460),
.Y(n_2675)
);

CKINVDCx20_ASAP7_75t_R g2676 ( 
.A(n_2455),
.Y(n_2676)
);

AND2x4_ASAP7_75t_L g2677 ( 
.A(n_2352),
.B(n_1990),
.Y(n_2677)
);

NOR2xp67_ASAP7_75t_L g2678 ( 
.A(n_2447),
.B(n_1307),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2389),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2463),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2340),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2391),
.Y(n_2682)
);

CKINVDCx5p33_ASAP7_75t_R g2683 ( 
.A(n_2503),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2354),
.Y(n_2684)
);

AND2x4_ASAP7_75t_L g2685 ( 
.A(n_2464),
.B(n_2017),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2364),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2405),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2406),
.Y(n_2688)
);

HB1xp67_ASAP7_75t_L g2689 ( 
.A(n_2390),
.Y(n_2689)
);

BUFx2_ASAP7_75t_L g2690 ( 
.A(n_2520),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2409),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2410),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_2535),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2293),
.B(n_1637),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2411),
.Y(n_2695)
);

XOR2xp5_ASAP7_75t_L g2696 ( 
.A(n_2559),
.B(n_1317),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2318),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2408),
.Y(n_2698)
);

INVxp67_ASAP7_75t_L g2699 ( 
.A(n_2543),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2414),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_2438),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2298),
.Y(n_2702)
);

CKINVDCx5p33_ASAP7_75t_R g2703 ( 
.A(n_2348),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2530),
.B(n_1869),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2301),
.Y(n_2705)
);

CKINVDCx5p33_ASAP7_75t_R g2706 ( 
.A(n_2544),
.Y(n_2706)
);

INVxp67_ASAP7_75t_L g2707 ( 
.A(n_2549),
.Y(n_2707)
);

AND2x4_ASAP7_75t_L g2708 ( 
.A(n_2533),
.B(n_2028),
.Y(n_2708)
);

AND2x4_ASAP7_75t_L g2709 ( 
.A(n_2534),
.B(n_2057),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2329),
.Y(n_2710)
);

CKINVDCx20_ASAP7_75t_R g2711 ( 
.A(n_2469),
.Y(n_2711)
);

HB1xp67_ASAP7_75t_L g2712 ( 
.A(n_2547),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2330),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2334),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2345),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2366),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2273),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2347),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2350),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2353),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2260),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2262),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_2498),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2264),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2349),
.B(n_1843),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2268),
.Y(n_2726)
);

CKINVDCx5p33_ASAP7_75t_R g2727 ( 
.A(n_2502),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2275),
.Y(n_2728)
);

NOR2xp33_ASAP7_75t_SL g2729 ( 
.A(n_2311),
.B(n_1583),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2280),
.Y(n_2730)
);

AND2x4_ASAP7_75t_L g2731 ( 
.A(n_2435),
.B(n_2089),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2281),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2289),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2426),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2349),
.B(n_1915),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2427),
.Y(n_2736)
);

BUFx3_ASAP7_75t_L g2737 ( 
.A(n_2517),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2450),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2475),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2476),
.Y(n_2740)
);

BUFx6f_ASAP7_75t_L g2741 ( 
.A(n_2556),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2477),
.Y(n_2742)
);

BUFx6f_ASAP7_75t_L g2743 ( 
.A(n_2265),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2546),
.B(n_1869),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2486),
.Y(n_2745)
);

INVx4_ASAP7_75t_L g2746 ( 
.A(n_2474),
.Y(n_2746)
);

CKINVDCx20_ASAP7_75t_R g2747 ( 
.A(n_2480),
.Y(n_2747)
);

CKINVDCx5p33_ASAP7_75t_R g2748 ( 
.A(n_2328),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_2361),
.Y(n_2749)
);

INVx3_ASAP7_75t_L g2750 ( 
.A(n_2507),
.Y(n_2750)
);

INVx3_ASAP7_75t_L g2751 ( 
.A(n_2510),
.Y(n_2751)
);

BUFx6f_ASAP7_75t_L g2752 ( 
.A(n_2270),
.Y(n_2752)
);

INVx1_ASAP7_75t_SL g2753 ( 
.A(n_2407),
.Y(n_2753)
);

CKINVDCx5p33_ASAP7_75t_R g2754 ( 
.A(n_2497),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2490),
.Y(n_2755)
);

BUFx6f_ASAP7_75t_L g2756 ( 
.A(n_2276),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2284),
.B(n_1942),
.Y(n_2757)
);

XNOR2xp5_ASAP7_75t_L g2758 ( 
.A(n_2525),
.B(n_1660),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2492),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2552),
.B(n_1933),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2494),
.Y(n_2761)
);

NOR2xp33_ASAP7_75t_L g2762 ( 
.A(n_2536),
.B(n_2541),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2430),
.B(n_1321),
.Y(n_2763)
);

NOR2xp67_ASAP7_75t_L g2764 ( 
.A(n_2573),
.B(n_2291),
.Y(n_2764)
);

INVxp33_ASAP7_75t_L g2765 ( 
.A(n_2279),
.Y(n_2765)
);

OR2x2_ASAP7_75t_L g2766 ( 
.A(n_2282),
.B(n_1680),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2545),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2553),
.Y(n_2768)
);

CKINVDCx20_ASAP7_75t_R g2769 ( 
.A(n_2548),
.Y(n_2769)
);

INVx4_ASAP7_75t_L g2770 ( 
.A(n_2512),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_2555),
.Y(n_2771)
);

NAND2xp33_ASAP7_75t_SL g2772 ( 
.A(n_2306),
.B(n_1318),
.Y(n_2772)
);

OR2x6_ASAP7_75t_L g2773 ( 
.A(n_2385),
.B(n_2417),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2562),
.B(n_1933),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2557),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2566),
.Y(n_2776)
);

CKINVDCx5p33_ASAP7_75t_R g2777 ( 
.A(n_2582),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2576),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2261),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2393),
.Y(n_2780)
);

NAND2x1_ASAP7_75t_L g2781 ( 
.A(n_2333),
.B(n_1357),
.Y(n_2781)
);

NOR2xp33_ASAP7_75t_L g2782 ( 
.A(n_2365),
.B(n_1736),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2292),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2383),
.B(n_1338),
.Y(n_2784)
);

INVxp67_ASAP7_75t_L g2785 ( 
.A(n_2574),
.Y(n_2785)
);

OA21x2_ASAP7_75t_L g2786 ( 
.A1(n_2442),
.A2(n_1353),
.B(n_1343),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2580),
.B(n_1988),
.Y(n_2787)
);

AND2x6_ASAP7_75t_L g2788 ( 
.A(n_2399),
.B(n_1366),
.Y(n_2788)
);

INVx1_ASAP7_75t_SL g2789 ( 
.A(n_2524),
.Y(n_2789)
);

CKINVDCx20_ASAP7_75t_R g2790 ( 
.A(n_2290),
.Y(n_2790)
);

CKINVDCx20_ASAP7_75t_R g2791 ( 
.A(n_2370),
.Y(n_2791)
);

AND2x6_ASAP7_75t_L g2792 ( 
.A(n_2392),
.B(n_1366),
.Y(n_2792)
);

BUFx6f_ASAP7_75t_L g2793 ( 
.A(n_2283),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2412),
.B(n_1354),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2303),
.Y(n_2795)
);

CKINVDCx20_ASAP7_75t_R g2796 ( 
.A(n_2365),
.Y(n_2796)
);

CKINVDCx20_ASAP7_75t_R g2797 ( 
.A(n_2323),
.Y(n_2797)
);

CKINVDCx20_ASAP7_75t_R g2798 ( 
.A(n_2362),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2416),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_SL g2800 ( 
.A(n_2467),
.B(n_1319),
.Y(n_2800)
);

CKINVDCx20_ASAP7_75t_R g2801 ( 
.A(n_2367),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2314),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2419),
.Y(n_2803)
);

BUFx2_ASAP7_75t_L g2804 ( 
.A(n_2529),
.Y(n_2804)
);

BUFx6f_ASAP7_75t_L g2805 ( 
.A(n_2285),
.Y(n_2805)
);

CKINVDCx6p67_ASAP7_75t_R g2806 ( 
.A(n_2573),
.Y(n_2806)
);

CKINVDCx5p33_ASAP7_75t_R g2807 ( 
.A(n_2540),
.Y(n_2807)
);

CKINVDCx5p33_ASAP7_75t_R g2808 ( 
.A(n_2564),
.Y(n_2808)
);

CKINVDCx5p33_ASAP7_75t_R g2809 ( 
.A(n_2424),
.Y(n_2809)
);

AND2x2_ASAP7_75t_L g2810 ( 
.A(n_2420),
.B(n_1988),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_2424),
.Y(n_2811)
);

BUFx3_ASAP7_75t_L g2812 ( 
.A(n_2342),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2356),
.Y(n_2813)
);

CKINVDCx5p33_ASAP7_75t_R g2814 ( 
.A(n_2470),
.Y(n_2814)
);

CKINVDCx20_ASAP7_75t_R g2815 ( 
.A(n_2436),
.Y(n_2815)
);

AND2x6_ASAP7_75t_L g2816 ( 
.A(n_2433),
.B(n_1366),
.Y(n_2816)
);

CKINVDCx5p33_ASAP7_75t_R g2817 ( 
.A(n_2539),
.Y(n_2817)
);

BUFx12f_ASAP7_75t_L g2818 ( 
.A(n_2563),
.Y(n_2818)
);

BUFx6f_ASAP7_75t_L g2819 ( 
.A(n_2299),
.Y(n_2819)
);

BUFx6f_ASAP7_75t_L g2820 ( 
.A(n_2302),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2358),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2359),
.Y(n_2822)
);

CKINVDCx5p33_ASAP7_75t_R g2823 ( 
.A(n_2565),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2432),
.Y(n_2824)
);

CKINVDCx20_ASAP7_75t_R g2825 ( 
.A(n_2484),
.Y(n_2825)
);

CKINVDCx20_ASAP7_75t_R g2826 ( 
.A(n_2567),
.Y(n_2826)
);

INVx3_ASAP7_75t_L g2827 ( 
.A(n_2380),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2377),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2373),
.Y(n_2829)
);

CKINVDCx5p33_ASAP7_75t_R g2830 ( 
.A(n_2516),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2481),
.B(n_1361),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2511),
.B(n_1378),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2585),
.Y(n_2833)
);

CKINVDCx5p33_ASAP7_75t_R g2834 ( 
.A(n_2310),
.Y(n_2834)
);

CKINVDCx5p33_ASAP7_75t_R g2835 ( 
.A(n_2384),
.Y(n_2835)
);

BUFx4f_ASAP7_75t_L g2836 ( 
.A(n_2402),
.Y(n_2836)
);

INVx1_ASAP7_75t_SL g2837 ( 
.A(n_2277),
.Y(n_2837)
);

AND2x4_ASAP7_75t_L g2838 ( 
.A(n_2425),
.B(n_1816),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2515),
.B(n_1381),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2444),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2456),
.Y(n_2841)
);

BUFx6f_ASAP7_75t_L g2842 ( 
.A(n_2308),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2446),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2415),
.B(n_1384),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2457),
.Y(n_2845)
);

AND2x4_ASAP7_75t_L g2846 ( 
.A(n_2448),
.B(n_1845),
.Y(n_2846)
);

CKINVDCx5p33_ASAP7_75t_R g2847 ( 
.A(n_2395),
.Y(n_2847)
);

BUFx6f_ASAP7_75t_L g2848 ( 
.A(n_2423),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2458),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_SL g2850 ( 
.A(n_2471),
.B(n_1322),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2466),
.Y(n_2851)
);

CKINVDCx5p33_ASAP7_75t_R g2852 ( 
.A(n_2394),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2449),
.Y(n_2853)
);

CKINVDCx5p33_ASAP7_75t_R g2854 ( 
.A(n_2402),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2479),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2518),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2523),
.B(n_1389),
.Y(n_2857)
);

CKINVDCx5p33_ASAP7_75t_R g2858 ( 
.A(n_2482),
.Y(n_2858)
);

BUFx6f_ASAP7_75t_L g2859 ( 
.A(n_2431),
.Y(n_2859)
);

CKINVDCx20_ASAP7_75t_R g2860 ( 
.A(n_2472),
.Y(n_2860)
);

CKINVDCx5p33_ASAP7_75t_R g2861 ( 
.A(n_2488),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2451),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2527),
.Y(n_2863)
);

INVx2_ASAP7_75t_SL g2864 ( 
.A(n_2537),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2272),
.Y(n_2865)
);

BUFx6f_ASAP7_75t_L g2866 ( 
.A(n_2437),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_R g2867 ( 
.A(n_2313),
.B(n_1396),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2274),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2335),
.B(n_2554),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2296),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2434),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2558),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2561),
.Y(n_2873)
);

INVx3_ASAP7_75t_L g2874 ( 
.A(n_2445),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2569),
.B(n_1397),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2578),
.Y(n_2876)
);

OAI21x1_ASAP7_75t_L g2877 ( 
.A1(n_2454),
.A2(n_1523),
.B(n_1464),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2363),
.B(n_2069),
.Y(n_2878)
);

CKINVDCx5p33_ASAP7_75t_R g2879 ( 
.A(n_2382),
.Y(n_2879)
);

BUFx6f_ASAP7_75t_L g2880 ( 
.A(n_2452),
.Y(n_2880)
);

CKINVDCx5p33_ASAP7_75t_R g2881 ( 
.A(n_2386),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2465),
.Y(n_2882)
);

INVx4_ASAP7_75t_L g2883 ( 
.A(n_2376),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2473),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2483),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2496),
.Y(n_2886)
);

CKINVDCx5p33_ASAP7_75t_R g2887 ( 
.A(n_2577),
.Y(n_2887)
);

HB1xp67_ASAP7_75t_L g2888 ( 
.A(n_2403),
.Y(n_2888)
);

CKINVDCx20_ASAP7_75t_R g2889 ( 
.A(n_2309),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2513),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2522),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2531),
.Y(n_2892)
);

OA21x2_ASAP7_75t_L g2893 ( 
.A1(n_2571),
.A2(n_1413),
.B(n_1407),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2572),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2579),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2453),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2461),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2485),
.Y(n_2898)
);

INVx2_ASAP7_75t_L g2899 ( 
.A(n_2622),
.Y(n_2899)
);

INVx3_ASAP7_75t_L g2900 ( 
.A(n_2588),
.Y(n_2900)
);

NAND2xp33_ASAP7_75t_SL g2901 ( 
.A(n_2661),
.B(n_1323),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2627),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2721),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2640),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2722),
.Y(n_2905)
);

INVx4_ASAP7_75t_L g2906 ( 
.A(n_2588),
.Y(n_2906)
);

NAND3xp33_ASAP7_75t_L g2907 ( 
.A(n_2748),
.B(n_1335),
.C(n_1331),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_SL g2908 ( 
.A(n_2668),
.B(n_1339),
.Y(n_2908)
);

NAND3xp33_ASAP7_75t_L g2909 ( 
.A(n_2749),
.B(n_1347),
.C(n_1345),
.Y(n_2909)
);

INVx8_ASAP7_75t_L g2910 ( 
.A(n_2773),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_L g2911 ( 
.A(n_2602),
.B(n_1733),
.Y(n_2911)
);

NOR2xp33_ASAP7_75t_L g2912 ( 
.A(n_2701),
.B(n_1768),
.Y(n_2912)
);

INVx3_ASAP7_75t_L g2913 ( 
.A(n_2620),
.Y(n_2913)
);

INVxp33_ASAP7_75t_SL g2914 ( 
.A(n_2680),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_SL g2915 ( 
.A(n_2836),
.B(n_1349),
.Y(n_2915)
);

BUFx3_ASAP7_75t_L g2916 ( 
.A(n_2633),
.Y(n_2916)
);

XOR2xp5_ASAP7_75t_R g2917 ( 
.A(n_2601),
.B(n_2608),
.Y(n_2917)
);

INVx4_ASAP7_75t_L g2918 ( 
.A(n_2613),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_2814),
.B(n_1351),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2647),
.B(n_2757),
.Y(n_2920)
);

INVx3_ASAP7_75t_L g2921 ( 
.A(n_2737),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2646),
.Y(n_2922)
);

HB1xp67_ASAP7_75t_L g2923 ( 
.A(n_2675),
.Y(n_2923)
);

OAI22xp5_ASAP7_75t_L g2924 ( 
.A1(n_2609),
.A2(n_1429),
.B1(n_1382),
.B2(n_1355),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_SL g2925 ( 
.A(n_2817),
.B(n_1352),
.Y(n_2925)
);

INVx2_ASAP7_75t_SL g2926 ( 
.A(n_2653),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2674),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2833),
.B(n_1892),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2681),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2724),
.Y(n_2930)
);

AOI21x1_ASAP7_75t_L g2931 ( 
.A1(n_2865),
.A2(n_1675),
.B(n_1665),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2684),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2686),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2690),
.B(n_2069),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2594),
.Y(n_2935)
);

NOR2xp33_ASAP7_75t_L g2936 ( 
.A(n_2699),
.B(n_1769),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2840),
.B(n_1949),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2726),
.Y(n_2938)
);

OR2x6_ASAP7_75t_L g2939 ( 
.A(n_2773),
.B(n_2052),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2730),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2607),
.Y(n_2941)
);

BUFx2_ASAP7_75t_L g2942 ( 
.A(n_2612),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2615),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2732),
.Y(n_2944)
);

AND3x2_ASAP7_75t_L g2945 ( 
.A(n_2707),
.B(n_1531),
.C(n_1529),
.Y(n_2945)
);

OR2x2_ASAP7_75t_L g2946 ( 
.A(n_2753),
.B(n_2766),
.Y(n_2946)
);

BUFx3_ASAP7_75t_L g2947 ( 
.A(n_2889),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2733),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2617),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2623),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2624),
.Y(n_2951)
);

OR2x2_ASAP7_75t_SL g2952 ( 
.A(n_2689),
.B(n_1549),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2734),
.Y(n_2953)
);

INVx5_ASAP7_75t_L g2954 ( 
.A(n_2818),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2631),
.Y(n_2955)
);

AO22x2_ASAP7_75t_L g2956 ( 
.A1(n_2590),
.A2(n_1803),
.B1(n_1806),
.B2(n_1795),
.Y(n_2956)
);

NOR2xp33_ASAP7_75t_L g2957 ( 
.A(n_2785),
.B(n_1829),
.Y(n_2957)
);

BUFx6f_ASAP7_75t_L g2958 ( 
.A(n_2616),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2810),
.B(n_2088),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2634),
.Y(n_2960)
);

AOI22xp33_ASAP7_75t_L g2961 ( 
.A1(n_2637),
.A2(n_1928),
.B1(n_2007),
.B2(n_1913),
.Y(n_2961)
);

AO22x2_ASAP7_75t_L g2962 ( 
.A1(n_2696),
.A2(n_2020),
.B1(n_2085),
.B2(n_1685),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2638),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2736),
.Y(n_2964)
);

NAND3xp33_ASAP7_75t_L g2965 ( 
.A(n_2611),
.B(n_1362),
.C(n_1358),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2739),
.Y(n_2966)
);

BUFx3_ASAP7_75t_L g2967 ( 
.A(n_2663),
.Y(n_2967)
);

NAND2xp33_ASAP7_75t_L g2968 ( 
.A(n_2823),
.B(n_1367),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2719),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2659),
.Y(n_2970)
);

BUFx6f_ASAP7_75t_L g2971 ( 
.A(n_2616),
.Y(n_2971)
);

AOI22xp5_ASAP7_75t_L g2972 ( 
.A1(n_2841),
.A2(n_1427),
.B1(n_1428),
.B2(n_1419),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2665),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2779),
.Y(n_2974)
);

NAND3xp33_ASAP7_75t_L g2975 ( 
.A(n_2807),
.B(n_1373),
.C(n_1370),
.Y(n_2975)
);

INVx4_ASAP7_75t_L g2976 ( 
.A(n_2628),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2783),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2740),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2795),
.Y(n_2979)
);

INVx4_ASAP7_75t_L g2980 ( 
.A(n_2630),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2802),
.Y(n_2981)
);

BUFx6f_ASAP7_75t_L g2982 ( 
.A(n_2618),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2824),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2843),
.Y(n_2984)
);

INVx3_ASAP7_75t_L g2985 ( 
.A(n_2618),
.Y(n_2985)
);

NOR2xp33_ASAP7_75t_L g2986 ( 
.A(n_2614),
.B(n_1383),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2853),
.Y(n_2987)
);

INVx2_ASAP7_75t_SL g2988 ( 
.A(n_2654),
.Y(n_2988)
);

OAI22x1_ASAP7_75t_L g2989 ( 
.A1(n_2598),
.A2(n_2758),
.B1(n_2706),
.B2(n_2754),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2845),
.B(n_1976),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2742),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_SL g2992 ( 
.A(n_2808),
.B(n_1386),
.Y(n_2992)
);

AOI22xp33_ASAP7_75t_L g2993 ( 
.A1(n_2702),
.A2(n_1611),
.B1(n_1654),
.B2(n_1570),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2862),
.Y(n_2994)
);

INVxp33_ASAP7_75t_L g2995 ( 
.A(n_2635),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2884),
.Y(n_2996)
);

INVx1_ASAP7_75t_SL g2997 ( 
.A(n_2815),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2894),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2728),
.Y(n_2999)
);

AOI22xp33_ASAP7_75t_L g3000 ( 
.A1(n_2705),
.A2(n_1741),
.B1(n_1763),
.B2(n_1702),
.Y(n_3000)
);

INVx2_ASAP7_75t_SL g3001 ( 
.A(n_2605),
.Y(n_3001)
);

BUFx6f_ASAP7_75t_L g3002 ( 
.A(n_2625),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2745),
.Y(n_3003)
);

AOI22xp33_ASAP7_75t_SL g3004 ( 
.A1(n_2672),
.A2(n_2088),
.B1(n_1390),
.B2(n_1394),
.Y(n_3004)
);

AOI21x1_ASAP7_75t_L g3005 ( 
.A1(n_2868),
.A2(n_1688),
.B(n_1681),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2738),
.Y(n_3006)
);

BUFx3_ASAP7_75t_L g3007 ( 
.A(n_2676),
.Y(n_3007)
);

INVx3_ASAP7_75t_L g3008 ( 
.A(n_2625),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2755),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2759),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_SL g3011 ( 
.A(n_2784),
.B(n_1387),
.Y(n_3011)
);

AO21x2_ASAP7_75t_L g3012 ( 
.A1(n_2829),
.A2(n_1696),
.B(n_1691),
.Y(n_3012)
);

CKINVDCx5p33_ASAP7_75t_R g3013 ( 
.A(n_2683),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_L g3014 ( 
.A(n_2645),
.B(n_2849),
.Y(n_3014)
);

NAND2xp33_ASAP7_75t_SL g3015 ( 
.A(n_2693),
.B(n_1401),
.Y(n_3015)
);

NOR2xp33_ASAP7_75t_L g3016 ( 
.A(n_2851),
.B(n_1403),
.Y(n_3016)
);

OAI22xp33_ASAP7_75t_L g3017 ( 
.A1(n_2729),
.A2(n_1405),
.B1(n_1406),
.B2(n_1404),
.Y(n_3017)
);

AOI22xp5_ASAP7_75t_L g3018 ( 
.A1(n_2855),
.A2(n_1450),
.B1(n_1459),
.B2(n_1436),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_SL g3019 ( 
.A(n_2746),
.B(n_1408),
.Y(n_3019)
);

OR2x6_ASAP7_75t_L g3020 ( 
.A(n_2864),
.B(n_2489),
.Y(n_3020)
);

AND2x2_ASAP7_75t_L g3021 ( 
.A(n_2771),
.B(n_2491),
.Y(n_3021)
);

NOR2xp33_ASAP7_75t_L g3022 ( 
.A(n_2856),
.B(n_1409),
.Y(n_3022)
);

NOR2xp33_ASAP7_75t_L g3023 ( 
.A(n_2863),
.B(n_1410),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_SL g3024 ( 
.A(n_2770),
.B(n_1414),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2761),
.Y(n_3025)
);

NAND2xp33_ASAP7_75t_L g3026 ( 
.A(n_2809),
.B(n_1415),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2768),
.Y(n_3027)
);

INVx3_ASAP7_75t_L g3028 ( 
.A(n_2741),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2844),
.B(n_1976),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2767),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2776),
.Y(n_3031)
);

OR2x6_ASAP7_75t_L g3032 ( 
.A(n_2712),
.B(n_2741),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2775),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_SL g3034 ( 
.A(n_2811),
.B(n_1416),
.Y(n_3034)
);

BUFx10_ASAP7_75t_L g3035 ( 
.A(n_2595),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2778),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2710),
.B(n_1978),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2713),
.Y(n_3038)
);

NAND3xp33_ASAP7_75t_L g3039 ( 
.A(n_2777),
.B(n_1421),
.C(n_1418),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2717),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2714),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2715),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2718),
.B(n_1978),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2720),
.Y(n_3044)
);

NAND2xp33_ASAP7_75t_L g3045 ( 
.A(n_2854),
.B(n_1422),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2882),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2885),
.Y(n_3047)
);

BUFx6f_ASAP7_75t_L g3048 ( 
.A(n_2743),
.Y(n_3048)
);

BUFx6f_ASAP7_75t_L g3049 ( 
.A(n_2743),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2698),
.Y(n_3050)
);

INVx4_ASAP7_75t_L g3051 ( 
.A(n_2632),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2700),
.Y(n_3052)
);

INVx4_ASAP7_75t_L g3053 ( 
.A(n_2636),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2886),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2762),
.B(n_1978),
.Y(n_3055)
);

AND2x2_ASAP7_75t_SL g3056 ( 
.A(n_2626),
.B(n_1764),
.Y(n_3056)
);

NOR2xp33_ASAP7_75t_L g3057 ( 
.A(n_2666),
.B(n_1423),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2890),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2891),
.Y(n_3059)
);

INVx2_ASAP7_75t_SL g3060 ( 
.A(n_2731),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_2892),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2895),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2813),
.Y(n_3063)
);

AND2x2_ASAP7_75t_SL g3064 ( 
.A(n_2629),
.B(n_1811),
.Y(n_3064)
);

NOR2xp33_ASAP7_75t_L g3065 ( 
.A(n_2837),
.B(n_1424),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2821),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_2822),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2697),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2716),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2831),
.B(n_2026),
.Y(n_3070)
);

OAI22xp33_ASAP7_75t_L g3071 ( 
.A1(n_2828),
.A2(n_1433),
.B1(n_1434),
.B2(n_1425),
.Y(n_3071)
);

AND2x2_ASAP7_75t_L g3072 ( 
.A(n_2650),
.B(n_2500),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2877),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2870),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2871),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2780),
.Y(n_3076)
);

OA22x2_ASAP7_75t_L g3077 ( 
.A1(n_2604),
.A2(n_1441),
.B1(n_1446),
.B2(n_1439),
.Y(n_3077)
);

AND3x2_ASAP7_75t_L g3078 ( 
.A(n_2670),
.B(n_1840),
.C(n_1817),
.Y(n_3078)
);

OAI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_2827),
.A2(n_2839),
.B1(n_2832),
.B2(n_2763),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2725),
.B(n_2026),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2799),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_SL g3082 ( 
.A(n_2789),
.B(n_1447),
.Y(n_3082)
);

NOR2x1p5_ASAP7_75t_L g3083 ( 
.A(n_2806),
.B(n_1449),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2872),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2735),
.B(n_2026),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2857),
.B(n_2072),
.Y(n_3086)
);

AO21x2_ASAP7_75t_L g3087 ( 
.A1(n_2873),
.A2(n_1707),
.B(n_1699),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2803),
.Y(n_3088)
);

INVxp33_ASAP7_75t_SL g3089 ( 
.A(n_2596),
.Y(n_3089)
);

INVx5_ASAP7_75t_L g3090 ( 
.A(n_2644),
.Y(n_3090)
);

INVx4_ASAP7_75t_L g3091 ( 
.A(n_2642),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_2876),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2812),
.Y(n_3093)
);

INVx1_ASAP7_75t_SL g3094 ( 
.A(n_2711),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2587),
.Y(n_3095)
);

BUFx3_ASAP7_75t_L g3096 ( 
.A(n_2621),
.Y(n_3096)
);

INVx2_ASAP7_75t_SL g3097 ( 
.A(n_2704),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_SL g3098 ( 
.A(n_2592),
.B(n_1452),
.Y(n_3098)
);

BUFx2_ASAP7_75t_L g3099 ( 
.A(n_2747),
.Y(n_3099)
);

BUFx6f_ASAP7_75t_SL g3100 ( 
.A(n_2603),
.Y(n_3100)
);

BUFx10_ASAP7_75t_L g3101 ( 
.A(n_2597),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2593),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2694),
.B(n_2072),
.Y(n_3103)
);

INVx3_ASAP7_75t_L g3104 ( 
.A(n_2752),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2591),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_SL g3106 ( 
.A(n_2804),
.B(n_2678),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2610),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2648),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2589),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2649),
.Y(n_3110)
);

INVx2_ASAP7_75t_SL g3111 ( 
.A(n_2744),
.Y(n_3111)
);

AO22x2_ASAP7_75t_L g3112 ( 
.A1(n_2765),
.A2(n_1709),
.B1(n_1713),
.B2(n_1708),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2651),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2655),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2658),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2662),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2664),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2667),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2669),
.Y(n_3119)
);

OR2x2_ASAP7_75t_L g3120 ( 
.A(n_2869),
.B(n_1722),
.Y(n_3120)
);

INVx4_ASAP7_75t_L g3121 ( 
.A(n_2643),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_2673),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_SL g3123 ( 
.A(n_2760),
.B(n_1455),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2679),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2788),
.B(n_2644),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_SL g3126 ( 
.A(n_2774),
.B(n_1456),
.Y(n_3126)
);

INVx4_ASAP7_75t_L g3127 ( 
.A(n_2657),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2682),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2687),
.Y(n_3129)
);

INVx2_ASAP7_75t_SL g3130 ( 
.A(n_2787),
.Y(n_3130)
);

INVx2_ASAP7_75t_SL g3131 ( 
.A(n_2858),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2688),
.Y(n_3132)
);

INVx2_ASAP7_75t_SL g3133 ( 
.A(n_2861),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2788),
.B(n_2072),
.Y(n_3134)
);

BUFx3_ASAP7_75t_L g3135 ( 
.A(n_2826),
.Y(n_3135)
);

OAI22xp5_ASAP7_75t_L g3136 ( 
.A1(n_2794),
.A2(n_1466),
.B1(n_1469),
.B2(n_1457),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2691),
.Y(n_3137)
);

INVx3_ASAP7_75t_L g3138 ( 
.A(n_2752),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2692),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2920),
.B(n_2788),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_3014),
.B(n_2879),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_SL g3142 ( 
.A(n_2988),
.B(n_2881),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2903),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2905),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2986),
.B(n_2644),
.Y(n_3145)
);

AO221x1_ASAP7_75t_L g3146 ( 
.A1(n_3017),
.A2(n_2671),
.B1(n_2750),
.B2(n_2619),
.C(n_2600),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_3016),
.B(n_2656),
.Y(n_3147)
);

OR2x6_ASAP7_75t_L g3148 ( 
.A(n_2910),
.B(n_2606),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_SL g3149 ( 
.A(n_2926),
.B(n_2769),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_3040),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2899),
.Y(n_3151)
);

INVx2_ASAP7_75t_SL g3152 ( 
.A(n_2923),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_3022),
.B(n_2656),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_3023),
.B(n_2656),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_2902),
.Y(n_3155)
);

AND2x6_ASAP7_75t_SL g3156 ( 
.A(n_2917),
.B(n_2797),
.Y(n_3156)
);

BUFx8_ASAP7_75t_L g3157 ( 
.A(n_3100),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2904),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2930),
.B(n_2751),
.Y(n_3159)
);

NOR2xp33_ASAP7_75t_L g3160 ( 
.A(n_2914),
.B(n_2860),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2938),
.B(n_2782),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2940),
.B(n_2878),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2944),
.B(n_2792),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_SL g3164 ( 
.A(n_3013),
.B(n_2875),
.Y(n_3164)
);

NOR2xp67_ASAP7_75t_L g3165 ( 
.A(n_2918),
.B(n_2660),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2922),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2927),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2948),
.B(n_2792),
.Y(n_3168)
);

INVx3_ASAP7_75t_L g3169 ( 
.A(n_3135),
.Y(n_3169)
);

AO221x1_ASAP7_75t_L g3170 ( 
.A1(n_2962),
.A2(n_2695),
.B1(n_1735),
.B2(n_1747),
.C(n_1739),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2953),
.Y(n_3171)
);

AND2x2_ASAP7_75t_L g3172 ( 
.A(n_2911),
.B(n_2838),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2929),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2964),
.Y(n_3174)
);

NAND3xp33_ASAP7_75t_L g3175 ( 
.A(n_2912),
.B(n_2772),
.C(n_2850),
.Y(n_3175)
);

BUFx5_ASAP7_75t_L g3176 ( 
.A(n_3063),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_SL g3177 ( 
.A(n_2995),
.B(n_2764),
.Y(n_3177)
);

NOR2xp33_ASAP7_75t_L g3178 ( 
.A(n_3056),
.B(n_2796),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2966),
.B(n_2792),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_2936),
.B(n_3064),
.Y(n_3180)
);

NOR3xp33_ASAP7_75t_L g3181 ( 
.A(n_3015),
.B(n_2800),
.C(n_1750),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2978),
.Y(n_3182)
);

BUFx6f_ASAP7_75t_L g3183 ( 
.A(n_3048),
.Y(n_3183)
);

NOR2xp33_ASAP7_75t_L g3184 ( 
.A(n_3094),
.B(n_2791),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_2991),
.B(n_2816),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_3003),
.B(n_2816),
.Y(n_3186)
);

HB1xp67_ASAP7_75t_L g3187 ( 
.A(n_2997),
.Y(n_3187)
);

NAND2xp33_ASAP7_75t_SL g3188 ( 
.A(n_2976),
.B(n_2790),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_SL g3189 ( 
.A(n_3001),
.B(n_2641),
.Y(n_3189)
);

NOR2xp33_ASAP7_75t_L g3190 ( 
.A(n_3097),
.B(n_2846),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_3111),
.B(n_2703),
.Y(n_3191)
);

NOR2xp33_ASAP7_75t_L g3192 ( 
.A(n_3130),
.B(n_2677),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_2959),
.B(n_2685),
.Y(n_3193)
);

BUFx6f_ASAP7_75t_SL g3194 ( 
.A(n_2916),
.Y(n_3194)
);

NOR2xp33_ASAP7_75t_L g3195 ( 
.A(n_2946),
.B(n_2708),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_3009),
.B(n_2816),
.Y(n_3196)
);

NOR2xp33_ASAP7_75t_L g3197 ( 
.A(n_2957),
.B(n_2709),
.Y(n_3197)
);

NOR2xp33_ASAP7_75t_L g3198 ( 
.A(n_3065),
.B(n_2887),
.Y(n_3198)
);

NOR2xp33_ASAP7_75t_L g3199 ( 
.A(n_3099),
.B(n_2825),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_2932),
.Y(n_3200)
);

AO21x2_ASAP7_75t_L g3201 ( 
.A1(n_3105),
.A2(n_2599),
.B(n_2639),
.Y(n_3201)
);

HB1xp67_ASAP7_75t_L g3202 ( 
.A(n_2942),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_3030),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2933),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3031),
.B(n_2786),
.Y(n_3205)
);

NOR2xp33_ASAP7_75t_L g3206 ( 
.A(n_3123),
.B(n_2723),
.Y(n_3206)
);

INVx2_ASAP7_75t_L g3207 ( 
.A(n_2969),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_2999),
.Y(n_3208)
);

BUFx3_ASAP7_75t_L g3209 ( 
.A(n_2967),
.Y(n_3209)
);

BUFx2_ASAP7_75t_R g3210 ( 
.A(n_3007),
.Y(n_3210)
);

AND2x2_ASAP7_75t_L g3211 ( 
.A(n_2934),
.B(n_2727),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_3036),
.B(n_2893),
.Y(n_3212)
);

NOR2xp33_ASAP7_75t_L g3213 ( 
.A(n_3126),
.B(n_2834),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3038),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3041),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_3042),
.B(n_1730),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_3006),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_3044),
.B(n_1754),
.Y(n_3218)
);

NOR3xp33_ASAP7_75t_L g3219 ( 
.A(n_3039),
.B(n_1759),
.C(n_1756),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_3010),
.Y(n_3220)
);

BUFx6f_ASAP7_75t_L g3221 ( 
.A(n_3048),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_3050),
.B(n_1776),
.Y(n_3222)
);

A2O1A1Ixp33_ASAP7_75t_L g3223 ( 
.A1(n_3057),
.A2(n_1801),
.B(n_1819),
.C(n_1785),
.Y(n_3223)
);

A2O1A1Ixp33_ASAP7_75t_L g3224 ( 
.A1(n_2961),
.A2(n_1822),
.B(n_1823),
.C(n_1821),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3052),
.Y(n_3225)
);

NAND2xp33_ASAP7_75t_L g3226 ( 
.A(n_3079),
.B(n_1470),
.Y(n_3226)
);

NOR3xp33_ASAP7_75t_L g3227 ( 
.A(n_2907),
.B(n_1836),
.C(n_1833),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_SL g3228 ( 
.A(n_3004),
.B(n_2867),
.Y(n_3228)
);

NOR2xp33_ASAP7_75t_L g3229 ( 
.A(n_3131),
.B(n_2798),
.Y(n_3229)
);

NOR2xp33_ASAP7_75t_L g3230 ( 
.A(n_3133),
.B(n_2801),
.Y(n_3230)
);

NOR2xp33_ASAP7_75t_L g3231 ( 
.A(n_2952),
.B(n_3011),
.Y(n_3231)
);

BUFx6f_ASAP7_75t_L g3232 ( 
.A(n_3049),
.Y(n_3232)
);

NOR2xp33_ASAP7_75t_L g3233 ( 
.A(n_2908),
.B(n_2896),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3025),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3027),
.Y(n_3235)
);

NAND2xp33_ASAP7_75t_L g3236 ( 
.A(n_3029),
.B(n_1473),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3033),
.Y(n_3237)
);

NOR2xp67_ASAP7_75t_L g3238 ( 
.A(n_2980),
.B(n_2888),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2935),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_SL g3240 ( 
.A(n_2913),
.B(n_1474),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_2928),
.B(n_1839),
.Y(n_3241)
);

NAND2xp33_ASAP7_75t_L g3242 ( 
.A(n_2901),
.B(n_1479),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2941),
.Y(n_3243)
);

OR2x6_ASAP7_75t_L g3244 ( 
.A(n_2910),
.B(n_2756),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_SL g3245 ( 
.A(n_2921),
.B(n_1485),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2937),
.B(n_1842),
.Y(n_3246)
);

NOR2xp33_ASAP7_75t_L g3247 ( 
.A(n_3060),
.B(n_2898),
.Y(n_3247)
);

AND2x2_ASAP7_75t_SL g3248 ( 
.A(n_3051),
.B(n_2756),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_SL g3249 ( 
.A(n_2958),
.B(n_1486),
.Y(n_3249)
);

NOR2xp33_ASAP7_75t_L g3250 ( 
.A(n_3089),
.B(n_2897),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_2943),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2949),
.B(n_1848),
.Y(n_3252)
);

INVxp67_ASAP7_75t_L g3253 ( 
.A(n_3021),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_SL g3254 ( 
.A(n_2958),
.B(n_1488),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_3072),
.B(n_2874),
.Y(n_3255)
);

NOR2xp33_ASAP7_75t_L g3256 ( 
.A(n_2992),
.B(n_1491),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_SL g3257 ( 
.A(n_2971),
.B(n_1495),
.Y(n_3257)
);

NAND2x1p5_ASAP7_75t_L g3258 ( 
.A(n_2906),
.B(n_2793),
.Y(n_3258)
);

AND2x2_ASAP7_75t_L g3259 ( 
.A(n_3112),
.B(n_2793),
.Y(n_3259)
);

NAND2xp33_ASAP7_75t_L g3260 ( 
.A(n_3070),
.B(n_2975),
.Y(n_3260)
);

AOI22xp5_ASAP7_75t_L g3261 ( 
.A1(n_2968),
.A2(n_1498),
.B1(n_1500),
.B2(n_1496),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2950),
.Y(n_3262)
);

NOR3xp33_ASAP7_75t_L g3263 ( 
.A(n_2909),
.B(n_1853),
.C(n_1849),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_2951),
.B(n_1859),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_2955),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_2960),
.B(n_1871),
.Y(n_3266)
);

INVxp67_ASAP7_75t_L g3267 ( 
.A(n_3096),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_2989),
.B(n_2805),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2963),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3055),
.B(n_1874),
.Y(n_3270)
);

AND2x2_ASAP7_75t_L g3271 ( 
.A(n_3120),
.B(n_2805),
.Y(n_3271)
);

INVxp33_ASAP7_75t_L g3272 ( 
.A(n_3049),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_3076),
.B(n_1889),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_3081),
.B(n_1893),
.Y(n_3274)
);

XNOR2xp5_ASAP7_75t_L g3275 ( 
.A(n_2947),
.B(n_2852),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3088),
.Y(n_3276)
);

CKINVDCx5p33_ASAP7_75t_R g3277 ( 
.A(n_3035),
.Y(n_3277)
);

NOR2xp33_ASAP7_75t_L g3278 ( 
.A(n_3068),
.B(n_1503),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3046),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_2970),
.Y(n_3280)
);

INVxp33_ASAP7_75t_L g3281 ( 
.A(n_2971),
.Y(n_3281)
);

NOR2xp33_ASAP7_75t_L g3282 ( 
.A(n_3069),
.B(n_1505),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_2919),
.B(n_1509),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_SL g3284 ( 
.A(n_2982),
.B(n_1510),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3047),
.Y(n_3285)
);

AOI22xp33_ASAP7_75t_L g3286 ( 
.A1(n_3012),
.A2(n_2652),
.B1(n_1968),
.B2(n_2015),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3066),
.B(n_1894),
.Y(n_3287)
);

NOR2xp33_ASAP7_75t_L g3288 ( 
.A(n_2925),
.B(n_1511),
.Y(n_3288)
);

NOR2xp33_ASAP7_75t_L g3289 ( 
.A(n_3082),
.B(n_1514),
.Y(n_3289)
);

INVx1_ASAP7_75t_SL g3290 ( 
.A(n_3032),
.Y(n_3290)
);

INVx5_ASAP7_75t_L g3291 ( 
.A(n_3101),
.Y(n_3291)
);

BUFx5_ASAP7_75t_L g3292 ( 
.A(n_3093),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3067),
.B(n_1898),
.Y(n_3293)
);

NOR2xp33_ASAP7_75t_L g3294 ( 
.A(n_2900),
.B(n_1520),
.Y(n_3294)
);

NOR2xp33_ASAP7_75t_L g3295 ( 
.A(n_3034),
.B(n_1521),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3143),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3144),
.Y(n_3297)
);

AND2x2_ASAP7_75t_L g3298 ( 
.A(n_3180),
.B(n_3032),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3171),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3174),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_3197),
.B(n_2972),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3141),
.B(n_3018),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_3198),
.B(n_3136),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3251),
.Y(n_3304)
);

AND2x4_ASAP7_75t_L g3305 ( 
.A(n_3244),
.B(n_2954),
.Y(n_3305)
);

AO22x2_ASAP7_75t_L g3306 ( 
.A1(n_3259),
.A2(n_2924),
.B1(n_3114),
.B2(n_3108),
.Y(n_3306)
);

AND2x4_ASAP7_75t_L g3307 ( 
.A(n_3244),
.B(n_2954),
.Y(n_3307)
);

NAND2x1p5_ASAP7_75t_L g3308 ( 
.A(n_3209),
.B(n_3053),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3182),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3203),
.B(n_3045),
.Y(n_3310)
);

NOR2xp33_ASAP7_75t_L g3311 ( 
.A(n_3172),
.B(n_3091),
.Y(n_3311)
);

AO22x2_ASAP7_75t_L g3312 ( 
.A1(n_3228),
.A2(n_3119),
.B1(n_3124),
.B2(n_3118),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3214),
.B(n_2973),
.Y(n_3313)
);

AND2x4_ASAP7_75t_L g3314 ( 
.A(n_3148),
.B(n_3121),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3265),
.Y(n_3315)
);

AO22x2_ASAP7_75t_L g3316 ( 
.A1(n_3268),
.A2(n_3128),
.B1(n_3110),
.B2(n_3115),
.Y(n_3316)
);

OAI22xp33_ASAP7_75t_SL g3317 ( 
.A1(n_3253),
.A2(n_2939),
.B1(n_2956),
.B2(n_2835),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3215),
.Y(n_3318)
);

AO22x2_ASAP7_75t_L g3319 ( 
.A1(n_3239),
.A2(n_3113),
.B1(n_3117),
.B2(n_3116),
.Y(n_3319)
);

OAI221xp5_ASAP7_75t_L g3320 ( 
.A1(n_3224),
.A2(n_2965),
.B1(n_3127),
.B2(n_3077),
.C(n_2939),
.Y(n_3320)
);

AOI22xp5_ASAP7_75t_L g3321 ( 
.A1(n_3160),
.A2(n_3026),
.B1(n_3071),
.B2(n_2982),
.Y(n_3321)
);

INVxp67_ASAP7_75t_L g3322 ( 
.A(n_3152),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_3150),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3225),
.Y(n_3324)
);

BUFx8_ASAP7_75t_L g3325 ( 
.A(n_3194),
.Y(n_3325)
);

NOR2xp67_ASAP7_75t_L g3326 ( 
.A(n_3291),
.B(n_3090),
.Y(n_3326)
);

AO22x2_ASAP7_75t_L g3327 ( 
.A1(n_3243),
.A2(n_3129),
.B1(n_3132),
.B2(n_3122),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3195),
.B(n_3002),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3276),
.Y(n_3329)
);

BUFx6f_ASAP7_75t_L g3330 ( 
.A(n_3183),
.Y(n_3330)
);

AOI22xp5_ASAP7_75t_L g3331 ( 
.A1(n_3211),
.A2(n_3002),
.B1(n_3008),
.B2(n_2985),
.Y(n_3331)
);

AND2x4_ASAP7_75t_L g3332 ( 
.A(n_3148),
.B(n_3028),
.Y(n_3332)
);

AO22x2_ASAP7_75t_L g3333 ( 
.A1(n_3262),
.A2(n_3139),
.B1(n_3137),
.B2(n_3102),
.Y(n_3333)
);

OAI221xp5_ASAP7_75t_L g3334 ( 
.A1(n_3223),
.A2(n_3106),
.B1(n_2993),
.B2(n_3000),
.C(n_2915),
.Y(n_3334)
);

AO22x2_ASAP7_75t_L g3335 ( 
.A1(n_3269),
.A2(n_3095),
.B1(n_3058),
.B2(n_3059),
.Y(n_3335)
);

INVxp67_ASAP7_75t_L g3336 ( 
.A(n_3187),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3279),
.Y(n_3337)
);

INVxp67_ASAP7_75t_L g3338 ( 
.A(n_3202),
.Y(n_3338)
);

BUFx3_ASAP7_75t_L g3339 ( 
.A(n_3157),
.Y(n_3339)
);

INVxp67_ASAP7_75t_SL g3340 ( 
.A(n_3271),
.Y(n_3340)
);

AOI22xp5_ASAP7_75t_L g3341 ( 
.A1(n_3149),
.A2(n_3083),
.B1(n_3020),
.B2(n_3024),
.Y(n_3341)
);

AOI22xp5_ASAP7_75t_L g3342 ( 
.A1(n_3193),
.A2(n_3020),
.B1(n_3019),
.B2(n_3098),
.Y(n_3342)
);

AO22x2_ASAP7_75t_L g3343 ( 
.A1(n_3285),
.A2(n_3061),
.B1(n_3062),
.B2(n_3054),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3161),
.B(n_3078),
.Y(n_3344)
);

INVxp67_ASAP7_75t_L g3345 ( 
.A(n_3210),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3234),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3235),
.Y(n_3347)
);

OAI221xp5_ASAP7_75t_L g3348 ( 
.A1(n_3283),
.A2(n_3138),
.B1(n_3104),
.B2(n_3107),
.C(n_2990),
.Y(n_3348)
);

AO22x2_ASAP7_75t_L g3349 ( 
.A1(n_3290),
.A2(n_3075),
.B1(n_3084),
.B2(n_3074),
.Y(n_3349)
);

CKINVDCx16_ASAP7_75t_R g3350 ( 
.A(n_3188),
.Y(n_3350)
);

BUFx2_ASAP7_75t_L g3351 ( 
.A(n_3169),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3237),
.Y(n_3352)
);

HB1xp67_ASAP7_75t_L g3353 ( 
.A(n_3267),
.Y(n_3353)
);

AND2x4_ASAP7_75t_L g3354 ( 
.A(n_3183),
.B(n_3090),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3162),
.B(n_2974),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3207),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3208),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_3217),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3231),
.B(n_2977),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3241),
.B(n_2979),
.Y(n_3360)
);

AO22x2_ASAP7_75t_L g3361 ( 
.A1(n_3220),
.A2(n_3092),
.B1(n_2981),
.B2(n_2984),
.Y(n_3361)
);

AND2x2_ASAP7_75t_L g3362 ( 
.A(n_3178),
.B(n_2847),
.Y(n_3362)
);

NOR2xp33_ASAP7_75t_L g3363 ( 
.A(n_3184),
.B(n_3125),
.Y(n_3363)
);

INVxp67_ASAP7_75t_L g3364 ( 
.A(n_3190),
.Y(n_3364)
);

NAND2x1p5_ASAP7_75t_L g3365 ( 
.A(n_3291),
.B(n_2819),
.Y(n_3365)
);

AO22x2_ASAP7_75t_L g3366 ( 
.A1(n_3280),
.A2(n_2987),
.B1(n_2994),
.B2(n_2983),
.Y(n_3366)
);

OAI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_3159),
.A2(n_3086),
.B1(n_3103),
.B2(n_3043),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3151),
.Y(n_3368)
);

AO22x2_ASAP7_75t_L g3369 ( 
.A1(n_3175),
.A2(n_2998),
.B1(n_2996),
.B2(n_3109),
.Y(n_3369)
);

AOI22xp5_ASAP7_75t_L g3370 ( 
.A1(n_3229),
.A2(n_3037),
.B1(n_3085),
.B2(n_3080),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3246),
.B(n_3087),
.Y(n_3371)
);

AO22x2_ASAP7_75t_L g3372 ( 
.A1(n_3189),
.A2(n_3073),
.B1(n_3134),
.B2(n_1902),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3155),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3176),
.B(n_2945),
.Y(n_3374)
);

HB1xp67_ASAP7_75t_L g3375 ( 
.A(n_3221),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3158),
.Y(n_3376)
);

NAND2x1p5_ASAP7_75t_L g3377 ( 
.A(n_3221),
.B(n_2819),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3166),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_3167),
.Y(n_3379)
);

NAND3xp33_ASAP7_75t_L g3380 ( 
.A(n_3226),
.B(n_1525),
.C(n_1522),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3173),
.Y(n_3381)
);

AO22x2_ASAP7_75t_L g3382 ( 
.A1(n_3200),
.A2(n_1910),
.B1(n_1926),
.B2(n_1918),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_3204),
.Y(n_3383)
);

AND2x4_ASAP7_75t_L g3384 ( 
.A(n_3232),
.B(n_2820),
.Y(n_3384)
);

INVx2_ASAP7_75t_L g3385 ( 
.A(n_3176),
.Y(n_3385)
);

NAND2x1p5_ASAP7_75t_L g3386 ( 
.A(n_3232),
.B(n_2820),
.Y(n_3386)
);

AOI22xp5_ASAP7_75t_L g3387 ( 
.A1(n_3230),
.A2(n_1537),
.B1(n_1538),
.B2(n_1527),
.Y(n_3387)
);

OAI22xp5_ASAP7_75t_L g3388 ( 
.A1(n_3140),
.A2(n_1540),
.B1(n_1541),
.B2(n_1539),
.Y(n_3388)
);

NOR2xp33_ASAP7_75t_L g3389 ( 
.A(n_3281),
.B(n_2842),
.Y(n_3389)
);

NAND2x1p5_ASAP7_75t_L g3390 ( 
.A(n_3248),
.B(n_2842),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_3176),
.Y(n_3391)
);

AO22x2_ASAP7_75t_L g3392 ( 
.A1(n_3170),
.A2(n_1927),
.B1(n_1943),
.B2(n_1929),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3252),
.Y(n_3393)
);

A2O1A1Ixp33_ASAP7_75t_L g3394 ( 
.A1(n_3147),
.A2(n_1958),
.B(n_1971),
.C(n_1963),
.Y(n_3394)
);

AOI22x1_ASAP7_75t_L g3395 ( 
.A1(n_3260),
.A2(n_1982),
.B1(n_1991),
.B2(n_1979),
.Y(n_3395)
);

NAND2x1p5_ASAP7_75t_L g3396 ( 
.A(n_3165),
.B(n_2848),
.Y(n_3396)
);

NAND2x1p5_ASAP7_75t_L g3397 ( 
.A(n_3255),
.B(n_3142),
.Y(n_3397)
);

NOR2xp67_ASAP7_75t_L g3398 ( 
.A(n_3191),
.B(n_2883),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3264),
.Y(n_3399)
);

AO22x2_ASAP7_75t_L g3400 ( 
.A1(n_3205),
.A2(n_3212),
.B1(n_3153),
.B2(n_3154),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3266),
.Y(n_3401)
);

BUFx8_ASAP7_75t_L g3402 ( 
.A(n_3156),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3287),
.Y(n_3403)
);

INVx2_ASAP7_75t_SL g3404 ( 
.A(n_3277),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3293),
.Y(n_3405)
);

OR2x2_ASAP7_75t_L g3406 ( 
.A(n_3199),
.B(n_2830),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_3176),
.Y(n_3407)
);

NOR2xp33_ASAP7_75t_L g3408 ( 
.A(n_3192),
.B(n_3272),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_SL g3409 ( 
.A(n_3145),
.B(n_2848),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3273),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_3292),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3274),
.Y(n_3412)
);

AO22x2_ASAP7_75t_L g3413 ( 
.A1(n_3227),
.A2(n_2003),
.B1(n_2013),
.B2(n_2012),
.Y(n_3413)
);

AOI22x1_ASAP7_75t_L g3414 ( 
.A1(n_3146),
.A2(n_2022),
.B1(n_2034),
.B2(n_2021),
.Y(n_3414)
);

NAND2x1p5_ASAP7_75t_L g3415 ( 
.A(n_3238),
.B(n_2859),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3216),
.Y(n_3416)
);

AO22x2_ASAP7_75t_L g3417 ( 
.A1(n_3263),
.A2(n_2039),
.B1(n_2040),
.B2(n_2035),
.Y(n_3417)
);

BUFx6f_ASAP7_75t_SL g3418 ( 
.A(n_3275),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3218),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3292),
.Y(n_3420)
);

INVx1_ASAP7_75t_SL g3421 ( 
.A(n_3258),
.Y(n_3421)
);

NAND2x1p5_ASAP7_75t_L g3422 ( 
.A(n_3177),
.B(n_2859),
.Y(n_3422)
);

AO22x2_ASAP7_75t_L g3423 ( 
.A1(n_3219),
.A2(n_2053),
.B1(n_2054),
.B2(n_2047),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3222),
.B(n_1542),
.Y(n_3424)
);

AO22x2_ASAP7_75t_L g3425 ( 
.A1(n_3249),
.A2(n_2066),
.B1(n_2070),
.B2(n_2056),
.Y(n_3425)
);

NAND3xp33_ASAP7_75t_L g3426 ( 
.A(n_3303),
.B(n_3395),
.C(n_3301),
.Y(n_3426)
);

AOI22xp5_ASAP7_75t_L g3427 ( 
.A1(n_3311),
.A2(n_3288),
.B1(n_3206),
.B2(n_3256),
.Y(n_3427)
);

NOR2x1_ASAP7_75t_SL g3428 ( 
.A(n_3385),
.B(n_3163),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_SL g3429 ( 
.A(n_3363),
.B(n_3292),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3410),
.B(n_3250),
.Y(n_3430)
);

BUFx4f_ASAP7_75t_L g3431 ( 
.A(n_3305),
.Y(n_3431)
);

O2A1O1Ixp5_ASAP7_75t_L g3432 ( 
.A1(n_3409),
.A2(n_3367),
.B(n_3394),
.C(n_3310),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3412),
.B(n_3213),
.Y(n_3433)
);

OAI22xp5_ASAP7_75t_L g3434 ( 
.A1(n_3302),
.A2(n_3289),
.B1(n_3261),
.B2(n_3164),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3416),
.B(n_3294),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3419),
.B(n_3278),
.Y(n_3436)
);

BUFx3_ASAP7_75t_L g3437 ( 
.A(n_3307),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3364),
.B(n_3282),
.Y(n_3438)
);

AOI21xp5_ASAP7_75t_L g3439 ( 
.A1(n_3391),
.A2(n_3236),
.B(n_3201),
.Y(n_3439)
);

AOI21xp5_ASAP7_75t_L g3440 ( 
.A1(n_3407),
.A2(n_3420),
.B(n_3411),
.Y(n_3440)
);

OAI22xp5_ASAP7_75t_L g3441 ( 
.A1(n_3321),
.A2(n_3295),
.B1(n_3233),
.B2(n_3179),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_SL g3442 ( 
.A(n_3328),
.B(n_3292),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3340),
.B(n_3247),
.Y(n_3443)
);

AOI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_3400),
.A2(n_3270),
.B(n_3168),
.Y(n_3444)
);

OAI22xp5_ASAP7_75t_L g3445 ( 
.A1(n_3380),
.A2(n_3185),
.B1(n_3196),
.B2(n_3186),
.Y(n_3445)
);

AOI21xp5_ASAP7_75t_L g3446 ( 
.A1(n_3371),
.A2(n_3242),
.B(n_3240),
.Y(n_3446)
);

AOI21xp5_ASAP7_75t_L g3447 ( 
.A1(n_3370),
.A2(n_3245),
.B(n_3286),
.Y(n_3447)
);

AO22x1_ASAP7_75t_L g3448 ( 
.A1(n_3402),
.A2(n_3181),
.B1(n_1546),
.B2(n_1548),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3393),
.B(n_3254),
.Y(n_3449)
);

NOR2xp33_ASAP7_75t_L g3450 ( 
.A(n_3338),
.B(n_3257),
.Y(n_3450)
);

BUFx6f_ASAP7_75t_L g3451 ( 
.A(n_3330),
.Y(n_3451)
);

AOI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_3348),
.A2(n_3284),
.B(n_2781),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3296),
.Y(n_3453)
);

NAND2xp33_ASAP7_75t_L g3454 ( 
.A(n_3414),
.B(n_3308),
.Y(n_3454)
);

NAND3xp33_ASAP7_75t_L g3455 ( 
.A(n_3387),
.B(n_1550),
.C(n_1545),
.Y(n_3455)
);

AOI22xp5_ASAP7_75t_L g3456 ( 
.A1(n_3408),
.A2(n_1558),
.B1(n_1563),
.B2(n_1557),
.Y(n_3456)
);

NOR2xp33_ASAP7_75t_L g3457 ( 
.A(n_3322),
.B(n_2866),
.Y(n_3457)
);

OAI22xp5_ASAP7_75t_L g3458 ( 
.A1(n_3424),
.A2(n_1572),
.B1(n_1578),
.B2(n_1565),
.Y(n_3458)
);

NOR2xp67_ASAP7_75t_SL g3459 ( 
.A(n_3339),
.B(n_2866),
.Y(n_3459)
);

BUFx3_ASAP7_75t_L g3460 ( 
.A(n_3330),
.Y(n_3460)
);

AOI21xp5_ASAP7_75t_L g3461 ( 
.A1(n_3355),
.A2(n_3401),
.B(n_3399),
.Y(n_3461)
);

AOI21xp5_ASAP7_75t_L g3462 ( 
.A1(n_3403),
.A2(n_1877),
.B(n_1609),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3304),
.Y(n_3463)
);

OAI21xp33_ASAP7_75t_L g3464 ( 
.A1(n_3388),
.A2(n_1580),
.B(n_1579),
.Y(n_3464)
);

OAI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_3405),
.A2(n_3005),
.B(n_2931),
.Y(n_3465)
);

O2A1O1Ixp33_ASAP7_75t_L g3466 ( 
.A1(n_3353),
.A2(n_2075),
.B(n_2081),
.C(n_2071),
.Y(n_3466)
);

AOI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_3297),
.A2(n_1877),
.B(n_1609),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3298),
.B(n_1581),
.Y(n_3468)
);

AOI21xp5_ASAP7_75t_L g3469 ( 
.A1(n_3299),
.A2(n_1877),
.B(n_1609),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3336),
.B(n_1582),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3300),
.Y(n_3471)
);

AOI22xp33_ASAP7_75t_SL g3472 ( 
.A1(n_3317),
.A2(n_2093),
.B1(n_1585),
.B2(n_1587),
.Y(n_3472)
);

AND2x4_ASAP7_75t_L g3473 ( 
.A(n_3314),
.B(n_2880),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_3309),
.A2(n_1993),
.B(n_1920),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_3360),
.B(n_1586),
.Y(n_3475)
);

AO22x1_ASAP7_75t_L g3476 ( 
.A1(n_3325),
.A2(n_3362),
.B1(n_3345),
.B2(n_3332),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3318),
.B(n_1588),
.Y(n_3477)
);

AOI21xp5_ASAP7_75t_L g3478 ( 
.A1(n_3324),
.A2(n_1993),
.B(n_1920),
.Y(n_3478)
);

OAI21xp33_ASAP7_75t_L g3479 ( 
.A1(n_3413),
.A2(n_1598),
.B(n_1594),
.Y(n_3479)
);

OAI21xp5_ASAP7_75t_L g3480 ( 
.A1(n_3359),
.A2(n_2019),
.B(n_1875),
.Y(n_3480)
);

NAND3xp33_ASAP7_75t_L g3481 ( 
.A(n_3334),
.B(n_1600),
.C(n_1599),
.Y(n_3481)
);

AOI21xp5_ASAP7_75t_L g3482 ( 
.A1(n_3329),
.A2(n_1993),
.B(n_1920),
.Y(n_3482)
);

NOR2xp33_ASAP7_75t_L g3483 ( 
.A(n_3350),
.B(n_2880),
.Y(n_3483)
);

A2O1A1Ixp33_ASAP7_75t_L g3484 ( 
.A1(n_3374),
.A2(n_2001),
.B(n_2005),
.C(n_1957),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3351),
.B(n_1605),
.Y(n_3485)
);

O2A1O1Ixp5_ASAP7_75t_L g3486 ( 
.A1(n_3344),
.A2(n_2080),
.B(n_2024),
.C(n_1802),
.Y(n_3486)
);

AOI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_3369),
.A2(n_1483),
.B(n_1482),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_3315),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3337),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_3421),
.B(n_1607),
.Y(n_3490)
);

AO32x1_ASAP7_75t_L g3491 ( 
.A1(n_3346),
.A2(n_3),
.A3(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3397),
.B(n_3306),
.Y(n_3492)
);

BUFx6f_ASAP7_75t_L g3493 ( 
.A(n_3354),
.Y(n_3493)
);

A2O1A1Ixp33_ASAP7_75t_L g3494 ( 
.A1(n_3342),
.A2(n_1615),
.B(n_1617),
.C(n_1613),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3331),
.B(n_1619),
.Y(n_3495)
);

AOI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_3312),
.A2(n_1518),
.B(n_1490),
.Y(n_3496)
);

OAI22xp5_ASAP7_75t_L g3497 ( 
.A1(n_3341),
.A2(n_1628),
.B1(n_1630),
.B2(n_1624),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_SL g3498 ( 
.A(n_3390),
.B(n_2501),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3323),
.Y(n_3499)
);

BUFx6f_ASAP7_75t_L g3500 ( 
.A(n_3365),
.Y(n_3500)
);

AOI21xp5_ASAP7_75t_L g3501 ( 
.A1(n_3313),
.A2(n_1526),
.B(n_1519),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3375),
.B(n_1633),
.Y(n_3502)
);

AOI21xp5_ASAP7_75t_L g3503 ( 
.A1(n_3343),
.A2(n_1536),
.B(n_1534),
.Y(n_3503)
);

AOI21xp5_ASAP7_75t_L g3504 ( 
.A1(n_3335),
.A2(n_1552),
.B(n_1547),
.Y(n_3504)
);

INVx2_ASAP7_75t_L g3505 ( 
.A(n_3358),
.Y(n_3505)
);

AOI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_3361),
.A2(n_1576),
.B(n_1575),
.Y(n_3506)
);

AND2x4_ASAP7_75t_L g3507 ( 
.A(n_3384),
.B(n_2504),
.Y(n_3507)
);

NAND2x1p5_ASAP7_75t_L g3508 ( 
.A(n_3326),
.B(n_2508),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_3319),
.A2(n_1596),
.B(n_1589),
.Y(n_3509)
);

O2A1O1Ixp5_ASAP7_75t_L g3510 ( 
.A1(n_3389),
.A2(n_1802),
.B(n_1458),
.C(n_1642),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3379),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3347),
.Y(n_3512)
);

AOI21xp5_ASAP7_75t_L g3513 ( 
.A1(n_3327),
.A2(n_1612),
.B(n_1610),
.Y(n_3513)
);

NOR2xp33_ASAP7_75t_L g3514 ( 
.A(n_3320),
.B(n_3404),
.Y(n_3514)
);

AOI21xp5_ASAP7_75t_L g3515 ( 
.A1(n_3333),
.A2(n_1618),
.B(n_1614),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_3382),
.B(n_3316),
.Y(n_3516)
);

AOI21xp5_ASAP7_75t_L g3517 ( 
.A1(n_3349),
.A2(n_1623),
.B(n_1620),
.Y(n_3517)
);

BUFx4f_ASAP7_75t_L g3518 ( 
.A(n_3377),
.Y(n_3518)
);

OAI22xp5_ASAP7_75t_L g3519 ( 
.A1(n_3398),
.A2(n_1641),
.B1(n_1646),
.B2(n_1645),
.Y(n_3519)
);

NOR2xp33_ASAP7_75t_L g3520 ( 
.A(n_3406),
.B(n_3386),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3383),
.Y(n_3521)
);

AOI22xp5_ASAP7_75t_L g3522 ( 
.A1(n_3417),
.A2(n_1650),
.B1(n_1653),
.B2(n_1647),
.Y(n_3522)
);

INVx2_ASAP7_75t_SL g3523 ( 
.A(n_3396),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_3352),
.B(n_1655),
.Y(n_3524)
);

OR2x2_ASAP7_75t_L g3525 ( 
.A(n_3356),
.B(n_2519),
.Y(n_3525)
);

AND2x2_ASAP7_75t_SL g3526 ( 
.A(n_3357),
.B(n_2521),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3368),
.B(n_1657),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3373),
.B(n_1659),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3376),
.B(n_1666),
.Y(n_3529)
);

NOR2xp33_ASAP7_75t_SL g3530 ( 
.A(n_3418),
.B(n_1625),
.Y(n_3530)
);

NOR2xp33_ASAP7_75t_L g3531 ( 
.A(n_3422),
.B(n_1672),
.Y(n_3531)
);

NOR2xp33_ASAP7_75t_L g3532 ( 
.A(n_3415),
.B(n_1674),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3378),
.B(n_3381),
.Y(n_3533)
);

NOR2xp67_ASAP7_75t_SL g3534 ( 
.A(n_3426),
.B(n_3438),
.Y(n_3534)
);

O2A1O1Ixp33_ASAP7_75t_L g3535 ( 
.A1(n_3434),
.A2(n_3441),
.B(n_3494),
.C(n_3435),
.Y(n_3535)
);

BUFx3_ASAP7_75t_L g3536 ( 
.A(n_3460),
.Y(n_3536)
);

INVx2_ASAP7_75t_SL g3537 ( 
.A(n_3431),
.Y(n_3537)
);

BUFx6f_ASAP7_75t_L g3538 ( 
.A(n_3518),
.Y(n_3538)
);

INVx3_ASAP7_75t_L g3539 ( 
.A(n_3451),
.Y(n_3539)
);

AOI21xp5_ASAP7_75t_L g3540 ( 
.A1(n_3429),
.A2(n_3366),
.B(n_3372),
.Y(n_3540)
);

AOI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_3446),
.A2(n_3392),
.B(n_3425),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3430),
.B(n_3423),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_3463),
.Y(n_3543)
);

AND2x4_ASAP7_75t_L g3544 ( 
.A(n_3437),
.B(n_2528),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3489),
.Y(n_3545)
);

BUFx2_ASAP7_75t_L g3546 ( 
.A(n_3451),
.Y(n_3546)
);

O2A1O1Ixp33_ASAP7_75t_L g3547 ( 
.A1(n_3466),
.A2(n_1678),
.B(n_1679),
.C(n_1677),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3453),
.Y(n_3548)
);

O2A1O1Ixp33_ASAP7_75t_L g3549 ( 
.A1(n_3458),
.A2(n_1684),
.B(n_1692),
.C(n_1683),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_SL g3550 ( 
.A(n_3427),
.B(n_3443),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3488),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3471),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3433),
.B(n_1697),
.Y(n_3553)
);

INVx3_ASAP7_75t_L g3554 ( 
.A(n_3493),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3512),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3436),
.B(n_1700),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3461),
.B(n_1703),
.Y(n_3557)
);

INVx2_ASAP7_75t_L g3558 ( 
.A(n_3499),
.Y(n_3558)
);

AOI22xp33_ASAP7_75t_L g3559 ( 
.A1(n_3479),
.A2(n_1704),
.B1(n_1712),
.B2(n_1705),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3505),
.Y(n_3560)
);

NAND2x1p5_ASAP7_75t_L g3561 ( 
.A(n_3459),
.B(n_2532),
.Y(n_3561)
);

O2A1O1Ixp33_ASAP7_75t_SL g3562 ( 
.A1(n_3514),
.A2(n_5),
.B(n_0),
.C(n_3),
.Y(n_3562)
);

INVx2_ASAP7_75t_L g3563 ( 
.A(n_3511),
.Y(n_3563)
);

INVx2_ASAP7_75t_SL g3564 ( 
.A(n_3493),
.Y(n_3564)
);

NOR2xp33_ASAP7_75t_L g3565 ( 
.A(n_3530),
.B(n_1714),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3533),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3520),
.B(n_1715),
.Y(n_3567)
);

INVx1_ASAP7_75t_SL g3568 ( 
.A(n_3473),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3521),
.Y(n_3569)
);

INVx2_ASAP7_75t_SL g3570 ( 
.A(n_3500),
.Y(n_3570)
);

INVx2_ASAP7_75t_L g3571 ( 
.A(n_3525),
.Y(n_3571)
);

BUFx4_ASAP7_75t_SL g3572 ( 
.A(n_3481),
.Y(n_3572)
);

BUFx6f_ASAP7_75t_L g3573 ( 
.A(n_3500),
.Y(n_3573)
);

BUFx2_ASAP7_75t_L g3574 ( 
.A(n_3492),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3526),
.B(n_1716),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3449),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3516),
.Y(n_3577)
);

O2A1O1Ixp33_ASAP7_75t_L g3578 ( 
.A1(n_3497),
.A2(n_1723),
.B(n_1725),
.C(n_1717),
.Y(n_3578)
);

AOI22xp33_ASAP7_75t_L g3579 ( 
.A1(n_3472),
.A2(n_1727),
.B1(n_1737),
.B2(n_1732),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3442),
.Y(n_3580)
);

OAI22xp5_ASAP7_75t_L g3581 ( 
.A1(n_3455),
.A2(n_1742),
.B1(n_1743),
.B2(n_1738),
.Y(n_3581)
);

CKINVDCx16_ASAP7_75t_R g3582 ( 
.A(n_3483),
.Y(n_3582)
);

AND2x2_ASAP7_75t_L g3583 ( 
.A(n_3468),
.B(n_1748),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3465),
.Y(n_3584)
);

BUFx6f_ASAP7_75t_L g3585 ( 
.A(n_3507),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_3523),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_SL g3587 ( 
.A(n_3432),
.B(n_2538),
.Y(n_3587)
);

NOR2xp33_ASAP7_75t_L g3588 ( 
.A(n_3450),
.B(n_1752),
.Y(n_3588)
);

A2O1A1Ixp33_ASAP7_75t_L g3589 ( 
.A1(n_3447),
.A2(n_3496),
.B(n_3480),
.C(n_3484),
.Y(n_3589)
);

BUFx6f_ASAP7_75t_L g3590 ( 
.A(n_3508),
.Y(n_3590)
);

INVx1_ASAP7_75t_SL g3591 ( 
.A(n_3476),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3428),
.Y(n_3592)
);

NOR2xp33_ASAP7_75t_L g3593 ( 
.A(n_3457),
.B(n_1757),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3475),
.B(n_1761),
.Y(n_3594)
);

NOR3xp33_ASAP7_75t_SL g3595 ( 
.A(n_3464),
.B(n_1772),
.C(n_1766),
.Y(n_3595)
);

A2O1A1Ixp33_ASAP7_75t_L g3596 ( 
.A1(n_3504),
.A2(n_1778),
.B(n_1779),
.C(n_1773),
.Y(n_3596)
);

INVx2_ASAP7_75t_L g3597 ( 
.A(n_3527),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3528),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3439),
.A2(n_1651),
.B(n_1648),
.Y(n_3599)
);

OAI22xp5_ASAP7_75t_L g3600 ( 
.A1(n_3456),
.A2(n_1782),
.B1(n_1787),
.B2(n_1780),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3529),
.Y(n_3601)
);

A2O1A1Ixp33_ASAP7_75t_L g3602 ( 
.A1(n_3515),
.A2(n_1790),
.B(n_1793),
.C(n_1788),
.Y(n_3602)
);

AOI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_3444),
.A2(n_1658),
.B(n_1652),
.Y(n_3603)
);

NOR2xp33_ASAP7_75t_L g3604 ( 
.A(n_3532),
.B(n_1794),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3440),
.Y(n_3605)
);

AOI21xp5_ASAP7_75t_L g3606 ( 
.A1(n_3454),
.A2(n_1662),
.B(n_1661),
.Y(n_3606)
);

INVx2_ASAP7_75t_L g3607 ( 
.A(n_3486),
.Y(n_3607)
);

BUFx6f_ASAP7_75t_L g3608 ( 
.A(n_3498),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3477),
.Y(n_3609)
);

O2A1O1Ixp33_ASAP7_75t_L g3610 ( 
.A1(n_3519),
.A2(n_3495),
.B(n_3485),
.C(n_3470),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_3524),
.Y(n_3611)
);

AOI21xp5_ASAP7_75t_L g3612 ( 
.A1(n_3452),
.A2(n_1664),
.B(n_1663),
.Y(n_3612)
);

BUFx2_ASAP7_75t_L g3613 ( 
.A(n_3502),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3491),
.Y(n_3614)
);

OAI21xp33_ASAP7_75t_L g3615 ( 
.A1(n_3522),
.A2(n_1797),
.B(n_1796),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_SL g3616 ( 
.A(n_3445),
.B(n_2568),
.Y(n_3616)
);

CKINVDCx5p33_ASAP7_75t_R g3617 ( 
.A(n_3490),
.Y(n_3617)
);

A2O1A1Ixp33_ASAP7_75t_L g3618 ( 
.A1(n_3517),
.A2(n_1808),
.B(n_1812),
.C(n_1807),
.Y(n_3618)
);

NOR3xp33_ASAP7_75t_SL g3619 ( 
.A(n_3531),
.B(n_1818),
.C(n_1813),
.Y(n_3619)
);

INVx3_ASAP7_75t_L g3620 ( 
.A(n_3448),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_SL g3621 ( 
.A(n_3503),
.B(n_2581),
.Y(n_3621)
);

OAI22xp5_ASAP7_75t_L g3622 ( 
.A1(n_3501),
.A2(n_1827),
.B1(n_1830),
.B2(n_1820),
.Y(n_3622)
);

NOR2xp33_ASAP7_75t_L g3623 ( 
.A(n_3509),
.B(n_1835),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3513),
.B(n_1841),
.Y(n_3624)
);

OAI21x1_ASAP7_75t_L g3625 ( 
.A1(n_3462),
.A2(n_1802),
.B(n_1458),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_3510),
.A2(n_3469),
.B(n_3467),
.Y(n_3626)
);

A2O1A1Ixp33_ASAP7_75t_L g3627 ( 
.A1(n_3487),
.A2(n_1850),
.B(n_1851),
.C(n_1844),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3506),
.B(n_1852),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_3491),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_3474),
.Y(n_3630)
);

AOI22xp5_ASAP7_75t_L g3631 ( 
.A1(n_3478),
.A2(n_1857),
.B1(n_1861),
.B2(n_1855),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3482),
.B(n_1863),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3430),
.B(n_1866),
.Y(n_3633)
);

CKINVDCx20_ASAP7_75t_R g3634 ( 
.A(n_3431),
.Y(n_3634)
);

NOR2xp33_ASAP7_75t_L g3635 ( 
.A(n_3427),
.B(n_1867),
.Y(n_3635)
);

NOR2xp33_ASAP7_75t_L g3636 ( 
.A(n_3427),
.B(n_1868),
.Y(n_3636)
);

O2A1O1Ixp5_ASAP7_75t_SL g3637 ( 
.A1(n_3429),
.A2(n_1802),
.B(n_1458),
.C(n_1870),
.Y(n_3637)
);

AOI22xp5_ASAP7_75t_L g3638 ( 
.A1(n_3427),
.A2(n_1873),
.B1(n_1879),
.B2(n_1872),
.Y(n_3638)
);

NOR3xp33_ASAP7_75t_L g3639 ( 
.A(n_3426),
.B(n_1883),
.C(n_1881),
.Y(n_3639)
);

OAI22xp33_ASAP7_75t_L g3640 ( 
.A1(n_3427),
.A2(n_1887),
.B1(n_1890),
.B2(n_1884),
.Y(n_3640)
);

O2A1O1Ixp33_ASAP7_75t_L g3641 ( 
.A1(n_3434),
.A2(n_1899),
.B(n_1901),
.C(n_1896),
.Y(n_3641)
);

AND2x4_ASAP7_75t_L g3642 ( 
.A(n_3437),
.B(n_2309),
.Y(n_3642)
);

NOR3xp33_ASAP7_75t_SL g3643 ( 
.A(n_3455),
.B(n_1908),
.C(n_1904),
.Y(n_3643)
);

NOR2xp33_ASAP7_75t_L g3644 ( 
.A(n_3427),
.B(n_1911),
.Y(n_3644)
);

NOR2xp33_ASAP7_75t_L g3645 ( 
.A(n_3427),
.B(n_1914),
.Y(n_3645)
);

AO31x2_ASAP7_75t_L g3646 ( 
.A1(n_3589),
.A2(n_1802),
.A3(n_1458),
.B(n_1671),
.Y(n_3646)
);

NOR4xp25_ASAP7_75t_L g3647 ( 
.A(n_3535),
.B(n_9),
.C(n_6),
.D(n_8),
.Y(n_3647)
);

AOI22xp33_ASAP7_75t_L g3648 ( 
.A1(n_3635),
.A2(n_1916),
.B1(n_1922),
.B2(n_1921),
.Y(n_3648)
);

OAI21x1_ASAP7_75t_SL g3649 ( 
.A1(n_3641),
.A2(n_8),
.B(n_9),
.Y(n_3649)
);

OAI21x1_ASAP7_75t_L g3650 ( 
.A1(n_3625),
.A2(n_1458),
.B(n_1048),
.Y(n_3650)
);

OAI21xp5_ASAP7_75t_L g3651 ( 
.A1(n_3645),
.A2(n_1945),
.B(n_1924),
.Y(n_3651)
);

OAI21x1_ASAP7_75t_L g3652 ( 
.A1(n_3626),
.A2(n_1051),
.B(n_1046),
.Y(n_3652)
);

BUFx10_ASAP7_75t_L g3653 ( 
.A(n_3538),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3550),
.B(n_1923),
.Y(n_3654)
);

BUFx3_ASAP7_75t_L g3655 ( 
.A(n_3536),
.Y(n_3655)
);

AOI221x1_ASAP7_75t_L g3656 ( 
.A1(n_3636),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.C(n_14),
.Y(n_3656)
);

OAI21x1_ASAP7_75t_L g3657 ( 
.A1(n_3630),
.A2(n_1053),
.B(n_1052),
.Y(n_3657)
);

AOI221x1_ASAP7_75t_L g3658 ( 
.A1(n_3644),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.C(n_14),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3576),
.B(n_1930),
.Y(n_3659)
);

OAI21x1_ASAP7_75t_SL g3660 ( 
.A1(n_3541),
.A2(n_15),
.B(n_16),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3566),
.B(n_1932),
.Y(n_3661)
);

AOI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3587),
.A2(n_2092),
.B(n_2091),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3534),
.B(n_1934),
.Y(n_3663)
);

A2O1A1Ixp33_ASAP7_75t_L g3664 ( 
.A1(n_3604),
.A2(n_1944),
.B(n_1948),
.C(n_1946),
.Y(n_3664)
);

NAND3xp33_ASAP7_75t_L g3665 ( 
.A(n_3588),
.B(n_3639),
.C(n_3638),
.Y(n_3665)
);

AO31x2_ASAP7_75t_L g3666 ( 
.A1(n_3540),
.A2(n_1673),
.A3(n_1676),
.B(n_1667),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3542),
.B(n_1936),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3548),
.B(n_1951),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3552),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3555),
.B(n_1953),
.Y(n_3670)
);

OAI21xp5_ASAP7_75t_L g3671 ( 
.A1(n_3603),
.A2(n_3640),
.B(n_3565),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3577),
.B(n_15),
.Y(n_3672)
);

INVxp67_ASAP7_75t_L g3673 ( 
.A(n_3613),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3545),
.Y(n_3674)
);

OAI21xp5_ASAP7_75t_L g3675 ( 
.A1(n_3616),
.A2(n_1975),
.B(n_1961),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3574),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3609),
.B(n_1956),
.Y(n_3677)
);

OAI21x1_ASAP7_75t_L g3678 ( 
.A1(n_3607),
.A2(n_1056),
.B(n_1054),
.Y(n_3678)
);

INVxp67_ASAP7_75t_SL g3679 ( 
.A(n_3605),
.Y(n_3679)
);

OAI21x1_ASAP7_75t_SL g3680 ( 
.A1(n_3610),
.A2(n_16),
.B(n_17),
.Y(n_3680)
);

AO31x2_ASAP7_75t_L g3681 ( 
.A1(n_3629),
.A2(n_1687),
.A3(n_1690),
.B(n_1686),
.Y(n_3681)
);

INVx4_ASAP7_75t_L g3682 ( 
.A(n_3538),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3611),
.B(n_1962),
.Y(n_3683)
);

OAI21xp5_ASAP7_75t_L g3684 ( 
.A1(n_3623),
.A2(n_2032),
.B(n_1981),
.Y(n_3684)
);

AO21x2_ASAP7_75t_L g3685 ( 
.A1(n_3599),
.A2(n_2082),
.B(n_2073),
.Y(n_3685)
);

OAI21x1_ASAP7_75t_L g3686 ( 
.A1(n_3637),
.A2(n_1059),
.B(n_1058),
.Y(n_3686)
);

AOI221x1_ASAP7_75t_L g3687 ( 
.A1(n_3557),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.C(n_20),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3543),
.Y(n_3688)
);

AOI221x1_ASAP7_75t_L g3689 ( 
.A1(n_3615),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.C(n_23),
.Y(n_3689)
);

OAI21x1_ASAP7_75t_L g3690 ( 
.A1(n_3584),
.A2(n_3592),
.B(n_3580),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_SL g3691 ( 
.A(n_3582),
.B(n_1693),
.Y(n_3691)
);

AOI21xp5_ASAP7_75t_L g3692 ( 
.A1(n_3612),
.A2(n_2094),
.B(n_1965),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3551),
.Y(n_3693)
);

AOI21x1_ASAP7_75t_SL g3694 ( 
.A1(n_3628),
.A2(n_21),
.B(n_22),
.Y(n_3694)
);

AOI21x1_ASAP7_75t_L g3695 ( 
.A1(n_3614),
.A2(n_1967),
.B(n_1964),
.Y(n_3695)
);

AND2x6_ASAP7_75t_L g3696 ( 
.A(n_3591),
.B(n_1063),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3597),
.B(n_1969),
.Y(n_3697)
);

OAI21x1_ASAP7_75t_L g3698 ( 
.A1(n_3621),
.A2(n_3560),
.B(n_3558),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3598),
.B(n_1972),
.Y(n_3699)
);

INVx3_ASAP7_75t_L g3700 ( 
.A(n_3573),
.Y(n_3700)
);

AO21x2_ASAP7_75t_L g3701 ( 
.A1(n_3632),
.A2(n_2090),
.B(n_2068),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3601),
.B(n_1973),
.Y(n_3702)
);

AOI21xp5_ASAP7_75t_L g3703 ( 
.A1(n_3562),
.A2(n_2079),
.B(n_2077),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3563),
.Y(n_3704)
);

OAI21x1_ASAP7_75t_L g3705 ( 
.A1(n_3569),
.A2(n_1066),
.B(n_1064),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3571),
.Y(n_3706)
);

OAI21x1_ASAP7_75t_L g3707 ( 
.A1(n_3631),
.A2(n_1069),
.B(n_1068),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3586),
.Y(n_3708)
);

AO21x2_ASAP7_75t_L g3709 ( 
.A1(n_3627),
.A2(n_2055),
.B(n_2043),
.Y(n_3709)
);

OAI21x1_ASAP7_75t_L g3710 ( 
.A1(n_3606),
.A2(n_1074),
.B(n_1073),
.Y(n_3710)
);

OAI21x1_ASAP7_75t_L g3711 ( 
.A1(n_3539),
.A2(n_1078),
.B(n_1076),
.Y(n_3711)
);

OAI22x1_ASAP7_75t_L g3712 ( 
.A1(n_3620),
.A2(n_1987),
.B1(n_1989),
.B2(n_1977),
.Y(n_3712)
);

AOI21xp5_ASAP7_75t_L g3713 ( 
.A1(n_3596),
.A2(n_2076),
.B(n_2067),
.Y(n_3713)
);

OAI21x1_ASAP7_75t_L g3714 ( 
.A1(n_3561),
.A2(n_1081),
.B(n_1080),
.Y(n_3714)
);

INVx2_ASAP7_75t_SL g3715 ( 
.A(n_3573),
.Y(n_3715)
);

OAI22xp5_ASAP7_75t_L g3716 ( 
.A1(n_3579),
.A2(n_2006),
.B1(n_2046),
.B2(n_1994),
.Y(n_3716)
);

OAI21x1_ASAP7_75t_L g3717 ( 
.A1(n_3624),
.A2(n_1087),
.B(n_1085),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3553),
.B(n_1983),
.Y(n_3718)
);

AOI21xp5_ASAP7_75t_L g3719 ( 
.A1(n_3602),
.A2(n_2045),
.B(n_2041),
.Y(n_3719)
);

O2A1O1Ixp33_ASAP7_75t_SL g3720 ( 
.A1(n_3578),
.A2(n_3618),
.B(n_3549),
.C(n_3547),
.Y(n_3720)
);

AO21x1_ASAP7_75t_L g3721 ( 
.A1(n_3593),
.A2(n_23),
.B(n_24),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3546),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3633),
.B(n_1992),
.Y(n_3723)
);

NOR3xp33_ASAP7_75t_SL g3724 ( 
.A(n_3622),
.B(n_1998),
.C(n_1997),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3570),
.Y(n_3725)
);

BUFx3_ASAP7_75t_L g3726 ( 
.A(n_3634),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3568),
.B(n_2000),
.Y(n_3727)
);

OAI21xp5_ASAP7_75t_L g3728 ( 
.A1(n_3595),
.A2(n_2033),
.B(n_2008),
.Y(n_3728)
);

OAI21x1_ASAP7_75t_L g3729 ( 
.A1(n_3554),
.A2(n_1091),
.B(n_1088),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3608),
.Y(n_3730)
);

OAI21x1_ASAP7_75t_L g3731 ( 
.A1(n_3559),
.A2(n_1094),
.B(n_1092),
.Y(n_3731)
);

OAI21x1_ASAP7_75t_L g3732 ( 
.A1(n_3567),
.A2(n_1097),
.B(n_1096),
.Y(n_3732)
);

AOI21xp5_ASAP7_75t_L g3733 ( 
.A1(n_3594),
.A2(n_2037),
.B(n_2031),
.Y(n_3733)
);

NAND2x1p5_ASAP7_75t_L g3734 ( 
.A(n_3537),
.B(n_3590),
.Y(n_3734)
);

AO32x2_ASAP7_75t_L g3735 ( 
.A1(n_3564),
.A2(n_26),
.A3(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3556),
.B(n_2004),
.Y(n_3736)
);

OAI21xp5_ASAP7_75t_L g3737 ( 
.A1(n_3600),
.A2(n_2023),
.B(n_2016),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3608),
.Y(n_3738)
);

OAI21x1_ASAP7_75t_L g3739 ( 
.A1(n_3575),
.A2(n_1101),
.B(n_1099),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3585),
.Y(n_3740)
);

AOI22xp5_ASAP7_75t_L g3741 ( 
.A1(n_3617),
.A2(n_2027),
.B1(n_2050),
.B2(n_2025),
.Y(n_3741)
);

AND2x2_ASAP7_75t_SL g3742 ( 
.A(n_3647),
.B(n_3590),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3669),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3674),
.Y(n_3744)
);

OAI21x1_ASAP7_75t_L g3745 ( 
.A1(n_3652),
.A2(n_3581),
.B(n_3572),
.Y(n_3745)
);

NOR2xp33_ASAP7_75t_L g3746 ( 
.A(n_3655),
.B(n_3583),
.Y(n_3746)
);

INVx2_ASAP7_75t_L g3747 ( 
.A(n_3704),
.Y(n_3747)
);

INVx3_ASAP7_75t_L g3748 ( 
.A(n_3700),
.Y(n_3748)
);

BUFx3_ASAP7_75t_L g3749 ( 
.A(n_3726),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3676),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3688),
.Y(n_3751)
);

OAI21x1_ASAP7_75t_L g3752 ( 
.A1(n_3650),
.A2(n_3643),
.B(n_3619),
.Y(n_3752)
);

OAI21x1_ASAP7_75t_L g3753 ( 
.A1(n_3690),
.A2(n_3544),
.B(n_3585),
.Y(n_3753)
);

OAI22xp5_ASAP7_75t_L g3754 ( 
.A1(n_3665),
.A2(n_2059),
.B1(n_2062),
.B2(n_2058),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3693),
.Y(n_3755)
);

NAND2x1p5_ASAP7_75t_L g3756 ( 
.A(n_3715),
.B(n_3642),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3706),
.Y(n_3757)
);

NAND3xp33_ASAP7_75t_L g3758 ( 
.A(n_3656),
.B(n_2086),
.C(n_2083),
.Y(n_3758)
);

NOR2xp33_ASAP7_75t_L g3759 ( 
.A(n_3682),
.B(n_25),
.Y(n_3759)
);

AOI21xp5_ASAP7_75t_L g3760 ( 
.A1(n_3679),
.A2(n_2087),
.B(n_1710),
.Y(n_3760)
);

OAI21x1_ASAP7_75t_L g3761 ( 
.A1(n_3678),
.A2(n_3657),
.B(n_3686),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3708),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3673),
.Y(n_3763)
);

AND2x4_ASAP7_75t_L g3764 ( 
.A(n_3722),
.B(n_1103),
.Y(n_3764)
);

OAI21x1_ASAP7_75t_L g3765 ( 
.A1(n_3694),
.A2(n_1106),
.B(n_1104),
.Y(n_3765)
);

OAI22xp5_ASAP7_75t_L g3766 ( 
.A1(n_3671),
.A2(n_1718),
.B1(n_1724),
.B2(n_1698),
.Y(n_3766)
);

NAND3xp33_ASAP7_75t_L g3767 ( 
.A(n_3658),
.B(n_1728),
.C(n_1726),
.Y(n_3767)
);

OAI21x1_ASAP7_75t_L g3768 ( 
.A1(n_3698),
.A2(n_1115),
.B(n_1112),
.Y(n_3768)
);

AO21x2_ASAP7_75t_L g3769 ( 
.A1(n_3660),
.A2(n_1749),
.B(n_1734),
.Y(n_3769)
);

BUFx3_ASAP7_75t_L g3770 ( 
.A(n_3653),
.Y(n_3770)
);

INVx3_ASAP7_75t_L g3771 ( 
.A(n_3734),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3730),
.Y(n_3772)
);

OAI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3689),
.A2(n_1755),
.B(n_1753),
.Y(n_3773)
);

AOI22xp33_ASAP7_75t_L g3774 ( 
.A1(n_3696),
.A2(n_3721),
.B1(n_3667),
.B2(n_3701),
.Y(n_3774)
);

CKINVDCx16_ASAP7_75t_R g3775 ( 
.A(n_3696),
.Y(n_3775)
);

BUFx12f_ASAP7_75t_L g3776 ( 
.A(n_3696),
.Y(n_3776)
);

OR2x2_ASAP7_75t_L g3777 ( 
.A(n_3738),
.B(n_28),
.Y(n_3777)
);

INVxp67_ASAP7_75t_SL g3778 ( 
.A(n_3725),
.Y(n_3778)
);

AO21x2_ASAP7_75t_L g3779 ( 
.A1(n_3695),
.A2(n_1767),
.B(n_1760),
.Y(n_3779)
);

AOI21xp5_ASAP7_75t_L g3780 ( 
.A1(n_3675),
.A2(n_1777),
.B(n_1774),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3672),
.B(n_28),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3740),
.Y(n_3782)
);

AOI22xp33_ASAP7_75t_L g3783 ( 
.A1(n_3685),
.A2(n_2036),
.B1(n_2038),
.B2(n_2030),
.Y(n_3783)
);

HB1xp67_ASAP7_75t_L g3784 ( 
.A(n_3646),
.Y(n_3784)
);

HB1xp67_ASAP7_75t_L g3785 ( 
.A(n_3646),
.Y(n_3785)
);

OAI21x1_ASAP7_75t_L g3786 ( 
.A1(n_3705),
.A2(n_1118),
.B(n_1117),
.Y(n_3786)
);

OAI211xp5_ASAP7_75t_L g3787 ( 
.A1(n_3648),
.A2(n_1805),
.B(n_1809),
.C(n_1800),
.Y(n_3787)
);

A2O1A1Ixp33_ASAP7_75t_L g3788 ( 
.A1(n_3703),
.A2(n_1919),
.B(n_1999),
.C(n_1858),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3735),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3735),
.Y(n_3790)
);

NAND2x1_ASAP7_75t_L g3791 ( 
.A(n_3680),
.B(n_29),
.Y(n_3791)
);

NAND2x1p5_ASAP7_75t_L g3792 ( 
.A(n_3717),
.B(n_1121),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3668),
.Y(n_3793)
);

OAI221xp5_ASAP7_75t_L g3794 ( 
.A1(n_3651),
.A2(n_1995),
.B1(n_1996),
.B2(n_1986),
.C(n_1955),
.Y(n_3794)
);

OAI21x1_ASAP7_75t_L g3795 ( 
.A1(n_3707),
.A2(n_1124),
.B(n_1123),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3670),
.Y(n_3796)
);

AOI22xp33_ASAP7_75t_SL g3797 ( 
.A1(n_3649),
.A2(n_1814),
.B1(n_1824),
.B2(n_1810),
.Y(n_3797)
);

NOR2xp67_ASAP7_75t_SL g3798 ( 
.A(n_3663),
.B(n_1828),
.Y(n_3798)
);

INVx3_ASAP7_75t_L g3799 ( 
.A(n_3729),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3691),
.B(n_29),
.Y(n_3800)
);

AOI22xp33_ASAP7_75t_SL g3801 ( 
.A1(n_3684),
.A2(n_1834),
.B1(n_1847),
.B2(n_1832),
.Y(n_3801)
);

OAI21x1_ASAP7_75t_SL g3802 ( 
.A1(n_3654),
.A2(n_3662),
.B(n_3661),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3681),
.Y(n_3803)
);

OAI21x1_ASAP7_75t_L g3804 ( 
.A1(n_3711),
.A2(n_1128),
.B(n_1127),
.Y(n_3804)
);

OAI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_3687),
.A2(n_1876),
.B(n_1862),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3681),
.Y(n_3806)
);

NOR2xp33_ASAP7_75t_L g3807 ( 
.A(n_3718),
.B(n_3741),
.Y(n_3807)
);

OA21x2_ASAP7_75t_L g3808 ( 
.A1(n_3739),
.A2(n_1891),
.B(n_1882),
.Y(n_3808)
);

OA21x2_ASAP7_75t_L g3809 ( 
.A1(n_3732),
.A2(n_1903),
.B(n_1897),
.Y(n_3809)
);

AOI22xp33_ASAP7_75t_L g3810 ( 
.A1(n_3709),
.A2(n_3697),
.B1(n_3699),
.B2(n_3683),
.Y(n_3810)
);

OA21x2_ASAP7_75t_L g3811 ( 
.A1(n_3731),
.A2(n_1935),
.B(n_1909),
.Y(n_3811)
);

OAI21x1_ASAP7_75t_L g3812 ( 
.A1(n_3710),
.A2(n_1133),
.B(n_1130),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3666),
.Y(n_3813)
);

INVx2_ASAP7_75t_SL g3814 ( 
.A(n_3727),
.Y(n_3814)
);

INVxp67_ASAP7_75t_SL g3815 ( 
.A(n_3659),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3666),
.Y(n_3816)
);

NOR2xp33_ASAP7_75t_L g3817 ( 
.A(n_3723),
.B(n_3736),
.Y(n_3817)
);

AO21x1_ASAP7_75t_L g3818 ( 
.A1(n_3677),
.A2(n_30),
.B(n_31),
.Y(n_3818)
);

OR2x2_ASAP7_75t_L g3819 ( 
.A(n_3702),
.B(n_3712),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3743),
.Y(n_3820)
);

INVx6_ASAP7_75t_L g3821 ( 
.A(n_3749),
.Y(n_3821)
);

AO21x1_ASAP7_75t_L g3822 ( 
.A1(n_3790),
.A2(n_3737),
.B(n_3728),
.Y(n_3822)
);

INVx2_ASAP7_75t_L g3823 ( 
.A(n_3744),
.Y(n_3823)
);

BUFx2_ASAP7_75t_R g3824 ( 
.A(n_3770),
.Y(n_3824)
);

INVx1_ASAP7_75t_SL g3825 ( 
.A(n_3814),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3750),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3751),
.Y(n_3827)
);

INVx2_ASAP7_75t_L g3828 ( 
.A(n_3755),
.Y(n_3828)
);

CKINVDCx11_ASAP7_75t_R g3829 ( 
.A(n_3776),
.Y(n_3829)
);

AOI21x1_ASAP7_75t_L g3830 ( 
.A1(n_3813),
.A2(n_3719),
.B(n_3713),
.Y(n_3830)
);

AOI22xp5_ASAP7_75t_L g3831 ( 
.A1(n_3775),
.A2(n_3720),
.B1(n_3724),
.B2(n_3714),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_3772),
.Y(n_3832)
);

AOI22xp33_ASAP7_75t_L g3833 ( 
.A1(n_3789),
.A2(n_3733),
.B1(n_3692),
.B2(n_3716),
.Y(n_3833)
);

AND2x2_ASAP7_75t_L g3834 ( 
.A(n_3763),
.B(n_3778),
.Y(n_3834)
);

AOI22xp33_ASAP7_75t_SL g3835 ( 
.A1(n_3742),
.A2(n_3664),
.B1(n_2011),
.B2(n_2014),
.Y(n_3835)
);

OAI22xp5_ASAP7_75t_L g3836 ( 
.A1(n_3774),
.A2(n_1947),
.B1(n_2060),
.B2(n_1937),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3762),
.Y(n_3837)
);

AND2x4_ASAP7_75t_L g3838 ( 
.A(n_3782),
.B(n_32),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3757),
.Y(n_3839)
);

BUFx2_ASAP7_75t_L g3840 ( 
.A(n_3748),
.Y(n_3840)
);

AOI22xp33_ASAP7_75t_L g3841 ( 
.A1(n_3818),
.A2(n_2065),
.B1(n_34),
.B2(n_32),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_3747),
.Y(n_3842)
);

BUFx6f_ASAP7_75t_L g3843 ( 
.A(n_3756),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3816),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3803),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3806),
.Y(n_3846)
);

INVxp67_ASAP7_75t_L g3847 ( 
.A(n_3815),
.Y(n_3847)
);

OAI21x1_ASAP7_75t_SL g3848 ( 
.A1(n_3802),
.A2(n_3760),
.B(n_3781),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3784),
.Y(n_3849)
);

BUFx2_ASAP7_75t_R g3850 ( 
.A(n_3771),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3785),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3793),
.Y(n_3852)
);

CKINVDCx11_ASAP7_75t_R g3853 ( 
.A(n_3796),
.Y(n_3853)
);

BUFx6f_ASAP7_75t_SL g3854 ( 
.A(n_3764),
.Y(n_3854)
);

BUFx2_ASAP7_75t_R g3855 ( 
.A(n_3819),
.Y(n_3855)
);

AOI22xp33_ASAP7_75t_SL g3856 ( 
.A1(n_3758),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_3856)
);

OAI22xp5_ASAP7_75t_L g3857 ( 
.A1(n_3767),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_3857)
);

BUFx3_ASAP7_75t_L g3858 ( 
.A(n_3746),
.Y(n_3858)
);

BUFx3_ASAP7_75t_L g3859 ( 
.A(n_3817),
.Y(n_3859)
);

AOI22xp33_ASAP7_75t_SL g3860 ( 
.A1(n_3811),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_3860)
);

INVx2_ASAP7_75t_SL g3861 ( 
.A(n_3777),
.Y(n_3861)
);

HB1xp67_ASAP7_75t_L g3862 ( 
.A(n_3799),
.Y(n_3862)
);

INVx2_ASAP7_75t_L g3863 ( 
.A(n_3753),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3768),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3765),
.Y(n_3865)
);

AOI22xp33_ASAP7_75t_L g3866 ( 
.A1(n_3807),
.A2(n_42),
.B1(n_38),
.B2(n_40),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3745),
.Y(n_3867)
);

BUFx12f_ASAP7_75t_L g3868 ( 
.A(n_3800),
.Y(n_3868)
);

OAI21x1_ASAP7_75t_L g3869 ( 
.A1(n_3761),
.A2(n_42),
.B(n_43),
.Y(n_3869)
);

INVx2_ASAP7_75t_L g3870 ( 
.A(n_3786),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3792),
.Y(n_3871)
);

AO21x2_ASAP7_75t_L g3872 ( 
.A1(n_3773),
.A2(n_43),
.B(n_45),
.Y(n_3872)
);

AOI21x1_ASAP7_75t_L g3873 ( 
.A1(n_3798),
.A2(n_3809),
.B(n_3808),
.Y(n_3873)
);

HB1xp67_ASAP7_75t_L g3874 ( 
.A(n_3811),
.Y(n_3874)
);

OAI22xp5_ASAP7_75t_L g3875 ( 
.A1(n_3791),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3759),
.Y(n_3876)
);

INVx1_ASAP7_75t_SL g3877 ( 
.A(n_3769),
.Y(n_3877)
);

AOI22xp33_ASAP7_75t_L g3878 ( 
.A1(n_3810),
.A2(n_50),
.B1(n_46),
.B2(n_48),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3795),
.Y(n_3879)
);

NAND2x1p5_ASAP7_75t_L g3880 ( 
.A(n_3752),
.B(n_48),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3804),
.Y(n_3881)
);

INVx2_ASAP7_75t_L g3882 ( 
.A(n_3812),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3779),
.Y(n_3883)
);

AO21x1_ASAP7_75t_SL g3884 ( 
.A1(n_3805),
.A2(n_51),
.B(n_52),
.Y(n_3884)
);

NAND2x1p5_ASAP7_75t_L g3885 ( 
.A(n_3780),
.B(n_52),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3754),
.Y(n_3886)
);

BUFx6f_ASAP7_75t_L g3887 ( 
.A(n_3787),
.Y(n_3887)
);

AOI22xp33_ASAP7_75t_L g3888 ( 
.A1(n_3766),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_3888)
);

INVx2_ASAP7_75t_L g3889 ( 
.A(n_3794),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3797),
.Y(n_3890)
);

AND2x2_ASAP7_75t_L g3891 ( 
.A(n_3783),
.B(n_53),
.Y(n_3891)
);

BUFx2_ASAP7_75t_SL g3892 ( 
.A(n_3801),
.Y(n_3892)
);

INVx6_ASAP7_75t_L g3893 ( 
.A(n_3788),
.Y(n_3893)
);

OAI22xp5_ASAP7_75t_L g3894 ( 
.A1(n_3774),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_3894)
);

INVx5_ASAP7_75t_L g3895 ( 
.A(n_3776),
.Y(n_3895)
);

AOI21x1_ASAP7_75t_L g3896 ( 
.A1(n_3813),
.A2(n_57),
.B(n_58),
.Y(n_3896)
);

AOI21x1_ASAP7_75t_L g3897 ( 
.A1(n_3813),
.A2(n_57),
.B(n_58),
.Y(n_3897)
);

BUFx2_ASAP7_75t_L g3898 ( 
.A(n_3748),
.Y(n_3898)
);

INVx6_ASAP7_75t_L g3899 ( 
.A(n_3749),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3750),
.B(n_59),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3743),
.Y(n_3901)
);

INVx4_ASAP7_75t_L g3902 ( 
.A(n_3749),
.Y(n_3902)
);

OAI22xp5_ASAP7_75t_L g3903 ( 
.A1(n_3831),
.A2(n_62),
.B1(n_59),
.B2(n_60),
.Y(n_3903)
);

AOI22xp33_ASAP7_75t_L g3904 ( 
.A1(n_3822),
.A2(n_66),
.B1(n_63),
.B2(n_64),
.Y(n_3904)
);

OAI21xp5_ASAP7_75t_SL g3905 ( 
.A1(n_3835),
.A2(n_3880),
.B(n_3841),
.Y(n_3905)
);

AOI22xp33_ASAP7_75t_L g3906 ( 
.A1(n_3889),
.A2(n_67),
.B1(n_63),
.B2(n_66),
.Y(n_3906)
);

INVx2_ASAP7_75t_SL g3907 ( 
.A(n_3821),
.Y(n_3907)
);

AOI22xp33_ASAP7_75t_L g3908 ( 
.A1(n_3892),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_3908)
);

OAI21xp5_ASAP7_75t_SL g3909 ( 
.A1(n_3866),
.A2(n_68),
.B(n_69),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3820),
.Y(n_3910)
);

OAI21xp5_ASAP7_75t_SL g3911 ( 
.A1(n_3875),
.A2(n_70),
.B(n_71),
.Y(n_3911)
);

OAI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_3876),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_3912)
);

AOI22xp33_ASAP7_75t_L g3913 ( 
.A1(n_3893),
.A2(n_75),
.B1(n_72),
.B2(n_73),
.Y(n_3913)
);

AND2x2_ASAP7_75t_L g3914 ( 
.A(n_3840),
.B(n_73),
.Y(n_3914)
);

OAI21xp5_ASAP7_75t_SL g3915 ( 
.A1(n_3885),
.A2(n_76),
.B(n_77),
.Y(n_3915)
);

AOI22xp33_ASAP7_75t_L g3916 ( 
.A1(n_3883),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3847),
.B(n_78),
.Y(n_3917)
);

INVx4_ASAP7_75t_L g3918 ( 
.A(n_3829),
.Y(n_3918)
);

AOI22xp33_ASAP7_75t_L g3919 ( 
.A1(n_3890),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_3919)
);

AOI22xp33_ASAP7_75t_L g3920 ( 
.A1(n_3877),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_3920)
);

BUFx6f_ASAP7_75t_L g3921 ( 
.A(n_3895),
.Y(n_3921)
);

BUFx12f_ASAP7_75t_L g3922 ( 
.A(n_3895),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3901),
.Y(n_3923)
);

AOI22xp5_ASAP7_75t_L g3924 ( 
.A1(n_3894),
.A2(n_85),
.B1(n_82),
.B2(n_83),
.Y(n_3924)
);

AOI22xp33_ASAP7_75t_L g3925 ( 
.A1(n_3860),
.A2(n_86),
.B1(n_82),
.B2(n_85),
.Y(n_3925)
);

OAI21xp33_ASAP7_75t_L g3926 ( 
.A1(n_3867),
.A2(n_3886),
.B(n_3874),
.Y(n_3926)
);

OAI22xp33_ASAP7_75t_L g3927 ( 
.A1(n_3859),
.A2(n_3861),
.B1(n_3871),
.B2(n_3825),
.Y(n_3927)
);

INVx6_ASAP7_75t_L g3928 ( 
.A(n_3902),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3898),
.B(n_86),
.Y(n_3929)
);

BUFx12f_ASAP7_75t_L g3930 ( 
.A(n_3899),
.Y(n_3930)
);

AOI22xp33_ASAP7_75t_SL g3931 ( 
.A1(n_3836),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3823),
.Y(n_3932)
);

AOI22xp33_ASAP7_75t_L g3933 ( 
.A1(n_3884),
.A2(n_91),
.B1(n_88),
.B2(n_90),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3852),
.B(n_91),
.Y(n_3934)
);

BUFx10_ASAP7_75t_L g3935 ( 
.A(n_3854),
.Y(n_3935)
);

AOI22xp33_ASAP7_75t_L g3936 ( 
.A1(n_3872),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_3936)
);

OAI22xp33_ASAP7_75t_L g3937 ( 
.A1(n_3868),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3837),
.Y(n_3938)
);

AOI22xp33_ASAP7_75t_SL g3939 ( 
.A1(n_3848),
.A2(n_99),
.B1(n_96),
.B2(n_98),
.Y(n_3939)
);

AOI22xp33_ASAP7_75t_SL g3940 ( 
.A1(n_3891),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_3940)
);

INVx6_ASAP7_75t_L g3941 ( 
.A(n_3843),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3834),
.B(n_100),
.Y(n_3942)
);

AND2x2_ASAP7_75t_L g3943 ( 
.A(n_3826),
.B(n_101),
.Y(n_3943)
);

AOI22xp33_ASAP7_75t_L g3944 ( 
.A1(n_3833),
.A2(n_3878),
.B1(n_3857),
.B2(n_3864),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3832),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3900),
.B(n_101),
.Y(n_3946)
);

INVxp67_ASAP7_75t_L g3947 ( 
.A(n_3858),
.Y(n_3947)
);

INVx5_ASAP7_75t_SL g3948 ( 
.A(n_3887),
.Y(n_3948)
);

OAI22xp5_ASAP7_75t_SL g3949 ( 
.A1(n_3855),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3844),
.B(n_102),
.Y(n_3950)
);

AOI22xp33_ASAP7_75t_L g3951 ( 
.A1(n_3870),
.A2(n_106),
.B1(n_103),
.B2(n_105),
.Y(n_3951)
);

OAI22xp5_ASAP7_75t_L g3952 ( 
.A1(n_3888),
.A2(n_109),
.B1(n_105),
.B2(n_108),
.Y(n_3952)
);

BUFx3_ASAP7_75t_L g3953 ( 
.A(n_3853),
.Y(n_3953)
);

AOI22xp33_ASAP7_75t_SL g3954 ( 
.A1(n_3838),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_3954)
);

OAI21xp33_ASAP7_75t_L g3955 ( 
.A1(n_3862),
.A2(n_110),
.B(n_111),
.Y(n_3955)
);

OR2x2_ASAP7_75t_L g3956 ( 
.A(n_3849),
.B(n_112),
.Y(n_3956)
);

AOI22xp33_ASAP7_75t_L g3957 ( 
.A1(n_3879),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_3957)
);

AOI22xp33_ASAP7_75t_SL g3958 ( 
.A1(n_3887),
.A2(n_116),
.B1(n_113),
.B2(n_115),
.Y(n_3958)
);

AOI22xp33_ASAP7_75t_L g3959 ( 
.A1(n_3881),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_3959)
);

NOR2xp33_ASAP7_75t_L g3960 ( 
.A(n_3824),
.B(n_117),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3850),
.B(n_118),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3851),
.Y(n_3962)
);

OAI21xp5_ASAP7_75t_SL g3963 ( 
.A1(n_3856),
.A2(n_118),
.B(n_119),
.Y(n_3963)
);

OAI21xp33_ASAP7_75t_L g3964 ( 
.A1(n_3865),
.A2(n_120),
.B(n_121),
.Y(n_3964)
);

BUFx12f_ASAP7_75t_L g3965 ( 
.A(n_3843),
.Y(n_3965)
);

INVx3_ASAP7_75t_L g3966 ( 
.A(n_3828),
.Y(n_3966)
);

OAI22xp5_ASAP7_75t_SL g3967 ( 
.A1(n_3882),
.A2(n_3863),
.B1(n_3873),
.B2(n_3839),
.Y(n_3967)
);

AOI22xp33_ASAP7_75t_L g3968 ( 
.A1(n_3827),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_3968)
);

AOI22xp33_ASAP7_75t_L g3969 ( 
.A1(n_3845),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_3969)
);

BUFx6f_ASAP7_75t_L g3970 ( 
.A(n_3869),
.Y(n_3970)
);

AOI22xp33_ASAP7_75t_SL g3971 ( 
.A1(n_3846),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_3971)
);

OR2x6_ASAP7_75t_L g3972 ( 
.A(n_3922),
.B(n_3896),
.Y(n_3972)
);

BUFx10_ASAP7_75t_L g3973 ( 
.A(n_3921),
.Y(n_3973)
);

AND2x4_ASAP7_75t_L g3974 ( 
.A(n_3947),
.B(n_3897),
.Y(n_3974)
);

AND2x4_ASAP7_75t_L g3975 ( 
.A(n_3918),
.B(n_3830),
.Y(n_3975)
);

NOR2xp33_ASAP7_75t_R g3976 ( 
.A(n_3953),
.B(n_125),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3942),
.B(n_3842),
.Y(n_3977)
);

INVx2_ASAP7_75t_L g3978 ( 
.A(n_3970),
.Y(n_3978)
);

NOR2xp33_ASAP7_75t_R g3979 ( 
.A(n_3921),
.B(n_126),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3910),
.Y(n_3980)
);

HB1xp67_ASAP7_75t_L g3981 ( 
.A(n_3923),
.Y(n_3981)
);

NOR2xp33_ASAP7_75t_R g3982 ( 
.A(n_3930),
.B(n_127),
.Y(n_3982)
);

NOR2xp33_ASAP7_75t_L g3983 ( 
.A(n_3928),
.B(n_128),
.Y(n_3983)
);

AND2x2_ASAP7_75t_L g3984 ( 
.A(n_3935),
.B(n_128),
.Y(n_3984)
);

INVxp67_ASAP7_75t_L g3985 ( 
.A(n_3960),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3938),
.Y(n_3986)
);

BUFx6f_ASAP7_75t_L g3987 ( 
.A(n_3965),
.Y(n_3987)
);

NAND2xp33_ASAP7_75t_R g3988 ( 
.A(n_3961),
.B(n_131),
.Y(n_3988)
);

AND2x4_ASAP7_75t_L g3989 ( 
.A(n_3907),
.B(n_129),
.Y(n_3989)
);

AND2x2_ASAP7_75t_L g3990 ( 
.A(n_3926),
.B(n_129),
.Y(n_3990)
);

NAND2xp33_ASAP7_75t_R g3991 ( 
.A(n_3914),
.B(n_3929),
.Y(n_3991)
);

NAND2xp33_ASAP7_75t_R g3992 ( 
.A(n_3943),
.B(n_3956),
.Y(n_3992)
);

CKINVDCx20_ASAP7_75t_R g3993 ( 
.A(n_3949),
.Y(n_3993)
);

XOR2xp5_ASAP7_75t_L g3994 ( 
.A(n_3903),
.B(n_131),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3928),
.B(n_132),
.Y(n_3995)
);

BUFx3_ASAP7_75t_L g3996 ( 
.A(n_3941),
.Y(n_3996)
);

XNOR2xp5_ASAP7_75t_L g3997 ( 
.A(n_3927),
.B(n_132),
.Y(n_3997)
);

BUFx10_ASAP7_75t_L g3998 ( 
.A(n_3941),
.Y(n_3998)
);

INVxp67_ASAP7_75t_L g3999 ( 
.A(n_3967),
.Y(n_3999)
);

INVx2_ASAP7_75t_L g4000 ( 
.A(n_3970),
.Y(n_4000)
);

NAND2xp33_ASAP7_75t_R g4001 ( 
.A(n_3917),
.B(n_134),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3945),
.Y(n_4002)
);

XNOR2xp5_ASAP7_75t_L g4003 ( 
.A(n_3937),
.B(n_133),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_L g4004 ( 
.A(n_3934),
.B(n_133),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3950),
.B(n_3946),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_SL g4006 ( 
.A(n_3962),
.B(n_134),
.Y(n_4006)
);

AND2x4_ASAP7_75t_L g4007 ( 
.A(n_3966),
.B(n_135),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_3932),
.Y(n_4008)
);

NOR2xp33_ASAP7_75t_L g4009 ( 
.A(n_3905),
.B(n_135),
.Y(n_4009)
);

NOR2xp33_ASAP7_75t_R g4010 ( 
.A(n_3933),
.B(n_136),
.Y(n_4010)
);

NOR2xp33_ASAP7_75t_R g4011 ( 
.A(n_3908),
.B(n_136),
.Y(n_4011)
);

AND2x4_ASAP7_75t_L g4012 ( 
.A(n_3944),
.B(n_137),
.Y(n_4012)
);

BUFx10_ASAP7_75t_L g4013 ( 
.A(n_3948),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3904),
.B(n_138),
.Y(n_4014)
);

NOR2xp33_ASAP7_75t_R g4015 ( 
.A(n_3913),
.B(n_138),
.Y(n_4015)
);

NAND2xp33_ASAP7_75t_R g4016 ( 
.A(n_3948),
.B(n_141),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_3955),
.B(n_140),
.Y(n_4017)
);

OR2x6_ASAP7_75t_L g4018 ( 
.A(n_3915),
.B(n_141),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3964),
.B(n_142),
.Y(n_4019)
);

HB1xp67_ASAP7_75t_L g4020 ( 
.A(n_3912),
.Y(n_4020)
);

OR2x6_ASAP7_75t_L g4021 ( 
.A(n_3911),
.B(n_142),
.Y(n_4021)
);

INVxp67_ASAP7_75t_L g4022 ( 
.A(n_3939),
.Y(n_4022)
);

NAND2xp33_ASAP7_75t_R g4023 ( 
.A(n_3963),
.B(n_144),
.Y(n_4023)
);

BUFx3_ASAP7_75t_L g4024 ( 
.A(n_3924),
.Y(n_4024)
);

CKINVDCx5p33_ASAP7_75t_R g4025 ( 
.A(n_3958),
.Y(n_4025)
);

NAND2xp33_ASAP7_75t_R g4026 ( 
.A(n_3909),
.B(n_144),
.Y(n_4026)
);

AND2x4_ASAP7_75t_L g4027 ( 
.A(n_3936),
.B(n_143),
.Y(n_4027)
);

NOR2xp33_ASAP7_75t_R g4028 ( 
.A(n_3919),
.B(n_143),
.Y(n_4028)
);

BUFx10_ASAP7_75t_L g4029 ( 
.A(n_3954),
.Y(n_4029)
);

CKINVDCx20_ASAP7_75t_R g4030 ( 
.A(n_3952),
.Y(n_4030)
);

NAND2xp33_ASAP7_75t_R g4031 ( 
.A(n_3940),
.B(n_147),
.Y(n_4031)
);

AND2x4_ASAP7_75t_L g4032 ( 
.A(n_3969),
.B(n_145),
.Y(n_4032)
);

NOR2xp33_ASAP7_75t_R g4033 ( 
.A(n_3959),
.B(n_147),
.Y(n_4033)
);

INVxp67_ASAP7_75t_L g4034 ( 
.A(n_3971),
.Y(n_4034)
);

NAND2xp33_ASAP7_75t_R g4035 ( 
.A(n_3931),
.B(n_149),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_3920),
.Y(n_4036)
);

BUFx10_ASAP7_75t_L g4037 ( 
.A(n_3951),
.Y(n_4037)
);

AND2x4_ASAP7_75t_L g4038 ( 
.A(n_3968),
.B(n_148),
.Y(n_4038)
);

AND2x4_ASAP7_75t_L g4039 ( 
.A(n_3957),
.B(n_148),
.Y(n_4039)
);

NAND2xp33_ASAP7_75t_R g4040 ( 
.A(n_3925),
.B(n_150),
.Y(n_4040)
);

CKINVDCx20_ASAP7_75t_R g4041 ( 
.A(n_3906),
.Y(n_4041)
);

NAND2xp33_ASAP7_75t_R g4042 ( 
.A(n_3916),
.B(n_150),
.Y(n_4042)
);

NAND2xp33_ASAP7_75t_R g4043 ( 
.A(n_3961),
.B(n_151),
.Y(n_4043)
);

NOR2xp33_ASAP7_75t_R g4044 ( 
.A(n_3922),
.B(n_149),
.Y(n_4044)
);

CKINVDCx20_ASAP7_75t_R g4045 ( 
.A(n_3953),
.Y(n_4045)
);

NAND2xp33_ASAP7_75t_R g4046 ( 
.A(n_3961),
.B(n_152),
.Y(n_4046)
);

OR2x6_ASAP7_75t_L g4047 ( 
.A(n_3922),
.B(n_151),
.Y(n_4047)
);

NOR2xp33_ASAP7_75t_R g4048 ( 
.A(n_3922),
.B(n_152),
.Y(n_4048)
);

INVxp67_ASAP7_75t_L g4049 ( 
.A(n_3960),
.Y(n_4049)
);

NAND2xp33_ASAP7_75t_R g4050 ( 
.A(n_3961),
.B(n_154),
.Y(n_4050)
);

NAND2xp33_ASAP7_75t_R g4051 ( 
.A(n_3961),
.B(n_154),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3926),
.B(n_153),
.Y(n_4052)
);

NAND2xp33_ASAP7_75t_R g4053 ( 
.A(n_3961),
.B(n_155),
.Y(n_4053)
);

NOR2xp33_ASAP7_75t_R g4054 ( 
.A(n_3922),
.B(n_153),
.Y(n_4054)
);

INVxp67_ASAP7_75t_L g4055 ( 
.A(n_3960),
.Y(n_4055)
);

NAND2xp33_ASAP7_75t_R g4056 ( 
.A(n_3961),
.B(n_156),
.Y(n_4056)
);

NAND2xp33_ASAP7_75t_R g4057 ( 
.A(n_3961),
.B(n_157),
.Y(n_4057)
);

INVx1_ASAP7_75t_SL g4058 ( 
.A(n_3953),
.Y(n_4058)
);

BUFx8_ASAP7_75t_SL g4059 ( 
.A(n_3922),
.Y(n_4059)
);

AND2x4_ASAP7_75t_L g4060 ( 
.A(n_3947),
.B(n_155),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3926),
.B(n_157),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3910),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3926),
.B(n_158),
.Y(n_4063)
);

NAND2xp33_ASAP7_75t_R g4064 ( 
.A(n_3961),
.B(n_159),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3970),
.Y(n_4065)
);

NAND2xp33_ASAP7_75t_R g4066 ( 
.A(n_3961),
.B(n_159),
.Y(n_4066)
);

AND2x4_ASAP7_75t_L g4067 ( 
.A(n_3947),
.B(n_158),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3910),
.Y(n_4068)
);

BUFx3_ASAP7_75t_L g4069 ( 
.A(n_3953),
.Y(n_4069)
);

NOR2xp33_ASAP7_75t_R g4070 ( 
.A(n_3922),
.B(n_160),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3910),
.Y(n_4071)
);

AND2x4_ASAP7_75t_L g4072 ( 
.A(n_3947),
.B(n_161),
.Y(n_4072)
);

NOR2xp33_ASAP7_75t_R g4073 ( 
.A(n_3922),
.B(n_161),
.Y(n_4073)
);

XOR2xp5_ASAP7_75t_L g4074 ( 
.A(n_3949),
.B(n_162),
.Y(n_4074)
);

NAND2xp33_ASAP7_75t_R g4075 ( 
.A(n_3961),
.B(n_164),
.Y(n_4075)
);

AND2x4_ASAP7_75t_L g4076 ( 
.A(n_3947),
.B(n_162),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3910),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3970),
.Y(n_4078)
);

NOR2xp33_ASAP7_75t_R g4079 ( 
.A(n_3922),
.B(n_165),
.Y(n_4079)
);

BUFx10_ASAP7_75t_L g4080 ( 
.A(n_3921),
.Y(n_4080)
);

NOR2xp33_ASAP7_75t_R g4081 ( 
.A(n_3922),
.B(n_165),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3926),
.B(n_166),
.Y(n_4082)
);

XNOR2xp5_ASAP7_75t_L g4083 ( 
.A(n_3949),
.B(n_166),
.Y(n_4083)
);

CKINVDCx5p33_ASAP7_75t_R g4084 ( 
.A(n_3930),
.Y(n_4084)
);

AND2x4_ASAP7_75t_L g4085 ( 
.A(n_3947),
.B(n_167),
.Y(n_4085)
);

INVxp67_ASAP7_75t_L g4086 ( 
.A(n_3960),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3910),
.Y(n_4087)
);

AND2x2_ASAP7_75t_L g4088 ( 
.A(n_3947),
.B(n_167),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3981),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3980),
.Y(n_4090)
);

INVx2_ASAP7_75t_L g4091 ( 
.A(n_3974),
.Y(n_4091)
);

AND2x2_ASAP7_75t_L g4092 ( 
.A(n_3975),
.B(n_168),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_3978),
.Y(n_4093)
);

OR2x2_ASAP7_75t_L g4094 ( 
.A(n_4002),
.B(n_168),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_4020),
.B(n_169),
.Y(n_4095)
);

AND2x2_ASAP7_75t_L g4096 ( 
.A(n_3996),
.B(n_170),
.Y(n_4096)
);

INVxp67_ASAP7_75t_L g4097 ( 
.A(n_3991),
.Y(n_4097)
);

AND2x2_ASAP7_75t_L g4098 ( 
.A(n_3998),
.B(n_170),
.Y(n_4098)
);

AND2x4_ASAP7_75t_L g4099 ( 
.A(n_4069),
.B(n_171),
.Y(n_4099)
);

AND2x4_ASAP7_75t_L g4100 ( 
.A(n_4007),
.B(n_4058),
.Y(n_4100)
);

INVx1_ASAP7_75t_SL g4101 ( 
.A(n_4045),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3986),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_3990),
.B(n_171),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_4062),
.Y(n_4104)
);

INVx2_ASAP7_75t_L g4105 ( 
.A(n_4000),
.Y(n_4105)
);

OR2x2_ASAP7_75t_L g4106 ( 
.A(n_4068),
.B(n_172),
.Y(n_4106)
);

HB1xp67_ASAP7_75t_L g4107 ( 
.A(n_4071),
.Y(n_4107)
);

AND2x2_ASAP7_75t_L g4108 ( 
.A(n_4005),
.B(n_172),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_4077),
.B(n_4087),
.Y(n_4109)
);

OR2x2_ASAP7_75t_L g4110 ( 
.A(n_4065),
.B(n_173),
.Y(n_4110)
);

AND2x4_ASAP7_75t_L g4111 ( 
.A(n_4078),
.B(n_173),
.Y(n_4111)
);

AND2x2_ASAP7_75t_L g4112 ( 
.A(n_3973),
.B(n_174),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_4052),
.B(n_4061),
.Y(n_4113)
);

OR2x2_ASAP7_75t_L g4114 ( 
.A(n_4063),
.B(n_174),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_4008),
.Y(n_4115)
);

INVxp67_ASAP7_75t_SL g4116 ( 
.A(n_3999),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_L g4117 ( 
.A(n_4082),
.B(n_175),
.Y(n_4117)
);

BUFx3_ASAP7_75t_L g4118 ( 
.A(n_4059),
.Y(n_4118)
);

INVx2_ASAP7_75t_L g4119 ( 
.A(n_3972),
.Y(n_4119)
);

AND2x2_ASAP7_75t_L g4120 ( 
.A(n_4080),
.B(n_175),
.Y(n_4120)
);

AND2x2_ASAP7_75t_L g4121 ( 
.A(n_4013),
.B(n_176),
.Y(n_4121)
);

INVx2_ASAP7_75t_L g4122 ( 
.A(n_3972),
.Y(n_4122)
);

OR2x2_ASAP7_75t_L g4123 ( 
.A(n_4024),
.B(n_177),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3977),
.Y(n_4124)
);

INVx2_ASAP7_75t_L g4125 ( 
.A(n_4036),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4004),
.Y(n_4126)
);

INVx2_ASAP7_75t_SL g4127 ( 
.A(n_3987),
.Y(n_4127)
);

OR2x2_ASAP7_75t_L g4128 ( 
.A(n_4022),
.B(n_177),
.Y(n_4128)
);

BUFx3_ASAP7_75t_L g4129 ( 
.A(n_4084),
.Y(n_4129)
);

OR2x2_ASAP7_75t_L g4130 ( 
.A(n_4021),
.B(n_178),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_4012),
.B(n_178),
.Y(n_4131)
);

INVx3_ASAP7_75t_L g4132 ( 
.A(n_3987),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_4006),
.Y(n_4133)
);

INVx2_ASAP7_75t_L g4134 ( 
.A(n_3995),
.Y(n_4134)
);

BUFx6f_ASAP7_75t_L g4135 ( 
.A(n_4047),
.Y(n_4135)
);

AND2x2_ASAP7_75t_L g4136 ( 
.A(n_4060),
.B(n_179),
.Y(n_4136)
);

OA21x2_ASAP7_75t_L g4137 ( 
.A1(n_3985),
.A2(n_179),
.B(n_180),
.Y(n_4137)
);

AOI22xp5_ASAP7_75t_L g4138 ( 
.A1(n_4026),
.A2(n_4023),
.B1(n_4042),
.B2(n_4009),
.Y(n_4138)
);

AND2x2_ASAP7_75t_L g4139 ( 
.A(n_4067),
.B(n_181),
.Y(n_4139)
);

AND2x2_ASAP7_75t_L g4140 ( 
.A(n_4072),
.B(n_181),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4088),
.Y(n_4141)
);

INVx2_ASAP7_75t_L g4142 ( 
.A(n_3989),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_4034),
.B(n_182),
.Y(n_4143)
);

INVx2_ASAP7_75t_SL g4144 ( 
.A(n_4076),
.Y(n_4144)
);

OR2x2_ASAP7_75t_L g4145 ( 
.A(n_4021),
.B(n_183),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_4037),
.Y(n_4146)
);

HB1xp67_ASAP7_75t_L g4147 ( 
.A(n_3992),
.Y(n_4147)
);

OR2x2_ASAP7_75t_L g4148 ( 
.A(n_4018),
.B(n_185),
.Y(n_4148)
);

INVx2_ASAP7_75t_L g4149 ( 
.A(n_4085),
.Y(n_4149)
);

AND2x4_ASAP7_75t_L g4150 ( 
.A(n_3984),
.B(n_185),
.Y(n_4150)
);

OR2x2_ASAP7_75t_L g4151 ( 
.A(n_4018),
.B(n_186),
.Y(n_4151)
);

BUFx2_ASAP7_75t_L g4152 ( 
.A(n_3976),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_4019),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_4017),
.Y(n_4154)
);

AND2x2_ASAP7_75t_L g4155 ( 
.A(n_3983),
.B(n_186),
.Y(n_4155)
);

AOI22xp33_ASAP7_75t_L g4156 ( 
.A1(n_4041),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_4156)
);

INVx2_ASAP7_75t_L g4157 ( 
.A(n_4029),
.Y(n_4157)
);

OAI211xp5_ASAP7_75t_SL g4158 ( 
.A1(n_4014),
.A2(n_192),
.B(n_189),
.C(n_191),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_4030),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_3997),
.B(n_193),
.Y(n_4160)
);

AND2x2_ASAP7_75t_L g4161 ( 
.A(n_4047),
.B(n_193),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_4049),
.B(n_194),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4003),
.Y(n_4163)
);

BUFx2_ASAP7_75t_L g4164 ( 
.A(n_3979),
.Y(n_4164)
);

AND2x2_ASAP7_75t_L g4165 ( 
.A(n_4055),
.B(n_194),
.Y(n_4165)
);

INVx2_ASAP7_75t_L g4166 ( 
.A(n_4086),
.Y(n_4166)
);

OAI22xp5_ASAP7_75t_L g4167 ( 
.A1(n_4025),
.A2(n_198),
.B1(n_195),
.B2(n_197),
.Y(n_4167)
);

INVx2_ASAP7_75t_L g4168 ( 
.A(n_4027),
.Y(n_4168)
);

INVx2_ASAP7_75t_L g4169 ( 
.A(n_4032),
.Y(n_4169)
);

AND2x2_ASAP7_75t_L g4170 ( 
.A(n_3982),
.B(n_195),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3994),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_4083),
.B(n_198),
.Y(n_4172)
);

AOI21xp5_ASAP7_75t_L g4173 ( 
.A1(n_4074),
.A2(n_199),
.B(n_202),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_L g4174 ( 
.A(n_4038),
.B(n_4039),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4010),
.Y(n_4175)
);

AND2x2_ASAP7_75t_L g4176 ( 
.A(n_4044),
.B(n_199),
.Y(n_4176)
);

INVx3_ASAP7_75t_L g4177 ( 
.A(n_4016),
.Y(n_4177)
);

AND2x2_ASAP7_75t_L g4178 ( 
.A(n_4048),
.B(n_202),
.Y(n_4178)
);

INVx2_ASAP7_75t_L g4179 ( 
.A(n_3993),
.Y(n_4179)
);

BUFx2_ASAP7_75t_L g4180 ( 
.A(n_4054),
.Y(n_4180)
);

HB1xp67_ASAP7_75t_L g4181 ( 
.A(n_4001),
.Y(n_4181)
);

OR2x2_ASAP7_75t_L g4182 ( 
.A(n_4035),
.B(n_203),
.Y(n_4182)
);

AND2x2_ASAP7_75t_L g4183 ( 
.A(n_4070),
.B(n_203),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4033),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_3988),
.Y(n_4185)
);

OR2x2_ASAP7_75t_L g4186 ( 
.A(n_4043),
.B(n_204),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_4073),
.B(n_204),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4015),
.Y(n_4188)
);

BUFx2_ASAP7_75t_L g4189 ( 
.A(n_4079),
.Y(n_4189)
);

INVx2_ASAP7_75t_L g4190 ( 
.A(n_4046),
.Y(n_4190)
);

AND2x4_ASAP7_75t_L g4191 ( 
.A(n_4081),
.B(n_4050),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_4028),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4011),
.Y(n_4193)
);

INVx3_ASAP7_75t_L g4194 ( 
.A(n_4051),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_4053),
.Y(n_4195)
);

AND2x4_ASAP7_75t_L g4196 ( 
.A(n_4056),
.B(n_4057),
.Y(n_4196)
);

AOI22xp33_ASAP7_75t_L g4197 ( 
.A1(n_4064),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_4197)
);

CKINVDCx5p33_ASAP7_75t_R g4198 ( 
.A(n_4066),
.Y(n_4198)
);

A2O1A1Ixp33_ASAP7_75t_L g4199 ( 
.A1(n_4075),
.A2(n_209),
.B(n_206),
.C(n_208),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4031),
.Y(n_4200)
);

HB1xp67_ASAP7_75t_L g4201 ( 
.A(n_4040),
.Y(n_4201)
);

INVx2_ASAP7_75t_L g4202 ( 
.A(n_3974),
.Y(n_4202)
);

OR2x2_ASAP7_75t_L g4203 ( 
.A(n_3981),
.B(n_208),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_3981),
.Y(n_4204)
);

INVx4_ASAP7_75t_L g4205 ( 
.A(n_4059),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_3981),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_3975),
.B(n_209),
.Y(n_4207)
);

AND2x2_ASAP7_75t_L g4208 ( 
.A(n_3975),
.B(n_210),
.Y(n_4208)
);

AND2x2_ASAP7_75t_L g4209 ( 
.A(n_3975),
.B(n_210),
.Y(n_4209)
);

OR2x2_ASAP7_75t_L g4210 ( 
.A(n_3981),
.B(n_211),
.Y(n_4210)
);

INVx2_ASAP7_75t_SL g4211 ( 
.A(n_4013),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_4020),
.B(n_211),
.Y(n_4212)
);

BUFx12f_ASAP7_75t_L g4213 ( 
.A(n_4047),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_3981),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_3981),
.Y(n_4215)
);

BUFx2_ASAP7_75t_SL g4216 ( 
.A(n_4045),
.Y(n_4216)
);

AND2x2_ASAP7_75t_L g4217 ( 
.A(n_3975),
.B(n_212),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_3981),
.Y(n_4218)
);

INVxp67_ASAP7_75t_L g4219 ( 
.A(n_3991),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4020),
.B(n_212),
.Y(n_4220)
);

OR2x2_ASAP7_75t_L g4221 ( 
.A(n_3981),
.B(n_213),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_3981),
.Y(n_4222)
);

BUFx2_ASAP7_75t_L g4223 ( 
.A(n_4059),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_3974),
.Y(n_4224)
);

AND2x2_ASAP7_75t_L g4225 ( 
.A(n_3975),
.B(n_213),
.Y(n_4225)
);

AND2x4_ASAP7_75t_L g4226 ( 
.A(n_3996),
.B(n_214),
.Y(n_4226)
);

BUFx2_ASAP7_75t_L g4227 ( 
.A(n_4059),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_3981),
.Y(n_4228)
);

INVx2_ASAP7_75t_SL g4229 ( 
.A(n_4013),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_3981),
.Y(n_4230)
);

HB1xp67_ASAP7_75t_L g4231 ( 
.A(n_3981),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_3981),
.Y(n_4232)
);

NAND3xp33_ASAP7_75t_L g4233 ( 
.A(n_4026),
.B(n_214),
.C(n_215),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_3981),
.Y(n_4234)
);

INVxp67_ASAP7_75t_L g4235 ( 
.A(n_3991),
.Y(n_4235)
);

BUFx2_ASAP7_75t_L g4236 ( 
.A(n_4059),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_3981),
.Y(n_4237)
);

OAI21xp5_ASAP7_75t_L g4238 ( 
.A1(n_4009),
.A2(n_216),
.B(n_217),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_3974),
.Y(n_4239)
);

NAND2x1p5_ASAP7_75t_L g4240 ( 
.A(n_4007),
.B(n_216),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_4020),
.B(n_218),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_3975),
.B(n_219),
.Y(n_4242)
);

AO21x2_ASAP7_75t_L g4243 ( 
.A1(n_3999),
.A2(n_220),
.B(n_221),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_3974),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_3981),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_3974),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_3981),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_3981),
.Y(n_4248)
);

OAI21xp33_ASAP7_75t_L g4249 ( 
.A1(n_4116),
.A2(n_220),
.B(n_223),
.Y(n_4249)
);

AND2x2_ASAP7_75t_L g4250 ( 
.A(n_4091),
.B(n_224),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4095),
.B(n_224),
.Y(n_4251)
);

AND2x4_ASAP7_75t_L g4252 ( 
.A(n_4211),
.B(n_226),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4107),
.Y(n_4253)
);

INVxp67_ASAP7_75t_SL g4254 ( 
.A(n_4181),
.Y(n_4254)
);

AND2x2_ASAP7_75t_L g4255 ( 
.A(n_4202),
.B(n_227),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_SL g4256 ( 
.A(n_4159),
.B(n_227),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_4109),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4090),
.Y(n_4258)
);

AND2x2_ASAP7_75t_L g4259 ( 
.A(n_4224),
.B(n_228),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_4166),
.B(n_229),
.Y(n_4260)
);

AOI22xp33_ASAP7_75t_SL g4261 ( 
.A1(n_4147),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_4126),
.B(n_230),
.Y(n_4262)
);

HB1xp67_ASAP7_75t_L g4263 ( 
.A(n_4231),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4102),
.Y(n_4264)
);

AND2x2_ASAP7_75t_L g4265 ( 
.A(n_4239),
.B(n_231),
.Y(n_4265)
);

AND2x2_ASAP7_75t_L g4266 ( 
.A(n_4244),
.B(n_232),
.Y(n_4266)
);

AND2x4_ASAP7_75t_L g4267 ( 
.A(n_4229),
.B(n_232),
.Y(n_4267)
);

INVx5_ASAP7_75t_L g4268 ( 
.A(n_4205),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4104),
.Y(n_4269)
);

INVx3_ASAP7_75t_L g4270 ( 
.A(n_4118),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_4194),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4089),
.Y(n_4272)
);

NOR2xp33_ASAP7_75t_L g4273 ( 
.A(n_4223),
.B(n_233),
.Y(n_4273)
);

OR2x2_ASAP7_75t_L g4274 ( 
.A(n_4204),
.B(n_233),
.Y(n_4274)
);

INVx2_ASAP7_75t_L g4275 ( 
.A(n_4185),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4206),
.Y(n_4276)
);

AND2x4_ASAP7_75t_L g4277 ( 
.A(n_4100),
.B(n_234),
.Y(n_4277)
);

OR2x2_ASAP7_75t_L g4278 ( 
.A(n_4214),
.B(n_234),
.Y(n_4278)
);

AND2x2_ASAP7_75t_L g4279 ( 
.A(n_4246),
.B(n_235),
.Y(n_4279)
);

BUFx3_ASAP7_75t_L g4280 ( 
.A(n_4227),
.Y(n_4280)
);

INVx1_ASAP7_75t_SL g4281 ( 
.A(n_4216),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4215),
.Y(n_4282)
);

AND2x4_ASAP7_75t_L g4283 ( 
.A(n_4144),
.B(n_4236),
.Y(n_4283)
);

INVx2_ASAP7_75t_L g4284 ( 
.A(n_4190),
.Y(n_4284)
);

AND2x2_ASAP7_75t_L g4285 ( 
.A(n_4141),
.B(n_235),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4119),
.B(n_236),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4122),
.B(n_236),
.Y(n_4287)
);

INVx2_ASAP7_75t_L g4288 ( 
.A(n_4195),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_4218),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4222),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4228),
.Y(n_4291)
);

AND2x2_ASAP7_75t_L g4292 ( 
.A(n_4092),
.B(n_4207),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4230),
.Y(n_4293)
);

INVx1_ASAP7_75t_SL g4294 ( 
.A(n_4101),
.Y(n_4294)
);

AND2x2_ASAP7_75t_L g4295 ( 
.A(n_4208),
.B(n_237),
.Y(n_4295)
);

INVxp67_ASAP7_75t_L g4296 ( 
.A(n_4152),
.Y(n_4296)
);

HB1xp67_ASAP7_75t_L g4297 ( 
.A(n_4232),
.Y(n_4297)
);

AND2x2_ASAP7_75t_L g4298 ( 
.A(n_4209),
.B(n_237),
.Y(n_4298)
);

INVx2_ASAP7_75t_L g4299 ( 
.A(n_4196),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_L g4300 ( 
.A(n_4108),
.B(n_4212),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4234),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_4220),
.B(n_238),
.Y(n_4302)
);

AND2x2_ASAP7_75t_L g4303 ( 
.A(n_4217),
.B(n_238),
.Y(n_4303)
);

HB1xp67_ASAP7_75t_L g4304 ( 
.A(n_4237),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4245),
.Y(n_4305)
);

AND2x2_ASAP7_75t_L g4306 ( 
.A(n_4225),
.B(n_239),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4247),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_4241),
.B(n_239),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_4242),
.B(n_240),
.Y(n_4309)
);

AND2x2_ASAP7_75t_L g4310 ( 
.A(n_4097),
.B(n_240),
.Y(n_4310)
);

INVx2_ASAP7_75t_L g4311 ( 
.A(n_4134),
.Y(n_4311)
);

AND2x2_ASAP7_75t_L g4312 ( 
.A(n_4219),
.B(n_4235),
.Y(n_4312)
);

OR2x2_ASAP7_75t_L g4313 ( 
.A(n_4248),
.B(n_241),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_4153),
.B(n_241),
.Y(n_4314)
);

AND2x2_ASAP7_75t_L g4315 ( 
.A(n_4149),
.B(n_4124),
.Y(n_4315)
);

INVx2_ASAP7_75t_L g4316 ( 
.A(n_4110),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_4154),
.B(n_242),
.Y(n_4317)
);

AND2x2_ASAP7_75t_L g4318 ( 
.A(n_4133),
.B(n_243),
.Y(n_4318)
);

AND2x2_ASAP7_75t_L g4319 ( 
.A(n_4132),
.B(n_244),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_L g4320 ( 
.A(n_4137),
.B(n_245),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4115),
.Y(n_4321)
);

AOI22xp33_ASAP7_75t_L g4322 ( 
.A1(n_4201),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_4322)
);

HB1xp67_ASAP7_75t_L g4323 ( 
.A(n_4094),
.Y(n_4323)
);

AND2x4_ASAP7_75t_L g4324 ( 
.A(n_4142),
.B(n_248),
.Y(n_4324)
);

OR2x2_ASAP7_75t_L g4325 ( 
.A(n_4113),
.B(n_4106),
.Y(n_4325)
);

NOR2xp67_ASAP7_75t_L g4326 ( 
.A(n_4177),
.B(n_250),
.Y(n_4326)
);

AOI22xp5_ASAP7_75t_L g4327 ( 
.A1(n_4138),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4203),
.Y(n_4328)
);

HB1xp67_ASAP7_75t_L g4329 ( 
.A(n_4210),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_4221),
.B(n_251),
.Y(n_4330)
);

OR2x2_ASAP7_75t_L g4331 ( 
.A(n_4093),
.B(n_252),
.Y(n_4331)
);

BUFx3_ASAP7_75t_L g4332 ( 
.A(n_4213),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4135),
.Y(n_4333)
);

AND2x2_ASAP7_75t_L g4334 ( 
.A(n_4127),
.B(n_255),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4168),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_L g4336 ( 
.A(n_4146),
.B(n_256),
.Y(n_4336)
);

INVx2_ASAP7_75t_L g4337 ( 
.A(n_4135),
.Y(n_4337)
);

OR2x2_ASAP7_75t_L g4338 ( 
.A(n_4105),
.B(n_257),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4169),
.Y(n_4339)
);

BUFx2_ASAP7_75t_L g4340 ( 
.A(n_4129),
.Y(n_4340)
);

AND2x2_ASAP7_75t_L g4341 ( 
.A(n_4112),
.B(n_257),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_SL g4342 ( 
.A(n_4157),
.B(n_258),
.Y(n_4342)
);

INVx2_ASAP7_75t_L g4343 ( 
.A(n_4243),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_4120),
.B(n_258),
.Y(n_4344)
);

AND2x4_ASAP7_75t_L g4345 ( 
.A(n_4096),
.B(n_259),
.Y(n_4345)
);

INVxp67_ASAP7_75t_L g4346 ( 
.A(n_4180),
.Y(n_4346)
);

OR2x2_ASAP7_75t_L g4347 ( 
.A(n_4114),
.B(n_259),
.Y(n_4347)
);

NAND2x1_ASAP7_75t_L g4348 ( 
.A(n_4098),
.B(n_261),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4128),
.Y(n_4349)
);

INVx2_ASAP7_75t_L g4350 ( 
.A(n_4123),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_4121),
.B(n_260),
.Y(n_4351)
);

HB1xp67_ASAP7_75t_L g4352 ( 
.A(n_4117),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_4103),
.B(n_260),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4125),
.Y(n_4354)
);

NOR2x1_ASAP7_75t_L g4355 ( 
.A(n_4233),
.B(n_261),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_L g4356 ( 
.A(n_4165),
.B(n_262),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4174),
.Y(n_4357)
);

AND2x2_ASAP7_75t_L g4358 ( 
.A(n_4179),
.B(n_262),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_4143),
.B(n_4111),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4162),
.Y(n_4360)
);

INVx2_ASAP7_75t_L g4361 ( 
.A(n_4186),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_L g4362 ( 
.A(n_4155),
.B(n_263),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4131),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4130),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_4238),
.B(n_263),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4145),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_4163),
.B(n_264),
.Y(n_4367)
);

OR2x2_ASAP7_75t_L g4368 ( 
.A(n_4148),
.B(n_4151),
.Y(n_4368)
);

INVx2_ASAP7_75t_L g4369 ( 
.A(n_4198),
.Y(n_4369)
);

AND2x2_ASAP7_75t_L g4370 ( 
.A(n_4099),
.B(n_264),
.Y(n_4370)
);

INVx2_ASAP7_75t_L g4371 ( 
.A(n_4150),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4171),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4182),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_4240),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_L g4375 ( 
.A(n_4200),
.B(n_265),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_4161),
.B(n_266),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4184),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4192),
.Y(n_4378)
);

AND2x4_ASAP7_75t_L g4379 ( 
.A(n_4226),
.B(n_267),
.Y(n_4379)
);

AND2x2_ASAP7_75t_L g4380 ( 
.A(n_4136),
.B(n_4139),
.Y(n_4380)
);

AND2x2_ASAP7_75t_L g4381 ( 
.A(n_4140),
.B(n_268),
.Y(n_4381)
);

AND2x2_ASAP7_75t_L g4382 ( 
.A(n_4164),
.B(n_268),
.Y(n_4382)
);

NAND2xp5_ASAP7_75t_L g4383 ( 
.A(n_4167),
.B(n_4173),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_4188),
.Y(n_4384)
);

INVx4_ASAP7_75t_L g4385 ( 
.A(n_4170),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4193),
.Y(n_4386)
);

AND2x2_ASAP7_75t_L g4387 ( 
.A(n_4189),
.B(n_269),
.Y(n_4387)
);

HB1xp67_ASAP7_75t_L g4388 ( 
.A(n_4175),
.Y(n_4388)
);

AND2x2_ASAP7_75t_SL g4389 ( 
.A(n_4191),
.B(n_269),
.Y(n_4389)
);

INVx2_ASAP7_75t_SL g4390 ( 
.A(n_4176),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4158),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_L g4392 ( 
.A(n_4199),
.B(n_270),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4178),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4160),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4183),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4187),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4172),
.Y(n_4397)
);

OR2x6_ASAP7_75t_L g4398 ( 
.A(n_4197),
.B(n_270),
.Y(n_4398)
);

AND2x2_ASAP7_75t_L g4399 ( 
.A(n_4156),
.B(n_272),
.Y(n_4399)
);

AND2x2_ASAP7_75t_L g4400 ( 
.A(n_4091),
.B(n_272),
.Y(n_4400)
);

AND2x4_ASAP7_75t_SL g4401 ( 
.A(n_4205),
.B(n_273),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_L g4402 ( 
.A(n_4095),
.B(n_273),
.Y(n_4402)
);

INVx4_ASAP7_75t_L g4403 ( 
.A(n_4118),
.Y(n_4403)
);

NOR2xp67_ASAP7_75t_L g4404 ( 
.A(n_4205),
.B(n_274),
.Y(n_4404)
);

AOI22xp33_ASAP7_75t_SL g4405 ( 
.A1(n_4147),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_4405)
);

HB1xp67_ASAP7_75t_L g4406 ( 
.A(n_4166),
.Y(n_4406)
);

AND2x2_ASAP7_75t_L g4407 ( 
.A(n_4091),
.B(n_278),
.Y(n_4407)
);

OR2x2_ASAP7_75t_L g4408 ( 
.A(n_4126),
.B(n_278),
.Y(n_4408)
);

INVx2_ASAP7_75t_L g4409 ( 
.A(n_4194),
.Y(n_4409)
);

AND2x2_ASAP7_75t_L g4410 ( 
.A(n_4091),
.B(n_279),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_4194),
.Y(n_4411)
);

AND2x2_ASAP7_75t_L g4412 ( 
.A(n_4091),
.B(n_280),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4107),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4091),
.B(n_280),
.Y(n_4414)
);

AND2x4_ASAP7_75t_L g4415 ( 
.A(n_4211),
.B(n_281),
.Y(n_4415)
);

NAND3xp33_ASAP7_75t_L g4416 ( 
.A(n_4233),
.B(n_281),
.C(n_282),
.Y(n_4416)
);

INVx1_ASAP7_75t_SL g4417 ( 
.A(n_4216),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_4194),
.Y(n_4418)
);

BUFx2_ASAP7_75t_L g4419 ( 
.A(n_4223),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4107),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4107),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_4107),
.Y(n_4422)
);

NAND2xp5_ASAP7_75t_L g4423 ( 
.A(n_4095),
.B(n_283),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4107),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4107),
.Y(n_4425)
);

INVx1_ASAP7_75t_L g4426 ( 
.A(n_4107),
.Y(n_4426)
);

HB1xp67_ASAP7_75t_L g4427 ( 
.A(n_4166),
.Y(n_4427)
);

AND2x2_ASAP7_75t_L g4428 ( 
.A(n_4091),
.B(n_283),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_4095),
.B(n_284),
.Y(n_4429)
);

HB1xp67_ASAP7_75t_L g4430 ( 
.A(n_4166),
.Y(n_4430)
);

OR2x2_ASAP7_75t_L g4431 ( 
.A(n_4126),
.B(n_285),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4091),
.B(n_285),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4107),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4095),
.B(n_286),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4107),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_4095),
.B(n_286),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4091),
.B(n_287),
.Y(n_4437)
);

BUFx2_ASAP7_75t_L g4438 ( 
.A(n_4223),
.Y(n_4438)
);

HB1xp67_ASAP7_75t_L g4439 ( 
.A(n_4166),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4107),
.Y(n_4440)
);

INVx2_ASAP7_75t_L g4441 ( 
.A(n_4194),
.Y(n_4441)
);

OR2x2_ASAP7_75t_L g4442 ( 
.A(n_4126),
.B(n_288),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_4194),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_4254),
.B(n_4323),
.Y(n_4444)
);

AND2x2_ASAP7_75t_L g4445 ( 
.A(n_4419),
.B(n_288),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4263),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_4329),
.B(n_289),
.Y(n_4447)
);

OR2x2_ASAP7_75t_L g4448 ( 
.A(n_4357),
.B(n_289),
.Y(n_4448)
);

INVx2_ASAP7_75t_L g4449 ( 
.A(n_4438),
.Y(n_4449)
);

AND2x2_ASAP7_75t_L g4450 ( 
.A(n_4292),
.B(n_290),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4297),
.Y(n_4451)
);

INVx3_ASAP7_75t_L g4452 ( 
.A(n_4403),
.Y(n_4452)
);

INVx2_ASAP7_75t_L g4453 ( 
.A(n_4281),
.Y(n_4453)
);

INVxp67_ASAP7_75t_L g4454 ( 
.A(n_4280),
.Y(n_4454)
);

AND2x2_ASAP7_75t_L g4455 ( 
.A(n_4283),
.B(n_290),
.Y(n_4455)
);

AND2x4_ASAP7_75t_L g4456 ( 
.A(n_4332),
.B(n_291),
.Y(n_4456)
);

OR2x2_ASAP7_75t_L g4457 ( 
.A(n_4372),
.B(n_291),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_4294),
.B(n_292),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_4391),
.B(n_292),
.Y(n_4459)
);

AND2x2_ASAP7_75t_L g4460 ( 
.A(n_4417),
.B(n_293),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4304),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_4258),
.Y(n_4462)
);

AND2x2_ASAP7_75t_L g4463 ( 
.A(n_4340),
.B(n_294),
.Y(n_4463)
);

HB1xp67_ASAP7_75t_L g4464 ( 
.A(n_4346),
.Y(n_4464)
);

AND2x2_ASAP7_75t_L g4465 ( 
.A(n_4380),
.B(n_294),
.Y(n_4465)
);

NAND4xp25_ASAP7_75t_L g4466 ( 
.A(n_4312),
.B(n_297),
.C(n_295),
.D(n_296),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4352),
.B(n_296),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4264),
.Y(n_4468)
);

AND2x2_ASAP7_75t_L g4469 ( 
.A(n_4270),
.B(n_298),
.Y(n_4469)
);

AND2x2_ASAP7_75t_L g4470 ( 
.A(n_4296),
.B(n_299),
.Y(n_4470)
);

AND2x4_ASAP7_75t_SL g4471 ( 
.A(n_4369),
.B(n_300),
.Y(n_4471)
);

AND2x4_ASAP7_75t_L g4472 ( 
.A(n_4299),
.B(n_300),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_L g4473 ( 
.A(n_4406),
.B(n_302),
.Y(n_4473)
);

OR2x2_ASAP7_75t_L g4474 ( 
.A(n_4328),
.B(n_303),
.Y(n_4474)
);

OR2x2_ASAP7_75t_L g4475 ( 
.A(n_4427),
.B(n_303),
.Y(n_4475)
);

AND2x4_ASAP7_75t_L g4476 ( 
.A(n_4271),
.B(n_304),
.Y(n_4476)
);

INVxp33_ASAP7_75t_L g4477 ( 
.A(n_4273),
.Y(n_4477)
);

AOI22xp5_ASAP7_75t_L g4478 ( 
.A1(n_4383),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.Y(n_4478)
);

HB1xp67_ASAP7_75t_L g4479 ( 
.A(n_4388),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_4430),
.B(n_305),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4269),
.Y(n_4481)
);

OR2x2_ASAP7_75t_L g4482 ( 
.A(n_4439),
.B(n_307),
.Y(n_4482)
);

OAI22xp5_ASAP7_75t_L g4483 ( 
.A1(n_4300),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_4483)
);

AND2x4_ASAP7_75t_L g4484 ( 
.A(n_4409),
.B(n_308),
.Y(n_4484)
);

OAI21xp33_ASAP7_75t_L g4485 ( 
.A1(n_4443),
.A2(n_309),
.B(n_311),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4321),
.Y(n_4486)
);

AND2x2_ASAP7_75t_L g4487 ( 
.A(n_4377),
.B(n_4378),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4384),
.B(n_312),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4386),
.B(n_312),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4268),
.B(n_313),
.Y(n_4490)
);

AND2x2_ASAP7_75t_L g4491 ( 
.A(n_4268),
.B(n_313),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_4397),
.B(n_314),
.Y(n_4492)
);

HB1xp67_ASAP7_75t_L g4493 ( 
.A(n_4411),
.Y(n_4493)
);

NOR2xp33_ASAP7_75t_L g4494 ( 
.A(n_4268),
.B(n_315),
.Y(n_4494)
);

INVx2_ASAP7_75t_L g4495 ( 
.A(n_4385),
.Y(n_4495)
);

AND2x2_ASAP7_75t_L g4496 ( 
.A(n_4315),
.B(n_315),
.Y(n_4496)
);

AND2x2_ASAP7_75t_L g4497 ( 
.A(n_4310),
.B(n_4252),
.Y(n_4497)
);

AND2x2_ASAP7_75t_L g4498 ( 
.A(n_4267),
.B(n_316),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_4394),
.B(n_316),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_4253),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4415),
.B(n_317),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4413),
.Y(n_4502)
);

NOR2xp33_ASAP7_75t_L g4503 ( 
.A(n_4348),
.B(n_317),
.Y(n_4503)
);

AND2x2_ASAP7_75t_L g4504 ( 
.A(n_4285),
.B(n_319),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4360),
.B(n_320),
.Y(n_4505)
);

AND2x2_ASAP7_75t_L g4506 ( 
.A(n_4319),
.B(n_320),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_L g4507 ( 
.A(n_4390),
.B(n_321),
.Y(n_4507)
);

AND2x2_ASAP7_75t_L g4508 ( 
.A(n_4374),
.B(n_322),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4420),
.Y(n_4509)
);

INVx3_ASAP7_75t_R g4510 ( 
.A(n_4345),
.Y(n_4510)
);

AOI22xp33_ASAP7_75t_L g4511 ( 
.A1(n_4275),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_4511)
);

AND2x2_ASAP7_75t_L g4512 ( 
.A(n_4334),
.B(n_325),
.Y(n_4512)
);

HB1xp67_ASAP7_75t_L g4513 ( 
.A(n_4418),
.Y(n_4513)
);

AND2x2_ASAP7_75t_L g4514 ( 
.A(n_4318),
.B(n_326),
.Y(n_4514)
);

AND3x2_ASAP7_75t_L g4515 ( 
.A(n_4343),
.B(n_326),
.C(n_327),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4421),
.Y(n_4516)
);

HB1xp67_ASAP7_75t_L g4517 ( 
.A(n_4441),
.Y(n_4517)
);

HB1xp67_ASAP7_75t_L g4518 ( 
.A(n_4364),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4422),
.Y(n_4519)
);

HB1xp67_ASAP7_75t_L g4520 ( 
.A(n_4366),
.Y(n_4520)
);

INVx1_ASAP7_75t_SL g4521 ( 
.A(n_4389),
.Y(n_4521)
);

AND2x2_ASAP7_75t_L g4522 ( 
.A(n_4257),
.B(n_327),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_L g4523 ( 
.A(n_4395),
.B(n_329),
.Y(n_4523)
);

NAND2xp5_ASAP7_75t_L g4524 ( 
.A(n_4396),
.B(n_331),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_L g4525 ( 
.A(n_4349),
.B(n_331),
.Y(n_4525)
);

INVx2_ASAP7_75t_L g4526 ( 
.A(n_4333),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4337),
.Y(n_4527)
);

HB1xp67_ASAP7_75t_L g4528 ( 
.A(n_4368),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4424),
.Y(n_4529)
);

AND2x2_ASAP7_75t_L g4530 ( 
.A(n_4425),
.B(n_332),
.Y(n_4530)
);

INVx3_ASAP7_75t_L g4531 ( 
.A(n_4277),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_4426),
.Y(n_4532)
);

INVx1_ASAP7_75t_L g4533 ( 
.A(n_4433),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4435),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_4440),
.B(n_333),
.Y(n_4535)
);

INVx1_ASAP7_75t_SL g4536 ( 
.A(n_4401),
.Y(n_4536)
);

AND2x2_ASAP7_75t_L g4537 ( 
.A(n_4336),
.B(n_4272),
.Y(n_4537)
);

INVx2_ASAP7_75t_L g4538 ( 
.A(n_4361),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4276),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4282),
.B(n_334),
.Y(n_4540)
);

OR2x2_ASAP7_75t_L g4541 ( 
.A(n_4363),
.B(n_334),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_SL g4542 ( 
.A(n_4325),
.B(n_4359),
.Y(n_4542)
);

AND2x2_ASAP7_75t_L g4543 ( 
.A(n_4289),
.B(n_335),
.Y(n_4543)
);

NAND2xp5_ASAP7_75t_L g4544 ( 
.A(n_4288),
.B(n_335),
.Y(n_4544)
);

AND2x4_ASAP7_75t_L g4545 ( 
.A(n_4371),
.B(n_336),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4290),
.B(n_339),
.Y(n_4546)
);

NOR2xp67_ASAP7_75t_L g4547 ( 
.A(n_4404),
.B(n_339),
.Y(n_4547)
);

AND2x2_ASAP7_75t_L g4548 ( 
.A(n_4291),
.B(n_340),
.Y(n_4548)
);

BUFx2_ASAP7_75t_SL g4549 ( 
.A(n_4326),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4293),
.Y(n_4550)
);

NAND2x1_ASAP7_75t_L g4551 ( 
.A(n_4301),
.B(n_341),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_4320),
.B(n_341),
.Y(n_4552)
);

INVx2_ASAP7_75t_L g4553 ( 
.A(n_4331),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_4305),
.Y(n_4554)
);

AND2x2_ASAP7_75t_L g4555 ( 
.A(n_4307),
.B(n_342),
.Y(n_4555)
);

NOR2xp33_ASAP7_75t_L g4556 ( 
.A(n_4408),
.B(n_342),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_4274),
.Y(n_4557)
);

AND2x4_ASAP7_75t_L g4558 ( 
.A(n_4358),
.B(n_343),
.Y(n_4558)
);

INVx2_ASAP7_75t_L g4559 ( 
.A(n_4338),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4278),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_4313),
.Y(n_4561)
);

AND2x4_ASAP7_75t_L g4562 ( 
.A(n_4250),
.B(n_344),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4284),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4335),
.Y(n_4564)
);

INVx2_ASAP7_75t_L g4565 ( 
.A(n_4393),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4339),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4431),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4442),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4347),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4314),
.Y(n_4570)
);

OR2x2_ASAP7_75t_L g4571 ( 
.A(n_4262),
.B(n_344),
.Y(n_4571)
);

HB1xp67_ASAP7_75t_L g4572 ( 
.A(n_4375),
.Y(n_4572)
);

INVx2_ASAP7_75t_SL g4573 ( 
.A(n_4382),
.Y(n_4573)
);

OR2x2_ASAP7_75t_L g4574 ( 
.A(n_4317),
.B(n_345),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4311),
.Y(n_4575)
);

BUFx2_ASAP7_75t_L g4576 ( 
.A(n_4387),
.Y(n_4576)
);

OR2x2_ASAP7_75t_L g4577 ( 
.A(n_4260),
.B(n_346),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4367),
.Y(n_4578)
);

AND2x4_ASAP7_75t_L g4579 ( 
.A(n_4255),
.B(n_347),
.Y(n_4579)
);

INVx2_ASAP7_75t_L g4580 ( 
.A(n_4350),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4316),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_4576),
.B(n_4261),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4528),
.Y(n_4583)
);

INVx3_ASAP7_75t_L g4584 ( 
.A(n_4452),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4479),
.Y(n_4585)
);

INVx2_ASAP7_75t_L g4586 ( 
.A(n_4497),
.Y(n_4586)
);

AND2x2_ASAP7_75t_L g4587 ( 
.A(n_4453),
.B(n_4295),
.Y(n_4587)
);

NAND2xp33_ASAP7_75t_R g4588 ( 
.A(n_4515),
.B(n_4392),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4459),
.Y(n_4589)
);

OR2x2_ASAP7_75t_L g4590 ( 
.A(n_4444),
.B(n_4251),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4464),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4447),
.Y(n_4592)
);

AND2x2_ASAP7_75t_L g4593 ( 
.A(n_4536),
.B(n_4298),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4467),
.Y(n_4594)
);

INVx2_ASAP7_75t_L g4595 ( 
.A(n_4472),
.Y(n_4595)
);

AND2x2_ASAP7_75t_L g4596 ( 
.A(n_4454),
.B(n_4303),
.Y(n_4596)
);

INVx2_ASAP7_75t_L g4597 ( 
.A(n_4450),
.Y(n_4597)
);

OR2x2_ASAP7_75t_L g4598 ( 
.A(n_4449),
.B(n_4402),
.Y(n_4598)
);

INVx3_ASAP7_75t_L g4599 ( 
.A(n_4456),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4518),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4520),
.Y(n_4601)
);

AND2x4_ASAP7_75t_L g4602 ( 
.A(n_4531),
.B(n_4379),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4446),
.Y(n_4603)
);

INVx2_ASAP7_75t_L g4604 ( 
.A(n_4465),
.Y(n_4604)
);

NAND2xp5_ASAP7_75t_L g4605 ( 
.A(n_4573),
.B(n_4405),
.Y(n_4605)
);

INVx2_ASAP7_75t_L g4606 ( 
.A(n_4490),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4475),
.Y(n_4607)
);

OR2x2_ASAP7_75t_L g4608 ( 
.A(n_4542),
.B(n_4423),
.Y(n_4608)
);

INVx2_ASAP7_75t_SL g4609 ( 
.A(n_4471),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4482),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4552),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4569),
.Y(n_4612)
);

AND2x2_ASAP7_75t_L g4613 ( 
.A(n_4537),
.B(n_4306),
.Y(n_4613)
);

AND2x2_ASAP7_75t_L g4614 ( 
.A(n_4445),
.B(n_4309),
.Y(n_4614)
);

OAI31xp33_ASAP7_75t_L g4615 ( 
.A1(n_4521),
.A2(n_4477),
.A3(n_4416),
.B(n_4249),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4495),
.B(n_4381),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_4530),
.B(n_4342),
.Y(n_4617)
);

AND2x2_ASAP7_75t_L g4618 ( 
.A(n_4535),
.B(n_4370),
.Y(n_4618)
);

INVx2_ASAP7_75t_L g4619 ( 
.A(n_4491),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4473),
.Y(n_4620)
);

OR2x2_ASAP7_75t_L g4621 ( 
.A(n_4557),
.B(n_4429),
.Y(n_4621)
);

INVx4_ASAP7_75t_L g4622 ( 
.A(n_4469),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4493),
.B(n_4259),
.Y(n_4623)
);

INVx2_ASAP7_75t_L g4624 ( 
.A(n_4551),
.Y(n_4624)
);

NAND2x1_ASAP7_75t_L g4625 ( 
.A(n_4451),
.B(n_4373),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4480),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_4572),
.B(n_4355),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4513),
.B(n_4265),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4474),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4517),
.B(n_4266),
.Y(n_4630)
);

INVx2_ASAP7_75t_L g4631 ( 
.A(n_4496),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4522),
.B(n_4327),
.Y(n_4632)
);

NOR2x1_ASAP7_75t_L g4633 ( 
.A(n_4466),
.B(n_4434),
.Y(n_4633)
);

OR2x2_ASAP7_75t_L g4634 ( 
.A(n_4560),
.B(n_4436),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4461),
.Y(n_4635)
);

NOR2xp33_ASAP7_75t_L g4636 ( 
.A(n_4510),
.B(n_4362),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4505),
.B(n_4279),
.Y(n_4637)
);

AND2x2_ASAP7_75t_L g4638 ( 
.A(n_4463),
.B(n_4455),
.Y(n_4638)
);

INVx2_ASAP7_75t_L g4639 ( 
.A(n_4558),
.Y(n_4639)
);

AND2x2_ASAP7_75t_L g4640 ( 
.A(n_4487),
.B(n_4400),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4581),
.Y(n_4641)
);

AND2x2_ASAP7_75t_L g4642 ( 
.A(n_4460),
.B(n_4407),
.Y(n_4642)
);

AND2x2_ASAP7_75t_L g4643 ( 
.A(n_4470),
.B(n_4488),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_4564),
.Y(n_4644)
);

AND2x2_ASAP7_75t_L g4645 ( 
.A(n_4489),
.B(n_4410),
.Y(n_4645)
);

AND2x2_ASAP7_75t_L g4646 ( 
.A(n_4540),
.B(n_4412),
.Y(n_4646)
);

AND2x2_ASAP7_75t_L g4647 ( 
.A(n_4543),
.B(n_4414),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4566),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4457),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4561),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_4462),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_4546),
.B(n_4548),
.Y(n_4652)
);

OR2x2_ASAP7_75t_L g4653 ( 
.A(n_4570),
.B(n_4302),
.Y(n_4653)
);

AND2x4_ASAP7_75t_SL g4654 ( 
.A(n_4458),
.B(n_4351),
.Y(n_4654)
);

AND2x2_ASAP7_75t_L g4655 ( 
.A(n_4555),
.B(n_4428),
.Y(n_4655)
);

AND2x2_ASAP7_75t_L g4656 ( 
.A(n_4494),
.B(n_4500),
.Y(n_4656)
);

OR2x2_ASAP7_75t_L g4657 ( 
.A(n_4525),
.B(n_4578),
.Y(n_4657)
);

OR2x2_ASAP7_75t_L g4658 ( 
.A(n_4492),
.B(n_4308),
.Y(n_4658)
);

INVx1_ASAP7_75t_SL g4659 ( 
.A(n_4549),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_4468),
.Y(n_4660)
);

BUFx3_ASAP7_75t_L g4661 ( 
.A(n_4512),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4481),
.Y(n_4662)
);

AND2x2_ASAP7_75t_L g4663 ( 
.A(n_4502),
.B(n_4432),
.Y(n_4663)
);

INVx2_ASAP7_75t_L g4664 ( 
.A(n_4476),
.Y(n_4664)
);

AND2x2_ASAP7_75t_L g4665 ( 
.A(n_4509),
.B(n_4437),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_L g4666 ( 
.A(n_4567),
.B(n_4322),
.Y(n_4666)
);

INVx3_ASAP7_75t_L g4667 ( 
.A(n_4484),
.Y(n_4667)
);

INVxp67_ASAP7_75t_L g4668 ( 
.A(n_4547),
.Y(n_4668)
);

AND2x2_ASAP7_75t_SL g4669 ( 
.A(n_4568),
.B(n_4341),
.Y(n_4669)
);

HB1xp67_ASAP7_75t_L g4670 ( 
.A(n_4526),
.Y(n_4670)
);

AND2x2_ASAP7_75t_L g4671 ( 
.A(n_4516),
.B(n_4344),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_4539),
.Y(n_4672)
);

NAND2xp5_ASAP7_75t_L g4673 ( 
.A(n_4556),
.B(n_4356),
.Y(n_4673)
);

AND2x2_ASAP7_75t_L g4674 ( 
.A(n_4519),
.B(n_4256),
.Y(n_4674)
);

OR2x2_ASAP7_75t_L g4675 ( 
.A(n_4499),
.B(n_4330),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4613),
.B(n_4478),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4583),
.Y(n_4677)
);

AND2x2_ASAP7_75t_L g4678 ( 
.A(n_4593),
.B(n_4529),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4587),
.B(n_4532),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4621),
.Y(n_4680)
);

OR2x6_ASAP7_75t_L g4681 ( 
.A(n_4609),
.B(n_4507),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_L g4682 ( 
.A(n_4661),
.B(n_4541),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_4634),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4671),
.B(n_4448),
.Y(n_4684)
);

OR2x2_ASAP7_75t_L g4685 ( 
.A(n_4591),
.B(n_4533),
.Y(n_4685)
);

INVx2_ASAP7_75t_SL g4686 ( 
.A(n_4618),
.Y(n_4686)
);

AND2x2_ASAP7_75t_L g4687 ( 
.A(n_4596),
.B(n_4534),
.Y(n_4687)
);

OR2x2_ASAP7_75t_L g4688 ( 
.A(n_4582),
.B(n_4523),
.Y(n_4688)
);

NAND2xp5_ASAP7_75t_L g4689 ( 
.A(n_4597),
.B(n_4514),
.Y(n_4689)
);

INVx2_ASAP7_75t_L g4690 ( 
.A(n_4654),
.Y(n_4690)
);

INVx2_ASAP7_75t_L g4691 ( 
.A(n_4642),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4670),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_4604),
.B(n_4504),
.Y(n_4693)
);

INVx2_ASAP7_75t_L g4694 ( 
.A(n_4614),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4653),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4585),
.Y(n_4696)
);

NAND2xp5_ASAP7_75t_L g4697 ( 
.A(n_4631),
.B(n_4527),
.Y(n_4697)
);

AND2x2_ASAP7_75t_L g4698 ( 
.A(n_4616),
.B(n_4550),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4600),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4601),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4589),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4657),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_L g4703 ( 
.A(n_4652),
.B(n_4565),
.Y(n_4703)
);

OR2x2_ASAP7_75t_L g4704 ( 
.A(n_4608),
.B(n_4524),
.Y(n_4704)
);

INVx1_ASAP7_75t_SL g4705 ( 
.A(n_4669),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4629),
.Y(n_4706)
);

INVxp67_ASAP7_75t_SL g4707 ( 
.A(n_4636),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_4640),
.B(n_4544),
.Y(n_4708)
);

INVxp67_ASAP7_75t_SL g4709 ( 
.A(n_4599),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4623),
.B(n_4628),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4649),
.Y(n_4711)
);

HB1xp67_ASAP7_75t_L g4712 ( 
.A(n_4630),
.Y(n_4712)
);

NAND2xp5_ASAP7_75t_L g4713 ( 
.A(n_4643),
.B(n_4663),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4607),
.Y(n_4714)
);

HB1xp67_ASAP7_75t_L g4715 ( 
.A(n_4625),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4610),
.Y(n_4716)
);

OR2x2_ASAP7_75t_L g4717 ( 
.A(n_4590),
.B(n_4554),
.Y(n_4717)
);

HB1xp67_ASAP7_75t_L g4718 ( 
.A(n_4638),
.Y(n_4718)
);

AND2x2_ASAP7_75t_L g4719 ( 
.A(n_4659),
.B(n_4508),
.Y(n_4719)
);

NAND2x1p5_ASAP7_75t_L g4720 ( 
.A(n_4584),
.B(n_4506),
.Y(n_4720)
);

OR2x2_ASAP7_75t_L g4721 ( 
.A(n_4598),
.B(n_4486),
.Y(n_4721)
);

OR2x2_ASAP7_75t_L g4722 ( 
.A(n_4586),
.B(n_4563),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_4611),
.Y(n_4723)
);

INVx2_ASAP7_75t_L g4724 ( 
.A(n_4645),
.Y(n_4724)
);

INVx2_ASAP7_75t_L g4725 ( 
.A(n_4646),
.Y(n_4725)
);

INVx1_ASAP7_75t_L g4726 ( 
.A(n_4650),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4665),
.B(n_4503),
.Y(n_4727)
);

AND2x2_ASAP7_75t_L g4728 ( 
.A(n_4602),
.B(n_4498),
.Y(n_4728)
);

OR2x2_ASAP7_75t_L g4729 ( 
.A(n_4612),
.B(n_4571),
.Y(n_4729)
);

AND2x2_ASAP7_75t_L g4730 ( 
.A(n_4674),
.B(n_4501),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4617),
.B(n_4574),
.Y(n_4731)
);

AND2x2_ASAP7_75t_L g4732 ( 
.A(n_4624),
.B(n_4545),
.Y(n_4732)
);

INVx1_ASAP7_75t_L g4733 ( 
.A(n_4594),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_4592),
.Y(n_4734)
);

NOR2xp33_ASAP7_75t_L g4735 ( 
.A(n_4622),
.B(n_4577),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_4712),
.Y(n_4736)
);

INVxp67_ASAP7_75t_SL g4737 ( 
.A(n_4718),
.Y(n_4737)
);

AND2x2_ASAP7_75t_L g4738 ( 
.A(n_4719),
.B(n_4656),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4713),
.Y(n_4739)
);

AND2x2_ASAP7_75t_L g4740 ( 
.A(n_4728),
.B(n_4647),
.Y(n_4740)
);

OAI22xp5_ASAP7_75t_L g4741 ( 
.A1(n_4705),
.A2(n_4720),
.B1(n_4707),
.B2(n_4710),
.Y(n_4741)
);

AND2x2_ASAP7_75t_L g4742 ( 
.A(n_4678),
.B(n_4655),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4729),
.Y(n_4743)
);

AND2x2_ASAP7_75t_L g4744 ( 
.A(n_4709),
.B(n_4603),
.Y(n_4744)
);

AND2x2_ASAP7_75t_L g4745 ( 
.A(n_4686),
.B(n_4635),
.Y(n_4745)
);

AND2x2_ASAP7_75t_L g4746 ( 
.A(n_4679),
.B(n_4633),
.Y(n_4746)
);

INVxp67_ASAP7_75t_L g4747 ( 
.A(n_4715),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4691),
.Y(n_4748)
);

INVx2_ASAP7_75t_L g4749 ( 
.A(n_4731),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4717),
.Y(n_4750)
);

INVx2_ASAP7_75t_L g4751 ( 
.A(n_4730),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4721),
.Y(n_4752)
);

NOR2x1_ASAP7_75t_L g4753 ( 
.A(n_4692),
.B(n_4605),
.Y(n_4753)
);

AND2x2_ASAP7_75t_L g4754 ( 
.A(n_4698),
.B(n_4667),
.Y(n_4754)
);

INVx2_ASAP7_75t_L g4755 ( 
.A(n_4724),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4725),
.Y(n_4756)
);

OR2x2_ASAP7_75t_L g4757 ( 
.A(n_4694),
.B(n_4627),
.Y(n_4757)
);

AND2x2_ASAP7_75t_L g4758 ( 
.A(n_4687),
.B(n_4644),
.Y(n_4758)
);

BUFx2_ASAP7_75t_L g4759 ( 
.A(n_4681),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4703),
.Y(n_4760)
);

AND2x2_ASAP7_75t_L g4761 ( 
.A(n_4690),
.B(n_4648),
.Y(n_4761)
);

INVx2_ASAP7_75t_L g4762 ( 
.A(n_4732),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4680),
.B(n_4606),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4704),
.Y(n_4764)
);

INVxp67_ASAP7_75t_L g4765 ( 
.A(n_4735),
.Y(n_4765)
);

OR2x2_ASAP7_75t_L g4766 ( 
.A(n_4683),
.B(n_4641),
.Y(n_4766)
);

OR2x2_ASAP7_75t_L g4767 ( 
.A(n_4702),
.B(n_4620),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4689),
.Y(n_4768)
);

OR2x2_ASAP7_75t_L g4769 ( 
.A(n_4695),
.B(n_4626),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_4693),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_L g4771 ( 
.A(n_4684),
.B(n_4619),
.Y(n_4771)
);

XNOR2x1_ASAP7_75t_L g4772 ( 
.A(n_4688),
.B(n_4658),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_L g4773 ( 
.A(n_4682),
.B(n_4639),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4681),
.B(n_4651),
.Y(n_4774)
);

NOR2x1_ASAP7_75t_L g4775 ( 
.A(n_4733),
.B(n_4483),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_4676),
.B(n_4673),
.Y(n_4776)
);

NAND2xp5_ASAP7_75t_L g4777 ( 
.A(n_4708),
.B(n_4637),
.Y(n_4777)
);

HB1xp67_ASAP7_75t_L g4778 ( 
.A(n_4727),
.Y(n_4778)
);

INVx2_ASAP7_75t_L g4779 ( 
.A(n_4722),
.Y(n_4779)
);

INVx2_ASAP7_75t_L g4780 ( 
.A(n_4685),
.Y(n_4780)
);

AND2x2_ASAP7_75t_L g4781 ( 
.A(n_4714),
.B(n_4660),
.Y(n_4781)
);

INVx1_ASAP7_75t_SL g4782 ( 
.A(n_4759),
.Y(n_4782)
);

NAND3xp33_ASAP7_75t_L g4783 ( 
.A(n_4753),
.B(n_4741),
.C(n_4747),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_L g4784 ( 
.A(n_4742),
.B(n_4664),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4737),
.Y(n_4785)
);

OAI21xp33_ASAP7_75t_SL g4786 ( 
.A1(n_4775),
.A2(n_4726),
.B(n_4716),
.Y(n_4786)
);

AOI22xp5_ASAP7_75t_L g4787 ( 
.A1(n_4746),
.A2(n_4588),
.B1(n_4668),
.B2(n_4632),
.Y(n_4787)
);

NAND2xp5_ASAP7_75t_L g4788 ( 
.A(n_4738),
.B(n_4615),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4772),
.Y(n_4789)
);

XOR2xp5_ASAP7_75t_L g4790 ( 
.A(n_4778),
.B(n_4562),
.Y(n_4790)
);

O2A1O1Ixp33_ASAP7_75t_L g4791 ( 
.A1(n_4780),
.A2(n_4696),
.B(n_4700),
.C(n_4699),
.Y(n_4791)
);

INVx2_ASAP7_75t_SL g4792 ( 
.A(n_4740),
.Y(n_4792)
);

AOI21xp5_ASAP7_75t_L g4793 ( 
.A1(n_4777),
.A2(n_4666),
.B(n_4776),
.Y(n_4793)
);

AOI21xp33_ASAP7_75t_L g4794 ( 
.A1(n_4771),
.A2(n_4697),
.B(n_4734),
.Y(n_4794)
);

AND2x2_ASAP7_75t_L g4795 ( 
.A(n_4754),
.B(n_4706),
.Y(n_4795)
);

XOR2x2_ASAP7_75t_L g4796 ( 
.A(n_4773),
.B(n_4675),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4749),
.Y(n_4797)
);

INVx2_ASAP7_75t_L g4798 ( 
.A(n_4751),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4758),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4744),
.Y(n_4800)
);

XNOR2x2_ASAP7_75t_L g4801 ( 
.A(n_4774),
.B(n_4677),
.Y(n_4801)
);

XOR2x2_ASAP7_75t_L g4802 ( 
.A(n_4764),
.B(n_4579),
.Y(n_4802)
);

AOI22xp33_ASAP7_75t_L g4803 ( 
.A1(n_4779),
.A2(n_4538),
.B1(n_4559),
.B2(n_4553),
.Y(n_4803)
);

OAI221xp5_ASAP7_75t_L g4804 ( 
.A1(n_4763),
.A2(n_4711),
.B1(n_4575),
.B2(n_4485),
.C(n_4723),
.Y(n_4804)
);

OAI211xp5_ASAP7_75t_L g4805 ( 
.A1(n_4736),
.A2(n_4701),
.B(n_4672),
.C(n_4662),
.Y(n_4805)
);

XNOR2x2_ASAP7_75t_L g4806 ( 
.A(n_4767),
.B(n_4353),
.Y(n_4806)
);

AND2x2_ASAP7_75t_L g4807 ( 
.A(n_4745),
.B(n_4761),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4750),
.Y(n_4808)
);

AOI211xp5_ASAP7_75t_L g4809 ( 
.A1(n_4743),
.A2(n_4365),
.B(n_4580),
.C(n_4376),
.Y(n_4809)
);

AND2x2_ASAP7_75t_L g4810 ( 
.A(n_4755),
.B(n_4595),
.Y(n_4810)
);

NAND2xp5_ASAP7_75t_L g4811 ( 
.A(n_4762),
.B(n_4286),
.Y(n_4811)
);

O2A1O1Ixp33_ASAP7_75t_L g4812 ( 
.A1(n_4752),
.A2(n_4398),
.B(n_4287),
.C(n_4399),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4769),
.Y(n_4813)
);

OAI22xp5_ASAP7_75t_L g4814 ( 
.A1(n_4765),
.A2(n_4511),
.B1(n_4324),
.B2(n_4354),
.Y(n_4814)
);

AOI22xp5_ASAP7_75t_L g4815 ( 
.A1(n_4760),
.A2(n_4398),
.B1(n_350),
.B2(n_348),
.Y(n_4815)
);

OAI21xp33_ASAP7_75t_L g4816 ( 
.A1(n_4739),
.A2(n_349),
.B(n_350),
.Y(n_4816)
);

O2A1O1Ixp33_ASAP7_75t_L g4817 ( 
.A1(n_4766),
.A2(n_352),
.B(n_349),
.C(n_351),
.Y(n_4817)
);

OAI21xp5_ASAP7_75t_L g4818 ( 
.A1(n_4748),
.A2(n_351),
.B(n_353),
.Y(n_4818)
);

OAI21xp33_ASAP7_75t_L g4819 ( 
.A1(n_4756),
.A2(n_353),
.B(n_354),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4781),
.Y(n_4820)
);

AOI21xp5_ASAP7_75t_L g4821 ( 
.A1(n_4757),
.A2(n_354),
.B(n_355),
.Y(n_4821)
);

HB1xp67_ASAP7_75t_L g4822 ( 
.A(n_4768),
.Y(n_4822)
);

AOI22xp33_ASAP7_75t_L g4823 ( 
.A1(n_4770),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_4737),
.Y(n_4824)
);

OAI21xp33_ASAP7_75t_L g4825 ( 
.A1(n_4753),
.A2(n_358),
.B(n_359),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4737),
.Y(n_4826)
);

XOR2x2_ASAP7_75t_L g4827 ( 
.A(n_4772),
.B(n_358),
.Y(n_4827)
);

AND2x2_ASAP7_75t_L g4828 ( 
.A(n_4807),
.B(n_359),
.Y(n_4828)
);

AOI332xp33_ASAP7_75t_L g4829 ( 
.A1(n_4785),
.A2(n_365),
.A3(n_364),
.B1(n_362),
.B2(n_366),
.B3(n_360),
.C1(n_361),
.C2(n_363),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4796),
.Y(n_4830)
);

OAI33xp33_ASAP7_75t_L g4831 ( 
.A1(n_4783),
.A2(n_362),
.A3(n_367),
.B1(n_360),
.B2(n_361),
.B3(n_364),
.Y(n_4831)
);

INVxp67_ASAP7_75t_L g4832 ( 
.A(n_4790),
.Y(n_4832)
);

AOI222xp33_ASAP7_75t_L g4833 ( 
.A1(n_4786),
.A2(n_369),
.B1(n_371),
.B2(n_367),
.C1(n_368),
.C2(n_370),
.Y(n_4833)
);

NAND2xp5_ASAP7_75t_L g4834 ( 
.A(n_4792),
.B(n_368),
.Y(n_4834)
);

AOI221xp5_ASAP7_75t_L g4835 ( 
.A1(n_4825),
.A2(n_387),
.B1(n_397),
.B2(n_378),
.C(n_370),
.Y(n_4835)
);

OAI321xp33_ASAP7_75t_L g4836 ( 
.A1(n_4787),
.A2(n_373),
.A3(n_375),
.B1(n_371),
.B2(n_372),
.C(n_374),
.Y(n_4836)
);

NAND3xp33_ASAP7_75t_SL g4837 ( 
.A(n_4782),
.B(n_373),
.C(n_374),
.Y(n_4837)
);

OR2x2_ASAP7_75t_L g4838 ( 
.A(n_4788),
.B(n_375),
.Y(n_4838)
);

OAI221xp5_ASAP7_75t_L g4839 ( 
.A1(n_4789),
.A2(n_379),
.B1(n_376),
.B2(n_377),
.C(n_381),
.Y(n_4839)
);

INVx2_ASAP7_75t_L g4840 ( 
.A(n_4802),
.Y(n_4840)
);

INVxp33_ASAP7_75t_L g4841 ( 
.A(n_4827),
.Y(n_4841)
);

INVxp67_ASAP7_75t_L g4842 ( 
.A(n_4806),
.Y(n_4842)
);

AND2x2_ASAP7_75t_L g4843 ( 
.A(n_4795),
.B(n_376),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4810),
.Y(n_4844)
);

AOI22xp5_ASAP7_75t_L g4845 ( 
.A1(n_4811),
.A2(n_389),
.B1(n_399),
.B2(n_377),
.Y(n_4845)
);

AND2x2_ASAP7_75t_L g4846 ( 
.A(n_4798),
.B(n_379),
.Y(n_4846)
);

INVx2_ASAP7_75t_L g4847 ( 
.A(n_4801),
.Y(n_4847)
);

AOI22xp5_ASAP7_75t_L g4848 ( 
.A1(n_4793),
.A2(n_392),
.B1(n_401),
.B2(n_381),
.Y(n_4848)
);

OAI22xp33_ASAP7_75t_L g4849 ( 
.A1(n_4815),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_4849)
);

AND2x2_ASAP7_75t_L g4850 ( 
.A(n_4799),
.B(n_382),
.Y(n_4850)
);

AOI211xp5_ASAP7_75t_L g4851 ( 
.A1(n_4794),
.A2(n_385),
.B(n_383),
.C(n_384),
.Y(n_4851)
);

NAND2xp5_ASAP7_75t_L g4852 ( 
.A(n_4820),
.B(n_385),
.Y(n_4852)
);

OAI21xp5_ASAP7_75t_L g4853 ( 
.A1(n_4784),
.A2(n_386),
.B(n_389),
.Y(n_4853)
);

INVx2_ASAP7_75t_L g4854 ( 
.A(n_4813),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4822),
.Y(n_4855)
);

AOI21xp5_ASAP7_75t_L g4856 ( 
.A1(n_4791),
.A2(n_394),
.B(n_393),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_L g4857 ( 
.A(n_4800),
.B(n_390),
.Y(n_4857)
);

NOR2xp33_ASAP7_75t_L g4858 ( 
.A(n_4824),
.B(n_394),
.Y(n_4858)
);

OAI22xp5_ASAP7_75t_L g4859 ( 
.A1(n_4797),
.A2(n_398),
.B1(n_395),
.B2(n_396),
.Y(n_4859)
);

AOI21xp33_ASAP7_75t_SL g4860 ( 
.A1(n_4826),
.A2(n_396),
.B(n_398),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4817),
.Y(n_4861)
);

OAI33xp33_ASAP7_75t_L g4862 ( 
.A1(n_4808),
.A2(n_402),
.A3(n_404),
.B1(n_399),
.B2(n_400),
.B3(n_403),
.Y(n_4862)
);

NAND2xp5_ASAP7_75t_L g4863 ( 
.A(n_4821),
.B(n_402),
.Y(n_4863)
);

INVxp67_ASAP7_75t_L g4864 ( 
.A(n_4804),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4816),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4819),
.Y(n_4866)
);

INVx2_ASAP7_75t_SL g4867 ( 
.A(n_4814),
.Y(n_4867)
);

AOI21xp5_ASAP7_75t_L g4868 ( 
.A1(n_4805),
.A2(n_407),
.B(n_406),
.Y(n_4868)
);

NAND4xp25_ASAP7_75t_L g4869 ( 
.A(n_4809),
.B(n_408),
.C(n_405),
.D(n_406),
.Y(n_4869)
);

OAI32xp33_ASAP7_75t_L g4870 ( 
.A1(n_4818),
.A2(n_409),
.A3(n_405),
.B1(n_408),
.B2(n_410),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4823),
.B(n_409),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4812),
.Y(n_4872)
);

INVx3_ASAP7_75t_L g4873 ( 
.A(n_4803),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4796),
.Y(n_4874)
);

XNOR2x1_ASAP7_75t_L g4875 ( 
.A(n_4827),
.B(n_410),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4796),
.Y(n_4876)
);

NAND4xp25_ASAP7_75t_SL g4877 ( 
.A(n_4786),
.B(n_414),
.C(n_411),
.D(n_413),
.Y(n_4877)
);

INVxp67_ASAP7_75t_L g4878 ( 
.A(n_4807),
.Y(n_4878)
);

AOI321xp33_ASAP7_75t_L g4879 ( 
.A1(n_4789),
.A2(n_415),
.A3(n_417),
.B1(n_413),
.B2(n_414),
.C(n_416),
.Y(n_4879)
);

AOI31xp33_ASAP7_75t_L g4880 ( 
.A1(n_4783),
.A2(n_417),
.A3(n_415),
.B(n_416),
.Y(n_4880)
);

OAI211xp5_ASAP7_75t_L g4881 ( 
.A1(n_4786),
.A2(n_420),
.B(n_418),
.C(n_419),
.Y(n_4881)
);

INVx2_ASAP7_75t_L g4882 ( 
.A(n_4828),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4843),
.Y(n_4883)
);

HB1xp67_ASAP7_75t_L g4884 ( 
.A(n_4847),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4838),
.Y(n_4885)
);

AND2x4_ASAP7_75t_L g4886 ( 
.A(n_4878),
.B(n_418),
.Y(n_4886)
);

OAI21xp33_ASAP7_75t_SL g4887 ( 
.A1(n_4877),
.A2(n_420),
.B(n_421),
.Y(n_4887)
);

OAI21xp5_ASAP7_75t_L g4888 ( 
.A1(n_4842),
.A2(n_421),
.B(n_422),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4844),
.Y(n_4889)
);

INVx2_ASAP7_75t_L g4890 ( 
.A(n_4875),
.Y(n_4890)
);

AOI32xp33_ASAP7_75t_L g4891 ( 
.A1(n_4830),
.A2(n_424),
.A3(n_422),
.B1(n_423),
.B2(n_425),
.Y(n_4891)
);

AND2x2_ASAP7_75t_L g4892 ( 
.A(n_4854),
.B(n_424),
.Y(n_4892)
);

INVx2_ASAP7_75t_L g4893 ( 
.A(n_4850),
.Y(n_4893)
);

A2O1A1Ixp33_ASAP7_75t_L g4894 ( 
.A1(n_4856),
.A2(n_428),
.B(n_426),
.C(n_427),
.Y(n_4894)
);

AND2x2_ASAP7_75t_L g4895 ( 
.A(n_4874),
.B(n_426),
.Y(n_4895)
);

AND2x2_ASAP7_75t_L g4896 ( 
.A(n_4876),
.B(n_427),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4846),
.Y(n_4897)
);

OAI32xp33_ASAP7_75t_L g4898 ( 
.A1(n_4832),
.A2(n_430),
.A3(n_428),
.B1(n_429),
.B2(n_431),
.Y(n_4898)
);

OAI22xp33_ASAP7_75t_L g4899 ( 
.A1(n_4873),
.A2(n_433),
.B1(n_429),
.B2(n_431),
.Y(n_4899)
);

NAND2xp5_ASAP7_75t_L g4900 ( 
.A(n_4833),
.B(n_433),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4879),
.Y(n_4901)
);

NAND2xp33_ASAP7_75t_SL g4902 ( 
.A(n_4855),
.B(n_434),
.Y(n_4902)
);

XOR2x2_ASAP7_75t_L g4903 ( 
.A(n_4837),
.B(n_434),
.Y(n_4903)
);

INVxp67_ASAP7_75t_L g4904 ( 
.A(n_4858),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4863),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4873),
.Y(n_4906)
);

NOR2x1_ASAP7_75t_SL g4907 ( 
.A(n_4881),
.B(n_435),
.Y(n_4907)
);

OAI32xp33_ASAP7_75t_L g4908 ( 
.A1(n_4841),
.A2(n_437),
.A3(n_435),
.B1(n_436),
.B2(n_438),
.Y(n_4908)
);

AOI221xp5_ASAP7_75t_L g4909 ( 
.A1(n_4880),
.A2(n_438),
.B1(n_436),
.B2(n_437),
.C(n_439),
.Y(n_4909)
);

A2O1A1Ixp33_ASAP7_75t_L g4910 ( 
.A1(n_4868),
.A2(n_441),
.B(n_439),
.C(n_440),
.Y(n_4910)
);

NOR2xp33_ASAP7_75t_L g4911 ( 
.A(n_4831),
.B(n_440),
.Y(n_4911)
);

AOI22xp5_ASAP7_75t_L g4912 ( 
.A1(n_4840),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4834),
.Y(n_4913)
);

INVx1_ASAP7_75t_L g4914 ( 
.A(n_4852),
.Y(n_4914)
);

BUFx3_ASAP7_75t_L g4915 ( 
.A(n_4857),
.Y(n_4915)
);

NAND2xp5_ASAP7_75t_L g4916 ( 
.A(n_4860),
.B(n_4851),
.Y(n_4916)
);

OR2x2_ASAP7_75t_L g4917 ( 
.A(n_4864),
.B(n_442),
.Y(n_4917)
);

OR2x2_ASAP7_75t_L g4918 ( 
.A(n_4869),
.B(n_443),
.Y(n_4918)
);

NAND3xp33_ASAP7_75t_L g4919 ( 
.A(n_4853),
.B(n_452),
.C(n_444),
.Y(n_4919)
);

NAND2xp5_ASAP7_75t_L g4920 ( 
.A(n_4861),
.B(n_445),
.Y(n_4920)
);

INVx2_ASAP7_75t_L g4921 ( 
.A(n_4867),
.Y(n_4921)
);

AND2x2_ASAP7_75t_L g4922 ( 
.A(n_4865),
.B(n_445),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4848),
.Y(n_4923)
);

AOI22xp33_ASAP7_75t_L g4924 ( 
.A1(n_4871),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.Y(n_4924)
);

OAI31xp33_ASAP7_75t_L g4925 ( 
.A1(n_4872),
.A2(n_450),
.A3(n_447),
.B(n_449),
.Y(n_4925)
);

AND2x2_ASAP7_75t_L g4926 ( 
.A(n_4866),
.B(n_450),
.Y(n_4926)
);

NAND2xp5_ASAP7_75t_L g4927 ( 
.A(n_4835),
.B(n_451),
.Y(n_4927)
);

NAND2xp5_ASAP7_75t_L g4928 ( 
.A(n_4845),
.B(n_451),
.Y(n_4928)
);

AND3x2_ASAP7_75t_L g4929 ( 
.A(n_4829),
.B(n_452),
.C(n_453),
.Y(n_4929)
);

AOI22xp33_ASAP7_75t_L g4930 ( 
.A1(n_4862),
.A2(n_455),
.B1(n_453),
.B2(n_454),
.Y(n_4930)
);

NAND2x1_ASAP7_75t_SL g4931 ( 
.A(n_4836),
.B(n_454),
.Y(n_4931)
);

NAND3xp33_ASAP7_75t_L g4932 ( 
.A(n_4839),
.B(n_466),
.C(n_456),
.Y(n_4932)
);

NAND2xp5_ASAP7_75t_L g4933 ( 
.A(n_4849),
.B(n_457),
.Y(n_4933)
);

OR2x2_ASAP7_75t_L g4934 ( 
.A(n_4859),
.B(n_458),
.Y(n_4934)
);

AOI21xp33_ASAP7_75t_SL g4935 ( 
.A1(n_4870),
.A2(n_458),
.B(n_460),
.Y(n_4935)
);

NOR4xp25_ASAP7_75t_SL g4936 ( 
.A(n_4830),
.B(n_462),
.C(n_460),
.D(n_461),
.Y(n_4936)
);

NAND3xp33_ASAP7_75t_L g4937 ( 
.A(n_4847),
.B(n_472),
.C(n_461),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4828),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4828),
.Y(n_4939)
);

NAND2xp5_ASAP7_75t_L g4940 ( 
.A(n_4828),
.B(n_464),
.Y(n_4940)
);

AOI21xp5_ASAP7_75t_L g4941 ( 
.A1(n_4847),
.A2(n_464),
.B(n_465),
.Y(n_4941)
);

AOI22xp33_ASAP7_75t_L g4942 ( 
.A1(n_4847),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_4942)
);

INVx2_ASAP7_75t_L g4943 ( 
.A(n_4828),
.Y(n_4943)
);

INVx2_ASAP7_75t_L g4944 ( 
.A(n_4828),
.Y(n_4944)
);

AND2x2_ASAP7_75t_L g4945 ( 
.A(n_4878),
.B(n_468),
.Y(n_4945)
);

AOI22xp5_ASAP7_75t_L g4946 ( 
.A1(n_4847),
.A2(n_472),
.B1(n_469),
.B2(n_470),
.Y(n_4946)
);

AND2x2_ASAP7_75t_L g4947 ( 
.A(n_4878),
.B(n_470),
.Y(n_4947)
);

NAND2xp5_ASAP7_75t_L g4948 ( 
.A(n_4828),
.B(n_473),
.Y(n_4948)
);

NOR2xp33_ASAP7_75t_L g4949 ( 
.A(n_4841),
.B(n_474),
.Y(n_4949)
);

OR2x2_ASAP7_75t_L g4950 ( 
.A(n_4847),
.B(n_474),
.Y(n_4950)
);

OAI21xp33_ASAP7_75t_SL g4951 ( 
.A1(n_4847),
.A2(n_476),
.B(n_477),
.Y(n_4951)
);

OAI322xp33_ASAP7_75t_L g4952 ( 
.A1(n_4847),
.A2(n_481),
.A3(n_480),
.B1(n_478),
.B2(n_476),
.C1(n_477),
.C2(n_479),
.Y(n_4952)
);

INVx1_ASAP7_75t_L g4953 ( 
.A(n_4828),
.Y(n_4953)
);

INVxp67_ASAP7_75t_L g4954 ( 
.A(n_4875),
.Y(n_4954)
);

AOI31xp33_ASAP7_75t_L g4955 ( 
.A1(n_4878),
.A2(n_480),
.A3(n_478),
.B(n_479),
.Y(n_4955)
);

A2O1A1Ixp33_ASAP7_75t_L g4956 ( 
.A1(n_4847),
.A2(n_483),
.B(n_481),
.C(n_482),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4828),
.Y(n_4957)
);

NOR2xp33_ASAP7_75t_L g4958 ( 
.A(n_4841),
.B(n_482),
.Y(n_4958)
);

OAI21xp33_ASAP7_75t_SL g4959 ( 
.A1(n_4847),
.A2(n_484),
.B(n_486),
.Y(n_4959)
);

NAND2xp5_ASAP7_75t_L g4960 ( 
.A(n_4828),
.B(n_484),
.Y(n_4960)
);

INVx3_ASAP7_75t_L g4961 ( 
.A(n_4844),
.Y(n_4961)
);

NAND2x1p5_ASAP7_75t_L g4962 ( 
.A(n_4844),
.B(n_487),
.Y(n_4962)
);

OAI22xp5_ASAP7_75t_L g4963 ( 
.A1(n_4847),
.A2(n_491),
.B1(n_488),
.B2(n_489),
.Y(n_4963)
);

AND2x4_ASAP7_75t_L g4964 ( 
.A(n_4878),
.B(n_488),
.Y(n_4964)
);

AND2x2_ASAP7_75t_L g4965 ( 
.A(n_4878),
.B(n_489),
.Y(n_4965)
);

INVx3_ASAP7_75t_L g4966 ( 
.A(n_4844),
.Y(n_4966)
);

INVx2_ASAP7_75t_L g4967 ( 
.A(n_4828),
.Y(n_4967)
);

NOR2xp33_ASAP7_75t_L g4968 ( 
.A(n_4841),
.B(n_492),
.Y(n_4968)
);

NOR3xp33_ASAP7_75t_L g4969 ( 
.A(n_4906),
.B(n_492),
.C(n_493),
.Y(n_4969)
);

AOI221xp5_ASAP7_75t_L g4970 ( 
.A1(n_4884),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.C(n_496),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4921),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4940),
.Y(n_4972)
);

NAND2xp33_ASAP7_75t_L g4973 ( 
.A(n_4950),
.B(n_495),
.Y(n_4973)
);

NAND2xp5_ASAP7_75t_L g4974 ( 
.A(n_4929),
.B(n_496),
.Y(n_4974)
);

NAND2xp5_ASAP7_75t_L g4975 ( 
.A(n_4901),
.B(n_497),
.Y(n_4975)
);

NOR2x1_ASAP7_75t_L g4976 ( 
.A(n_4937),
.B(n_497),
.Y(n_4976)
);

AOI221xp5_ASAP7_75t_L g4977 ( 
.A1(n_4951),
.A2(n_501),
.B1(n_498),
.B2(n_500),
.C(n_503),
.Y(n_4977)
);

INVx2_ASAP7_75t_L g4978 ( 
.A(n_4962),
.Y(n_4978)
);

NOR3xp33_ASAP7_75t_SL g4979 ( 
.A(n_4959),
.B(n_498),
.C(n_500),
.Y(n_4979)
);

NOR3x1_ASAP7_75t_L g4980 ( 
.A(n_4963),
.B(n_501),
.C(n_503),
.Y(n_4980)
);

INVxp67_ASAP7_75t_SL g4981 ( 
.A(n_4931),
.Y(n_4981)
);

INVx1_ASAP7_75t_SL g4982 ( 
.A(n_4902),
.Y(n_4982)
);

NAND3xp33_ASAP7_75t_SL g4983 ( 
.A(n_4936),
.B(n_504),
.C(n_505),
.Y(n_4983)
);

AOI221xp5_ASAP7_75t_SL g4984 ( 
.A1(n_4956),
.A2(n_506),
.B1(n_504),
.B2(n_505),
.C(n_507),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4948),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_4960),
.Y(n_4986)
);

AOI221xp5_ASAP7_75t_L g4987 ( 
.A1(n_4941),
.A2(n_509),
.B1(n_507),
.B2(n_508),
.C(n_510),
.Y(n_4987)
);

NAND2xp5_ASAP7_75t_SL g4988 ( 
.A(n_4887),
.B(n_508),
.Y(n_4988)
);

HB1xp67_ASAP7_75t_L g4989 ( 
.A(n_4903),
.Y(n_4989)
);

NOR3xp33_ASAP7_75t_SL g4990 ( 
.A(n_4888),
.B(n_509),
.C(n_510),
.Y(n_4990)
);

NAND2xp5_ASAP7_75t_SL g4991 ( 
.A(n_4909),
.B(n_511),
.Y(n_4991)
);

NAND2xp5_ASAP7_75t_L g4992 ( 
.A(n_4955),
.B(n_512),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4907),
.Y(n_4993)
);

XOR2x2_ASAP7_75t_L g4994 ( 
.A(n_4938),
.B(n_512),
.Y(n_4994)
);

OAI211xp5_ASAP7_75t_SL g4995 ( 
.A1(n_4942),
.A2(n_515),
.B(n_513),
.C(n_514),
.Y(n_4995)
);

NAND2xp5_ASAP7_75t_L g4996 ( 
.A(n_4882),
.B(n_513),
.Y(n_4996)
);

NOR4xp75_ASAP7_75t_L g4997 ( 
.A(n_4952),
.B(n_519),
.C(n_516),
.D(n_517),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_4943),
.B(n_516),
.Y(n_4998)
);

NAND3xp33_ASAP7_75t_SL g4999 ( 
.A(n_4946),
.B(n_520),
.C(n_521),
.Y(n_4999)
);

NAND2xp5_ASAP7_75t_L g5000 ( 
.A(n_4944),
.B(n_521),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4967),
.Y(n_5001)
);

AOI22xp5_ASAP7_75t_L g5002 ( 
.A1(n_4911),
.A2(n_524),
.B1(n_522),
.B2(n_523),
.Y(n_5002)
);

NAND2xp5_ASAP7_75t_L g5003 ( 
.A(n_4939),
.B(n_523),
.Y(n_5003)
);

AOI21xp5_ASAP7_75t_L g5004 ( 
.A1(n_4910),
.A2(n_524),
.B(n_525),
.Y(n_5004)
);

NAND3xp33_ASAP7_75t_SL g5005 ( 
.A(n_4925),
.B(n_526),
.C(n_528),
.Y(n_5005)
);

NOR3xp33_ASAP7_75t_SL g5006 ( 
.A(n_4889),
.B(n_530),
.C(n_531),
.Y(n_5006)
);

NAND3xp33_ASAP7_75t_L g5007 ( 
.A(n_4891),
.B(n_531),
.C(n_532),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4953),
.Y(n_5008)
);

BUFx12f_ASAP7_75t_L g5009 ( 
.A(n_4895),
.Y(n_5009)
);

OR2x2_ASAP7_75t_L g5010 ( 
.A(n_4961),
.B(n_532),
.Y(n_5010)
);

NAND3xp33_ASAP7_75t_L g5011 ( 
.A(n_4954),
.B(n_533),
.C(n_534),
.Y(n_5011)
);

NOR2xp33_ASAP7_75t_L g5012 ( 
.A(n_4957),
.B(n_535),
.Y(n_5012)
);

AOI22xp5_ASAP7_75t_L g5013 ( 
.A1(n_4905),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_5013)
);

NAND2xp5_ASAP7_75t_L g5014 ( 
.A(n_4883),
.B(n_536),
.Y(n_5014)
);

AOI21xp5_ASAP7_75t_L g5015 ( 
.A1(n_4916),
.A2(n_539),
.B(n_540),
.Y(n_5015)
);

INVx1_ASAP7_75t_SL g5016 ( 
.A(n_4892),
.Y(n_5016)
);

INVxp67_ASAP7_75t_L g5017 ( 
.A(n_4949),
.Y(n_5017)
);

INVx2_ASAP7_75t_L g5018 ( 
.A(n_4915),
.Y(n_5018)
);

NOR3xp33_ASAP7_75t_SL g5019 ( 
.A(n_4958),
.B(n_540),
.C(n_541),
.Y(n_5019)
);

HB1xp67_ASAP7_75t_L g5020 ( 
.A(n_4890),
.Y(n_5020)
);

AOI22xp5_ASAP7_75t_L g5021 ( 
.A1(n_4914),
.A2(n_545),
.B1(n_541),
.B2(n_543),
.Y(n_5021)
);

NAND2xp5_ASAP7_75t_L g5022 ( 
.A(n_4886),
.B(n_545),
.Y(n_5022)
);

NAND3xp33_ASAP7_75t_SL g5023 ( 
.A(n_4935),
.B(n_546),
.C(n_547),
.Y(n_5023)
);

INVxp67_ASAP7_75t_L g5024 ( 
.A(n_4968),
.Y(n_5024)
);

NOR2xp33_ASAP7_75t_SL g5025 ( 
.A(n_4922),
.B(n_546),
.Y(n_5025)
);

HB1xp67_ASAP7_75t_L g5026 ( 
.A(n_4964),
.Y(n_5026)
);

NAND3xp33_ASAP7_75t_L g5027 ( 
.A(n_4912),
.B(n_548),
.C(n_549),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_4885),
.Y(n_5028)
);

NOR3xp33_ASAP7_75t_L g5029 ( 
.A(n_4920),
.B(n_550),
.C(n_551),
.Y(n_5029)
);

NAND4xp25_ASAP7_75t_L g5030 ( 
.A(n_4896),
.B(n_553),
.C(n_554),
.D(n_552),
.Y(n_5030)
);

NOR2xp33_ASAP7_75t_L g5031 ( 
.A(n_4908),
.B(n_550),
.Y(n_5031)
);

NOR2xp67_ASAP7_75t_L g5032 ( 
.A(n_4966),
.B(n_552),
.Y(n_5032)
);

NOR2x1_ASAP7_75t_SL g5033 ( 
.A(n_4945),
.B(n_555),
.Y(n_5033)
);

AOI221xp5_ASAP7_75t_L g5034 ( 
.A1(n_4913),
.A2(n_4930),
.B1(n_4904),
.B2(n_4923),
.C(n_4897),
.Y(n_5034)
);

OAI221xp5_ASAP7_75t_SL g5035 ( 
.A1(n_4917),
.A2(n_558),
.B1(n_556),
.B2(n_557),
.C(n_560),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_4947),
.Y(n_5036)
);

NAND2xp5_ASAP7_75t_L g5037 ( 
.A(n_4893),
.B(n_556),
.Y(n_5037)
);

NOR2xp33_ASAP7_75t_L g5038 ( 
.A(n_4898),
.B(n_558),
.Y(n_5038)
);

AND2x2_ASAP7_75t_L g5039 ( 
.A(n_4965),
.B(n_4926),
.Y(n_5039)
);

AOI211xp5_ASAP7_75t_L g5040 ( 
.A1(n_4899),
.A2(n_562),
.B(n_560),
.C(n_561),
.Y(n_5040)
);

AOI22x1_ASAP7_75t_L g5041 ( 
.A1(n_4934),
.A2(n_563),
.B1(n_561),
.B2(n_562),
.Y(n_5041)
);

NOR3x1_ASAP7_75t_L g5042 ( 
.A(n_4919),
.B(n_563),
.C(n_564),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_4894),
.B(n_564),
.Y(n_5043)
);

NAND3xp33_ASAP7_75t_SL g5044 ( 
.A(n_4900),
.B(n_565),
.C(n_566),
.Y(n_5044)
);

BUFx2_ASAP7_75t_L g5045 ( 
.A(n_4918),
.Y(n_5045)
);

AND2x2_ASAP7_75t_L g5046 ( 
.A(n_4927),
.B(n_565),
.Y(n_5046)
);

INVxp67_ASAP7_75t_L g5047 ( 
.A(n_4933),
.Y(n_5047)
);

NAND3xp33_ASAP7_75t_L g5048 ( 
.A(n_4924),
.B(n_566),
.C(n_567),
.Y(n_5048)
);

AOI211xp5_ASAP7_75t_L g5049 ( 
.A1(n_4932),
.A2(n_571),
.B(n_568),
.C(n_569),
.Y(n_5049)
);

OAI21xp5_ASAP7_75t_L g5050 ( 
.A1(n_4928),
.A2(n_573),
.B(n_572),
.Y(n_5050)
);

NAND2xp5_ASAP7_75t_L g5051 ( 
.A(n_4929),
.B(n_571),
.Y(n_5051)
);

INVx2_ASAP7_75t_L g5052 ( 
.A(n_4962),
.Y(n_5052)
);

NOR2xp67_ASAP7_75t_L g5053 ( 
.A(n_4971),
.B(n_5018),
.Y(n_5053)
);

OAI221xp5_ASAP7_75t_SL g5054 ( 
.A1(n_4982),
.A2(n_575),
.B1(n_572),
.B2(n_574),
.C(n_578),
.Y(n_5054)
);

OAI22xp5_ASAP7_75t_L g5055 ( 
.A1(n_5008),
.A2(n_578),
.B1(n_574),
.B2(n_575),
.Y(n_5055)
);

AOI21xp33_ASAP7_75t_L g5056 ( 
.A1(n_4993),
.A2(n_579),
.B(n_580),
.Y(n_5056)
);

NOR3xp33_ASAP7_75t_L g5057 ( 
.A(n_5020),
.B(n_579),
.C(n_581),
.Y(n_5057)
);

NOR2xp33_ASAP7_75t_L g5058 ( 
.A(n_4983),
.B(n_581),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_L g5059 ( 
.A(n_4981),
.B(n_5033),
.Y(n_5059)
);

AOI21xp33_ASAP7_75t_SL g5060 ( 
.A1(n_4974),
.A2(n_5051),
.B(n_4992),
.Y(n_5060)
);

AOI21xp5_ASAP7_75t_L g5061 ( 
.A1(n_4988),
.A2(n_582),
.B(n_583),
.Y(n_5061)
);

NOR2xp33_ASAP7_75t_R g5062 ( 
.A(n_5028),
.B(n_584),
.Y(n_5062)
);

OAI211xp5_ASAP7_75t_SL g5063 ( 
.A1(n_5001),
.A2(n_586),
.B(n_584),
.C(n_585),
.Y(n_5063)
);

NAND3xp33_ASAP7_75t_L g5064 ( 
.A(n_4973),
.B(n_588),
.C(n_587),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_SL g5065 ( 
.A(n_4984),
.B(n_586),
.Y(n_5065)
);

OAI221xp5_ASAP7_75t_L g5066 ( 
.A1(n_5002),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.C(n_591),
.Y(n_5066)
);

AOI221xp5_ASAP7_75t_L g5067 ( 
.A1(n_5045),
.A2(n_592),
.B1(n_589),
.B2(n_591),
.C(n_594),
.Y(n_5067)
);

AND2x2_ASAP7_75t_L g5068 ( 
.A(n_5026),
.B(n_592),
.Y(n_5068)
);

NAND3xp33_ASAP7_75t_L g5069 ( 
.A(n_5025),
.B(n_596),
.C(n_595),
.Y(n_5069)
);

NAND3xp33_ASAP7_75t_L g5070 ( 
.A(n_5006),
.B(n_597),
.C(n_595),
.Y(n_5070)
);

OAI21xp5_ASAP7_75t_L g5071 ( 
.A1(n_5015),
.A2(n_594),
.B(n_597),
.Y(n_5071)
);

OAI222xp33_ASAP7_75t_L g5072 ( 
.A1(n_4976),
.A2(n_600),
.B1(n_602),
.B2(n_598),
.C1(n_599),
.C2(n_601),
.Y(n_5072)
);

NOR3xp33_ASAP7_75t_L g5073 ( 
.A(n_5034),
.B(n_599),
.C(n_600),
.Y(n_5073)
);

AND2x2_ASAP7_75t_L g5074 ( 
.A(n_4978),
.B(n_604),
.Y(n_5074)
);

NAND3xp33_ASAP7_75t_SL g5075 ( 
.A(n_5016),
.B(n_604),
.C(n_605),
.Y(n_5075)
);

NAND2xp5_ASAP7_75t_L g5076 ( 
.A(n_5032),
.B(n_605),
.Y(n_5076)
);

NAND3xp33_ASAP7_75t_SL g5077 ( 
.A(n_4997),
.B(n_606),
.C(n_607),
.Y(n_5077)
);

OAI21xp33_ASAP7_75t_L g5078 ( 
.A1(n_4975),
.A2(n_606),
.B(n_607),
.Y(n_5078)
);

OAI21xp5_ASAP7_75t_L g5079 ( 
.A1(n_5007),
.A2(n_608),
.B(n_609),
.Y(n_5079)
);

OAI221xp5_ASAP7_75t_L g5080 ( 
.A1(n_5052),
.A2(n_611),
.B1(n_609),
.B2(n_610),
.C(n_612),
.Y(n_5080)
);

NAND3xp33_ASAP7_75t_SL g5081 ( 
.A(n_4977),
.B(n_610),
.C(n_611),
.Y(n_5081)
);

INVx2_ASAP7_75t_L g5082 ( 
.A(n_5041),
.Y(n_5082)
);

AOI211xp5_ASAP7_75t_L g5083 ( 
.A1(n_5023),
.A2(n_616),
.B(n_613),
.C(n_614),
.Y(n_5083)
);

NAND2xp5_ASAP7_75t_L g5084 ( 
.A(n_5039),
.B(n_4990),
.Y(n_5084)
);

NAND4xp25_ASAP7_75t_L g5085 ( 
.A(n_5042),
.B(n_619),
.C(n_617),
.D(n_618),
.Y(n_5085)
);

NAND2xp5_ASAP7_75t_L g5086 ( 
.A(n_5012),
.B(n_617),
.Y(n_5086)
);

AOI211x1_ASAP7_75t_L g5087 ( 
.A1(n_4991),
.A2(n_5005),
.B(n_5044),
.C(n_5050),
.Y(n_5087)
);

OAI21xp33_ASAP7_75t_SL g5088 ( 
.A1(n_5036),
.A2(n_618),
.B(n_619),
.Y(n_5088)
);

AOI211xp5_ASAP7_75t_SL g5089 ( 
.A1(n_4989),
.A2(n_622),
.B(n_620),
.C(n_621),
.Y(n_5089)
);

NAND2xp5_ASAP7_75t_L g5090 ( 
.A(n_5029),
.B(n_620),
.Y(n_5090)
);

NOR4xp25_ASAP7_75t_L g5091 ( 
.A(n_5047),
.B(n_5024),
.C(n_5017),
.D(n_4985),
.Y(n_5091)
);

AOI22xp5_ASAP7_75t_L g5092 ( 
.A1(n_5009),
.A2(n_625),
.B1(n_621),
.B2(n_624),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4994),
.Y(n_5093)
);

OAI22xp5_ASAP7_75t_L g5094 ( 
.A1(n_5010),
.A2(n_626),
.B1(n_624),
.B2(n_625),
.Y(n_5094)
);

AOI222xp33_ASAP7_75t_L g5095 ( 
.A1(n_4972),
.A2(n_629),
.B1(n_633),
.B2(n_627),
.C1(n_628),
.C2(n_632),
.Y(n_5095)
);

NAND4xp25_ASAP7_75t_L g5096 ( 
.A(n_4980),
.B(n_629),
.C(n_627),
.D(n_628),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_5022),
.Y(n_5097)
);

AND3x1_ASAP7_75t_L g5098 ( 
.A(n_4979),
.B(n_632),
.C(n_633),
.Y(n_5098)
);

NAND2xp5_ASAP7_75t_L g5099 ( 
.A(n_4986),
.B(n_634),
.Y(n_5099)
);

AOI22xp5_ASAP7_75t_L g5100 ( 
.A1(n_5046),
.A2(n_636),
.B1(n_634),
.B2(n_635),
.Y(n_5100)
);

AOI221xp5_ASAP7_75t_L g5101 ( 
.A1(n_4999),
.A2(n_638),
.B1(n_636),
.B2(n_637),
.C(n_640),
.Y(n_5101)
);

AOI22xp33_ASAP7_75t_L g5102 ( 
.A1(n_4995),
.A2(n_642),
.B1(n_640),
.B2(n_641),
.Y(n_5102)
);

AOI22xp33_ASAP7_75t_SL g5103 ( 
.A1(n_5031),
.A2(n_643),
.B1(n_641),
.B2(n_642),
.Y(n_5103)
);

O2A1O1Ixp33_ASAP7_75t_SL g5104 ( 
.A1(n_5003),
.A2(n_647),
.B(n_645),
.C(n_646),
.Y(n_5104)
);

AOI221xp5_ASAP7_75t_L g5105 ( 
.A1(n_5004),
.A2(n_648),
.B1(n_645),
.B2(n_647),
.C(n_649),
.Y(n_5105)
);

NAND4xp25_ASAP7_75t_L g5106 ( 
.A(n_5049),
.B(n_651),
.C(n_649),
.D(n_650),
.Y(n_5106)
);

NOR2xp33_ASAP7_75t_L g5107 ( 
.A(n_5030),
.B(n_650),
.Y(n_5107)
);

OAI211xp5_ASAP7_75t_SL g5108 ( 
.A1(n_4970),
.A2(n_654),
.B(n_652),
.C(n_653),
.Y(n_5108)
);

AND2x2_ASAP7_75t_L g5109 ( 
.A(n_5038),
.B(n_652),
.Y(n_5109)
);

NOR2xp33_ASAP7_75t_L g5110 ( 
.A(n_5035),
.B(n_653),
.Y(n_5110)
);

NAND2xp5_ASAP7_75t_L g5111 ( 
.A(n_5019),
.B(n_654),
.Y(n_5111)
);

AOI21xp5_ASAP7_75t_SL g5112 ( 
.A1(n_5014),
.A2(n_665),
.B(n_656),
.Y(n_5112)
);

OAI221xp5_ASAP7_75t_L g5113 ( 
.A1(n_4996),
.A2(n_659),
.B1(n_656),
.B2(n_658),
.C(n_660),
.Y(n_5113)
);

AOI211xp5_ASAP7_75t_L g5114 ( 
.A1(n_5027),
.A2(n_661),
.B(n_659),
.C(n_660),
.Y(n_5114)
);

AOI22xp5_ASAP7_75t_L g5115 ( 
.A1(n_4998),
.A2(n_664),
.B1(n_662),
.B2(n_663),
.Y(n_5115)
);

AOI211xp5_ASAP7_75t_SL g5116 ( 
.A1(n_5000),
.A2(n_665),
.B(n_662),
.C(n_663),
.Y(n_5116)
);

OAI21xp5_ASAP7_75t_SL g5117 ( 
.A1(n_5037),
.A2(n_666),
.B(n_668),
.Y(n_5117)
);

XNOR2xp5_ASAP7_75t_L g5118 ( 
.A(n_5040),
.B(n_670),
.Y(n_5118)
);

NAND2xp5_ASAP7_75t_L g5119 ( 
.A(n_4969),
.B(n_668),
.Y(n_5119)
);

NOR2xp33_ASAP7_75t_L g5120 ( 
.A(n_5011),
.B(n_670),
.Y(n_5120)
);

AOI221xp5_ASAP7_75t_L g5121 ( 
.A1(n_4987),
.A2(n_5048),
.B1(n_5043),
.B2(n_5013),
.C(n_5021),
.Y(n_5121)
);

NOR3xp33_ASAP7_75t_L g5122 ( 
.A(n_5020),
.B(n_671),
.C(n_672),
.Y(n_5122)
);

AND2x2_ASAP7_75t_L g5123 ( 
.A(n_4971),
.B(n_671),
.Y(n_5123)
);

OAI221xp5_ASAP7_75t_SL g5124 ( 
.A1(n_4982),
.A2(n_675),
.B1(n_673),
.B2(n_674),
.C(n_676),
.Y(n_5124)
);

AOI322xp5_ASAP7_75t_L g5125 ( 
.A1(n_4993),
.A2(n_682),
.A3(n_681),
.B1(n_679),
.B2(n_675),
.C1(n_677),
.C2(n_680),
.Y(n_5125)
);

NOR3xp33_ASAP7_75t_L g5126 ( 
.A(n_5020),
.B(n_679),
.C(n_681),
.Y(n_5126)
);

AOI222xp33_ASAP7_75t_L g5127 ( 
.A1(n_4993),
.A2(n_684),
.B1(n_686),
.B2(n_682),
.C1(n_683),
.C2(n_685),
.Y(n_5127)
);

O2A1O1Ixp33_ASAP7_75t_L g5128 ( 
.A1(n_4981),
.A2(n_686),
.B(n_684),
.C(n_685),
.Y(n_5128)
);

OAI221xp5_ASAP7_75t_SL g5129 ( 
.A1(n_4982),
.A2(n_689),
.B1(n_687),
.B2(n_688),
.C(n_690),
.Y(n_5129)
);

NAND4xp75_ASAP7_75t_L g5130 ( 
.A(n_4976),
.B(n_691),
.C(n_687),
.D(n_689),
.Y(n_5130)
);

A2O1A1Ixp33_ASAP7_75t_L g5131 ( 
.A1(n_4993),
.A2(n_699),
.B(n_708),
.C(n_691),
.Y(n_5131)
);

OAI211xp5_ASAP7_75t_L g5132 ( 
.A1(n_4971),
.A2(n_694),
.B(n_692),
.C(n_693),
.Y(n_5132)
);

OAI21xp33_ASAP7_75t_L g5133 ( 
.A1(n_4971),
.A2(n_694),
.B(n_695),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_5020),
.Y(n_5134)
);

AOI21xp33_ASAP7_75t_SL g5135 ( 
.A1(n_4993),
.A2(n_695),
.B(n_696),
.Y(n_5135)
);

O2A1O1Ixp33_ASAP7_75t_L g5136 ( 
.A1(n_4981),
.A2(n_699),
.B(n_697),
.C(n_698),
.Y(n_5136)
);

OAI31xp33_ASAP7_75t_L g5137 ( 
.A1(n_4993),
.A2(n_708),
.A3(n_716),
.B(n_698),
.Y(n_5137)
);

AOI21xp5_ASAP7_75t_L g5138 ( 
.A1(n_4971),
.A2(n_700),
.B(n_702),
.Y(n_5138)
);

O2A1O1Ixp33_ASAP7_75t_L g5139 ( 
.A1(n_5059),
.A2(n_705),
.B(n_703),
.C(n_704),
.Y(n_5139)
);

OAI221xp5_ASAP7_75t_L g5140 ( 
.A1(n_5134),
.A2(n_706),
.B1(n_703),
.B2(n_705),
.C(n_707),
.Y(n_5140)
);

OAI211xp5_ASAP7_75t_L g5141 ( 
.A1(n_5053),
.A2(n_710),
.B(n_707),
.C(n_709),
.Y(n_5141)
);

OAI211xp5_ASAP7_75t_L g5142 ( 
.A1(n_5088),
.A2(n_711),
.B(n_709),
.C(n_710),
.Y(n_5142)
);

AOI21xp5_ASAP7_75t_L g5143 ( 
.A1(n_5131),
.A2(n_711),
.B(n_712),
.Y(n_5143)
);

A2O1A1O1Ixp25_ASAP7_75t_L g5144 ( 
.A1(n_5093),
.A2(n_715),
.B(n_713),
.C(n_714),
.D(n_716),
.Y(n_5144)
);

NAND4xp25_ASAP7_75t_L g5145 ( 
.A(n_5103),
.B(n_717),
.C(n_713),
.D(n_715),
.Y(n_5145)
);

AOI22xp33_ASAP7_75t_SL g5146 ( 
.A1(n_5109),
.A2(n_5058),
.B1(n_5068),
.B2(n_5084),
.Y(n_5146)
);

NAND2xp5_ASAP7_75t_SL g5147 ( 
.A(n_5135),
.B(n_717),
.Y(n_5147)
);

OAI211xp5_ASAP7_75t_L g5148 ( 
.A1(n_5137),
.A2(n_721),
.B(n_718),
.C(n_719),
.Y(n_5148)
);

AOI22xp33_ASAP7_75t_L g5149 ( 
.A1(n_5077),
.A2(n_722),
.B1(n_718),
.B2(n_719),
.Y(n_5149)
);

O2A1O1Ixp33_ASAP7_75t_L g5150 ( 
.A1(n_5060),
.A2(n_727),
.B(n_724),
.C(n_725),
.Y(n_5150)
);

NAND2xp5_ASAP7_75t_SL g5151 ( 
.A(n_5127),
.B(n_724),
.Y(n_5151)
);

OAI211xp5_ASAP7_75t_L g5152 ( 
.A1(n_5065),
.A2(n_729),
.B(n_725),
.C(n_728),
.Y(n_5152)
);

NAND2xp5_ASAP7_75t_L g5153 ( 
.A(n_5089),
.B(n_730),
.Y(n_5153)
);

NAND2xp5_ASAP7_75t_L g5154 ( 
.A(n_5116),
.B(n_730),
.Y(n_5154)
);

NOR3xp33_ASAP7_75t_L g5155 ( 
.A(n_5099),
.B(n_729),
.C(n_731),
.Y(n_5155)
);

AOI321xp33_ASAP7_75t_L g5156 ( 
.A1(n_5091),
.A2(n_734),
.A3(n_736),
.B1(n_732),
.B2(n_733),
.C(n_735),
.Y(n_5156)
);

AOI221xp5_ASAP7_75t_L g5157 ( 
.A1(n_5061),
.A2(n_738),
.B1(n_734),
.B2(n_737),
.C(n_739),
.Y(n_5157)
);

AOI221xp5_ASAP7_75t_L g5158 ( 
.A1(n_5121),
.A2(n_739),
.B1(n_737),
.B2(n_738),
.C(n_740),
.Y(n_5158)
);

OAI21xp33_ASAP7_75t_L g5159 ( 
.A1(n_5085),
.A2(n_740),
.B(n_741),
.Y(n_5159)
);

NAND2xp5_ASAP7_75t_L g5160 ( 
.A(n_5123),
.B(n_742),
.Y(n_5160)
);

OAI221xp5_ASAP7_75t_L g5161 ( 
.A1(n_5133),
.A2(n_744),
.B1(n_741),
.B2(n_743),
.C(n_745),
.Y(n_5161)
);

O2A1O1Ixp33_ASAP7_75t_L g5162 ( 
.A1(n_5072),
.A2(n_745),
.B(n_743),
.C(n_744),
.Y(n_5162)
);

AOI221x1_ASAP7_75t_L g5163 ( 
.A1(n_5073),
.A2(n_750),
.B1(n_746),
.B2(n_748),
.C(n_751),
.Y(n_5163)
);

AO21x1_ASAP7_75t_L g5164 ( 
.A1(n_5110),
.A2(n_746),
.B(n_748),
.Y(n_5164)
);

AOI21xp5_ASAP7_75t_L g5165 ( 
.A1(n_5128),
.A2(n_750),
.B(n_752),
.Y(n_5165)
);

NAND2xp5_ASAP7_75t_SL g5166 ( 
.A(n_5095),
.B(n_752),
.Y(n_5166)
);

AOI221xp5_ASAP7_75t_L g5167 ( 
.A1(n_5071),
.A2(n_5097),
.B1(n_5087),
.B2(n_5098),
.C(n_5075),
.Y(n_5167)
);

NAND2xp5_ASAP7_75t_L g5168 ( 
.A(n_5082),
.B(n_754),
.Y(n_5168)
);

AOI21xp33_ASAP7_75t_L g5169 ( 
.A1(n_5070),
.A2(n_753),
.B(n_756),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_5076),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_L g5171 ( 
.A(n_5102),
.B(n_757),
.Y(n_5171)
);

AOI22xp5_ASAP7_75t_L g5172 ( 
.A1(n_5107),
.A2(n_758),
.B1(n_756),
.B2(n_757),
.Y(n_5172)
);

AOI21xp5_ASAP7_75t_L g5173 ( 
.A1(n_5136),
.A2(n_759),
.B(n_760),
.Y(n_5173)
);

O2A1O1Ixp33_ASAP7_75t_L g5174 ( 
.A1(n_5056),
.A2(n_762),
.B(n_760),
.C(n_761),
.Y(n_5174)
);

OAI311xp33_ASAP7_75t_L g5175 ( 
.A1(n_5096),
.A2(n_764),
.A3(n_762),
.B1(n_763),
.C1(n_765),
.Y(n_5175)
);

AOI22xp5_ASAP7_75t_L g5176 ( 
.A1(n_5120),
.A2(n_768),
.B1(n_763),
.B2(n_767),
.Y(n_5176)
);

AOI21xp5_ASAP7_75t_L g5177 ( 
.A1(n_5104),
.A2(n_767),
.B(n_768),
.Y(n_5177)
);

AOI221x1_ASAP7_75t_L g5178 ( 
.A1(n_5057),
.A2(n_771),
.B1(n_769),
.B2(n_770),
.C(n_772),
.Y(n_5178)
);

OAI21xp33_ASAP7_75t_L g5179 ( 
.A1(n_5106),
.A2(n_769),
.B(n_770),
.Y(n_5179)
);

AOI21xp5_ASAP7_75t_L g5180 ( 
.A1(n_5138),
.A2(n_771),
.B(n_772),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_5074),
.B(n_774),
.Y(n_5181)
);

OAI211xp5_ASAP7_75t_SL g5182 ( 
.A1(n_5079),
.A2(n_775),
.B(n_773),
.C(n_774),
.Y(n_5182)
);

OAI221xp5_ASAP7_75t_L g5183 ( 
.A1(n_5117),
.A2(n_777),
.B1(n_773),
.B2(n_776),
.C(n_778),
.Y(n_5183)
);

NAND2xp5_ASAP7_75t_L g5184 ( 
.A(n_5083),
.B(n_777),
.Y(n_5184)
);

NAND2xp5_ASAP7_75t_SL g5185 ( 
.A(n_5101),
.B(n_776),
.Y(n_5185)
);

OAI211xp5_ASAP7_75t_SL g5186 ( 
.A1(n_5112),
.A2(n_782),
.B(n_778),
.C(n_781),
.Y(n_5186)
);

AOI22xp5_ASAP7_75t_L g5187 ( 
.A1(n_5086),
.A2(n_785),
.B1(n_783),
.B2(n_784),
.Y(n_5187)
);

INVxp67_ASAP7_75t_SL g5188 ( 
.A(n_5111),
.Y(n_5188)
);

AOI221x1_ASAP7_75t_L g5189 ( 
.A1(n_5122),
.A2(n_786),
.B1(n_783),
.B2(n_785),
.C(n_788),
.Y(n_5189)
);

NOR3xp33_ASAP7_75t_L g5190 ( 
.A(n_5126),
.B(n_789),
.C(n_790),
.Y(n_5190)
);

OAI221xp5_ASAP7_75t_L g5191 ( 
.A1(n_5114),
.A2(n_792),
.B1(n_789),
.B2(n_791),
.C(n_793),
.Y(n_5191)
);

OR2x2_ASAP7_75t_L g5192 ( 
.A(n_5119),
.B(n_791),
.Y(n_5192)
);

OAI21xp33_ASAP7_75t_L g5193 ( 
.A1(n_5108),
.A2(n_792),
.B(n_794),
.Y(n_5193)
);

AOI222xp33_ASAP7_75t_L g5194 ( 
.A1(n_5081),
.A2(n_796),
.B1(n_799),
.B2(n_800),
.C1(n_795),
.C2(n_797),
.Y(n_5194)
);

OAI211xp5_ASAP7_75t_L g5195 ( 
.A1(n_5132),
.A2(n_797),
.B(n_794),
.C(n_795),
.Y(n_5195)
);

OAI211xp5_ASAP7_75t_L g5196 ( 
.A1(n_5067),
.A2(n_803),
.B(n_801),
.C(n_802),
.Y(n_5196)
);

AOI22xp5_ASAP7_75t_L g5197 ( 
.A1(n_5078),
.A2(n_805),
.B1(n_802),
.B2(n_804),
.Y(n_5197)
);

AOI211xp5_ASAP7_75t_L g5198 ( 
.A1(n_5054),
.A2(n_808),
.B(n_804),
.C(n_806),
.Y(n_5198)
);

OAI21xp5_ASAP7_75t_L g5199 ( 
.A1(n_5064),
.A2(n_808),
.B(n_809),
.Y(n_5199)
);

AOI221xp5_ASAP7_75t_L g5200 ( 
.A1(n_5066),
.A2(n_813),
.B1(n_810),
.B2(n_811),
.C(n_814),
.Y(n_5200)
);

NAND2xp5_ASAP7_75t_L g5201 ( 
.A(n_5125),
.B(n_811),
.Y(n_5201)
);

AOI322xp5_ASAP7_75t_L g5202 ( 
.A1(n_5090),
.A2(n_818),
.A3(n_817),
.B1(n_815),
.B2(n_810),
.C1(n_814),
.C2(n_816),
.Y(n_5202)
);

AOI221x1_ASAP7_75t_L g5203 ( 
.A1(n_5094),
.A2(n_817),
.B1(n_815),
.B2(n_816),
.C(n_818),
.Y(n_5203)
);

NOR2xp67_ASAP7_75t_L g5204 ( 
.A(n_5092),
.B(n_820),
.Y(n_5204)
);

AND4x1_ASAP7_75t_L g5205 ( 
.A(n_5105),
.B(n_822),
.C(n_819),
.D(n_821),
.Y(n_5205)
);

NAND3xp33_ASAP7_75t_SL g5206 ( 
.A(n_5062),
.B(n_821),
.C(n_823),
.Y(n_5206)
);

AOI221xp5_ASAP7_75t_L g5207 ( 
.A1(n_5113),
.A2(n_825),
.B1(n_823),
.B2(n_824),
.C(n_826),
.Y(n_5207)
);

NAND2xp33_ASAP7_75t_SL g5208 ( 
.A(n_5118),
.B(n_825),
.Y(n_5208)
);

OAI221xp5_ASAP7_75t_L g5209 ( 
.A1(n_5124),
.A2(n_828),
.B1(n_826),
.B2(n_827),
.C(n_829),
.Y(n_5209)
);

OAI211xp5_ASAP7_75t_SL g5210 ( 
.A1(n_5080),
.A2(n_5115),
.B(n_5100),
.C(n_5069),
.Y(n_5210)
);

AOI21xp5_ASAP7_75t_L g5211 ( 
.A1(n_5129),
.A2(n_5055),
.B(n_5063),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_5130),
.Y(n_5212)
);

INVx3_ASAP7_75t_L g5213 ( 
.A(n_5134),
.Y(n_5213)
);

A2O1A1Ixp33_ASAP7_75t_L g5214 ( 
.A1(n_5134),
.A2(n_831),
.B(n_827),
.C(n_829),
.Y(n_5214)
);

AND2x2_ASAP7_75t_L g5215 ( 
.A(n_5134),
.B(n_831),
.Y(n_5215)
);

AOI22xp5_ASAP7_75t_L g5216 ( 
.A1(n_5188),
.A2(n_834),
.B1(n_832),
.B2(n_833),
.Y(n_5216)
);

NAND3x1_ASAP7_75t_SL g5217 ( 
.A(n_5158),
.B(n_843),
.C(n_833),
.Y(n_5217)
);

OAI221xp5_ASAP7_75t_SL g5218 ( 
.A1(n_5149),
.A2(n_837),
.B1(n_839),
.B2(n_836),
.C(n_838),
.Y(n_5218)
);

NAND2xp5_ASAP7_75t_SL g5219 ( 
.A(n_5156),
.B(n_835),
.Y(n_5219)
);

AOI21xp5_ASAP7_75t_L g5220 ( 
.A1(n_5168),
.A2(n_836),
.B(n_840),
.Y(n_5220)
);

OAI22xp5_ASAP7_75t_L g5221 ( 
.A1(n_5213),
.A2(n_844),
.B1(n_840),
.B2(n_841),
.Y(n_5221)
);

AOI21xp5_ASAP7_75t_L g5222 ( 
.A1(n_5139),
.A2(n_841),
.B(n_844),
.Y(n_5222)
);

OAI211xp5_ASAP7_75t_SL g5223 ( 
.A1(n_5167),
.A2(n_847),
.B(n_845),
.C(n_846),
.Y(n_5223)
);

AOI22xp5_ASAP7_75t_L g5224 ( 
.A1(n_5213),
.A2(n_847),
.B1(n_845),
.B2(n_846),
.Y(n_5224)
);

AND2x2_ASAP7_75t_L g5225 ( 
.A(n_5215),
.B(n_848),
.Y(n_5225)
);

NOR2xp33_ASAP7_75t_L g5226 ( 
.A(n_5142),
.B(n_849),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_5154),
.Y(n_5227)
);

AOI221x1_ASAP7_75t_L g5228 ( 
.A1(n_5201),
.A2(n_851),
.B1(n_849),
.B2(n_850),
.C(n_852),
.Y(n_5228)
);

AOI221xp5_ASAP7_75t_L g5229 ( 
.A1(n_5169),
.A2(n_852),
.B1(n_850),
.B2(n_851),
.C(n_853),
.Y(n_5229)
);

NAND2xp5_ASAP7_75t_L g5230 ( 
.A(n_5177),
.B(n_853),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_5153),
.Y(n_5231)
);

AND4x2_ASAP7_75t_L g5232 ( 
.A(n_5211),
.B(n_856),
.C(n_857),
.D(n_855),
.Y(n_5232)
);

AOI221x1_ASAP7_75t_L g5233 ( 
.A1(n_5159),
.A2(n_858),
.B1(n_854),
.B2(n_855),
.C(n_859),
.Y(n_5233)
);

OR2x2_ASAP7_75t_L g5234 ( 
.A(n_5147),
.B(n_854),
.Y(n_5234)
);

OAI21xp33_ASAP7_75t_L g5235 ( 
.A1(n_5179),
.A2(n_858),
.B(n_860),
.Y(n_5235)
);

A2O1A1Ixp33_ASAP7_75t_L g5236 ( 
.A1(n_5150),
.A2(n_864),
.B(n_862),
.C(n_863),
.Y(n_5236)
);

OA211x2_ASAP7_75t_L g5237 ( 
.A1(n_5157),
.A2(n_865),
.B(n_863),
.C(n_864),
.Y(n_5237)
);

NAND4xp75_ASAP7_75t_L g5238 ( 
.A(n_5164),
.B(n_867),
.C(n_865),
.D(n_866),
.Y(n_5238)
);

AOI222xp33_ASAP7_75t_L g5239 ( 
.A1(n_5208),
.A2(n_5212),
.B1(n_5151),
.B2(n_5166),
.C1(n_5170),
.C2(n_5206),
.Y(n_5239)
);

NAND4xp75_ASAP7_75t_L g5240 ( 
.A(n_5204),
.B(n_871),
.C(n_868),
.D(n_869),
.Y(n_5240)
);

AOI21xp5_ASAP7_75t_L g5241 ( 
.A1(n_5214),
.A2(n_868),
.B(n_869),
.Y(n_5241)
);

OAI22xp33_ASAP7_75t_L g5242 ( 
.A1(n_5172),
.A2(n_873),
.B1(n_871),
.B2(n_872),
.Y(n_5242)
);

NAND2xp5_ASAP7_75t_L g5243 ( 
.A(n_5146),
.B(n_873),
.Y(n_5243)
);

AOI22xp5_ASAP7_75t_L g5244 ( 
.A1(n_5152),
.A2(n_877),
.B1(n_874),
.B2(n_875),
.Y(n_5244)
);

AOI211xp5_ASAP7_75t_L g5245 ( 
.A1(n_5175),
.A2(n_880),
.B(n_875),
.C(n_879),
.Y(n_5245)
);

NAND2xp33_ASAP7_75t_SL g5246 ( 
.A(n_5184),
.B(n_880),
.Y(n_5246)
);

AOI22xp5_ASAP7_75t_L g5247 ( 
.A1(n_5182),
.A2(n_883),
.B1(n_881),
.B2(n_882),
.Y(n_5247)
);

AOI22xp5_ASAP7_75t_L g5248 ( 
.A1(n_5155),
.A2(n_884),
.B1(n_881),
.B2(n_882),
.Y(n_5248)
);

OAI211xp5_ASAP7_75t_SL g5249 ( 
.A1(n_5194),
.A2(n_887),
.B(n_885),
.C(n_886),
.Y(n_5249)
);

OAI221xp5_ASAP7_75t_L g5250 ( 
.A1(n_5209),
.A2(n_888),
.B1(n_886),
.B2(n_887),
.C(n_889),
.Y(n_5250)
);

OAI211xp5_ASAP7_75t_SL g5251 ( 
.A1(n_5185),
.A2(n_891),
.B(n_888),
.C(n_890),
.Y(n_5251)
);

OAI22xp33_ASAP7_75t_L g5252 ( 
.A1(n_5176),
.A2(n_892),
.B1(n_890),
.B2(n_891),
.Y(n_5252)
);

AOI21xp5_ASAP7_75t_L g5253 ( 
.A1(n_5162),
.A2(n_893),
.B(n_894),
.Y(n_5253)
);

AOI221xp5_ASAP7_75t_L g5254 ( 
.A1(n_5210),
.A2(n_5173),
.B1(n_5165),
.B2(n_5143),
.C(n_5193),
.Y(n_5254)
);

NAND2xp33_ASAP7_75t_L g5255 ( 
.A(n_5190),
.B(n_895),
.Y(n_5255)
);

OAI211xp5_ASAP7_75t_SL g5256 ( 
.A1(n_5198),
.A2(n_899),
.B(n_896),
.C(n_898),
.Y(n_5256)
);

OAI222xp33_ASAP7_75t_L g5257 ( 
.A1(n_5171),
.A2(n_5180),
.B1(n_5192),
.B2(n_5183),
.C1(n_5191),
.C2(n_5197),
.Y(n_5257)
);

AOI32xp33_ASAP7_75t_L g5258 ( 
.A1(n_5186),
.A2(n_899),
.A3(n_896),
.B1(n_898),
.B2(n_900),
.Y(n_5258)
);

AOI221xp5_ASAP7_75t_SL g5259 ( 
.A1(n_5174),
.A2(n_902),
.B1(n_900),
.B2(n_901),
.C(n_904),
.Y(n_5259)
);

OAI22xp33_ASAP7_75t_L g5260 ( 
.A1(n_5160),
.A2(n_904),
.B1(n_901),
.B2(n_902),
.Y(n_5260)
);

OAI211xp5_ASAP7_75t_SL g5261 ( 
.A1(n_5207),
.A2(n_907),
.B(n_905),
.C(n_906),
.Y(n_5261)
);

AOI33xp33_ASAP7_75t_L g5262 ( 
.A1(n_5200),
.A2(n_908),
.A3(n_911),
.B1(n_905),
.B2(n_906),
.B3(n_910),
.Y(n_5262)
);

AOI21xp5_ASAP7_75t_L g5263 ( 
.A1(n_5161),
.A2(n_908),
.B(n_911),
.Y(n_5263)
);

AOI221xp5_ASAP7_75t_L g5264 ( 
.A1(n_5199),
.A2(n_915),
.B1(n_912),
.B2(n_914),
.C(n_916),
.Y(n_5264)
);

AOI211x1_ASAP7_75t_SL g5265 ( 
.A1(n_5145),
.A2(n_5181),
.B(n_5144),
.C(n_5148),
.Y(n_5265)
);

AOI221xp5_ASAP7_75t_L g5266 ( 
.A1(n_5195),
.A2(n_917),
.B1(n_912),
.B2(n_916),
.C(n_919),
.Y(n_5266)
);

AOI211xp5_ASAP7_75t_L g5267 ( 
.A1(n_5196),
.A2(n_921),
.B(n_919),
.C(n_920),
.Y(n_5267)
);

NAND3xp33_ASAP7_75t_SL g5268 ( 
.A(n_5141),
.B(n_5205),
.C(n_5187),
.Y(n_5268)
);

A2O1A1Ixp33_ASAP7_75t_L g5269 ( 
.A1(n_5202),
.A2(n_923),
.B(n_921),
.C(n_922),
.Y(n_5269)
);

NAND2xp5_ASAP7_75t_L g5270 ( 
.A(n_5178),
.B(n_923),
.Y(n_5270)
);

AOI221xp5_ASAP7_75t_L g5271 ( 
.A1(n_5140),
.A2(n_926),
.B1(n_924),
.B2(n_925),
.C(n_927),
.Y(n_5271)
);

AOI21xp5_ASAP7_75t_L g5272 ( 
.A1(n_5219),
.A2(n_5189),
.B(n_5203),
.Y(n_5272)
);

NAND4xp75_ASAP7_75t_L g5273 ( 
.A(n_5228),
.B(n_5163),
.C(n_927),
.D(n_925),
.Y(n_5273)
);

INVx1_ASAP7_75t_L g5274 ( 
.A(n_5232),
.Y(n_5274)
);

NAND4xp75_ASAP7_75t_L g5275 ( 
.A(n_5243),
.B(n_929),
.C(n_926),
.D(n_928),
.Y(n_5275)
);

INVx1_ASAP7_75t_L g5276 ( 
.A(n_5238),
.Y(n_5276)
);

NAND2xp5_ASAP7_75t_L g5277 ( 
.A(n_5245),
.B(n_930),
.Y(n_5277)
);

AND2x2_ASAP7_75t_L g5278 ( 
.A(n_5225),
.B(n_931),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5270),
.Y(n_5279)
);

NOR4xp75_ASAP7_75t_L g5280 ( 
.A(n_5230),
.B(n_935),
.C(n_931),
.D(n_932),
.Y(n_5280)
);

NOR2xp33_ASAP7_75t_L g5281 ( 
.A(n_5223),
.B(n_932),
.Y(n_5281)
);

NAND4xp75_ASAP7_75t_L g5282 ( 
.A(n_5227),
.B(n_937),
.C(n_935),
.D(n_936),
.Y(n_5282)
);

XOR2x1_ASAP7_75t_L g5283 ( 
.A(n_5237),
.B(n_936),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_5240),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_5217),
.Y(n_5285)
);

NAND3xp33_ASAP7_75t_L g5286 ( 
.A(n_5239),
.B(n_937),
.C(n_938),
.Y(n_5286)
);

INVx1_ASAP7_75t_L g5287 ( 
.A(n_5265),
.Y(n_5287)
);

INVx1_ASAP7_75t_L g5288 ( 
.A(n_5234),
.Y(n_5288)
);

NOR3xp33_ASAP7_75t_L g5289 ( 
.A(n_5231),
.B(n_939),
.C(n_940),
.Y(n_5289)
);

NAND4xp75_ASAP7_75t_L g5290 ( 
.A(n_5233),
.B(n_941),
.C(n_939),
.D(n_940),
.Y(n_5290)
);

NAND2xp5_ASAP7_75t_L g5291 ( 
.A(n_5258),
.B(n_942),
.Y(n_5291)
);

INVxp67_ASAP7_75t_L g5292 ( 
.A(n_5226),
.Y(n_5292)
);

NAND3xp33_ASAP7_75t_L g5293 ( 
.A(n_5246),
.B(n_942),
.C(n_943),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_5247),
.Y(n_5294)
);

NOR2x1_ASAP7_75t_L g5295 ( 
.A(n_5221),
.B(n_5260),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_5262),
.Y(n_5296)
);

AOI22xp5_ASAP7_75t_L g5297 ( 
.A1(n_5235),
.A2(n_947),
.B1(n_944),
.B2(n_945),
.Y(n_5297)
);

NOR2xp33_ASAP7_75t_L g5298 ( 
.A(n_5256),
.B(n_944),
.Y(n_5298)
);

INVx1_ASAP7_75t_L g5299 ( 
.A(n_5244),
.Y(n_5299)
);

INVx1_ASAP7_75t_L g5300 ( 
.A(n_5268),
.Y(n_5300)
);

HB1xp67_ASAP7_75t_L g5301 ( 
.A(n_5267),
.Y(n_5301)
);

INVx2_ASAP7_75t_L g5302 ( 
.A(n_5248),
.Y(n_5302)
);

NOR3xp33_ASAP7_75t_L g5303 ( 
.A(n_5249),
.B(n_945),
.C(n_948),
.Y(n_5303)
);

NOR3xp33_ASAP7_75t_L g5304 ( 
.A(n_5255),
.B(n_948),
.C(n_949),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_5251),
.Y(n_5305)
);

NOR2xp33_ASAP7_75t_L g5306 ( 
.A(n_5257),
.B(n_5261),
.Y(n_5306)
);

INVxp67_ASAP7_75t_L g5307 ( 
.A(n_5278),
.Y(n_5307)
);

NOR3xp33_ASAP7_75t_L g5308 ( 
.A(n_5287),
.B(n_5229),
.C(n_5218),
.Y(n_5308)
);

INVx2_ASAP7_75t_L g5309 ( 
.A(n_5283),
.Y(n_5309)
);

AND2x4_ASAP7_75t_L g5310 ( 
.A(n_5300),
.B(n_5269),
.Y(n_5310)
);

NOR2xp67_ASAP7_75t_L g5311 ( 
.A(n_5286),
.B(n_5216),
.Y(n_5311)
);

NOR3xp33_ASAP7_75t_L g5312 ( 
.A(n_5279),
.B(n_5220),
.C(n_5254),
.Y(n_5312)
);

NAND2xp5_ASAP7_75t_L g5313 ( 
.A(n_5274),
.B(n_5259),
.Y(n_5313)
);

NAND3xp33_ASAP7_75t_L g5314 ( 
.A(n_5306),
.B(n_5266),
.C(n_5264),
.Y(n_5314)
);

NAND3xp33_ASAP7_75t_L g5315 ( 
.A(n_5276),
.B(n_5271),
.C(n_5253),
.Y(n_5315)
);

INVx1_ASAP7_75t_L g5316 ( 
.A(n_5273),
.Y(n_5316)
);

NOR2xp33_ASAP7_75t_L g5317 ( 
.A(n_5277),
.B(n_5250),
.Y(n_5317)
);

NOR3x2_ASAP7_75t_L g5318 ( 
.A(n_5282),
.B(n_5236),
.C(n_5252),
.Y(n_5318)
);

OAI21xp5_ASAP7_75t_L g5319 ( 
.A1(n_5272),
.A2(n_5222),
.B(n_5241),
.Y(n_5319)
);

AND2x2_ASAP7_75t_L g5320 ( 
.A(n_5285),
.B(n_5263),
.Y(n_5320)
);

OR2x2_ASAP7_75t_L g5321 ( 
.A(n_5293),
.B(n_5242),
.Y(n_5321)
);

NOR3xp33_ASAP7_75t_L g5322 ( 
.A(n_5292),
.B(n_5224),
.C(n_949),
.Y(n_5322)
);

AOI22xp5_ASAP7_75t_L g5323 ( 
.A1(n_5288),
.A2(n_953),
.B1(n_950),
.B2(n_951),
.Y(n_5323)
);

NOR2xp67_ASAP7_75t_L g5324 ( 
.A(n_5323),
.B(n_5297),
.Y(n_5324)
);

AOI221xp5_ASAP7_75t_L g5325 ( 
.A1(n_5309),
.A2(n_5296),
.B1(n_5305),
.B2(n_5299),
.C(n_5301),
.Y(n_5325)
);

AOI22xp5_ASAP7_75t_L g5326 ( 
.A1(n_5312),
.A2(n_5281),
.B1(n_5298),
.B2(n_5303),
.Y(n_5326)
);

NOR2x1_ASAP7_75t_L g5327 ( 
.A(n_5310),
.B(n_5275),
.Y(n_5327)
);

NAND4xp25_ASAP7_75t_L g5328 ( 
.A(n_5316),
.B(n_5304),
.C(n_5284),
.D(n_5295),
.Y(n_5328)
);

NOR2xp67_ASAP7_75t_L g5329 ( 
.A(n_5314),
.B(n_5291),
.Y(n_5329)
);

OAI221xp5_ASAP7_75t_L g5330 ( 
.A1(n_5313),
.A2(n_5308),
.B1(n_5319),
.B2(n_5322),
.C(n_5315),
.Y(n_5330)
);

OR3x1_ASAP7_75t_L g5331 ( 
.A(n_5317),
.B(n_5294),
.C(n_5290),
.Y(n_5331)
);

NOR2x1_ASAP7_75t_L g5332 ( 
.A(n_5320),
.B(n_5302),
.Y(n_5332)
);

INVx1_ASAP7_75t_L g5333 ( 
.A(n_5307),
.Y(n_5333)
);

NOR3xp33_ASAP7_75t_L g5334 ( 
.A(n_5311),
.B(n_5289),
.C(n_5280),
.Y(n_5334)
);

NAND2xp5_ASAP7_75t_L g5335 ( 
.A(n_5332),
.B(n_5321),
.Y(n_5335)
);

NOR2xp33_ASAP7_75t_R g5336 ( 
.A(n_5333),
.B(n_5327),
.Y(n_5336)
);

NAND3xp33_ASAP7_75t_SL g5337 ( 
.A(n_5325),
.B(n_5318),
.C(n_950),
.Y(n_5337)
);

NAND2xp33_ASAP7_75t_SL g5338 ( 
.A(n_5330),
.B(n_954),
.Y(n_5338)
);

NOR2xp33_ASAP7_75t_R g5339 ( 
.A(n_5331),
.B(n_955),
.Y(n_5339)
);

NOR2xp33_ASAP7_75t_R g5340 ( 
.A(n_5328),
.B(n_955),
.Y(n_5340)
);

NAND2xp5_ASAP7_75t_L g5341 ( 
.A(n_5334),
.B(n_957),
.Y(n_5341)
);

OAI22xp5_ASAP7_75t_L g5342 ( 
.A1(n_5335),
.A2(n_5326),
.B1(n_5329),
.B2(n_5324),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_5339),
.Y(n_5343)
);

INVx2_ASAP7_75t_L g5344 ( 
.A(n_5341),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_5336),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_5337),
.Y(n_5346)
);

AO22x2_ASAP7_75t_L g5347 ( 
.A1(n_5342),
.A2(n_5338),
.B1(n_5340),
.B2(n_960),
.Y(n_5347)
);

XNOR2xp5_ASAP7_75t_L g5348 ( 
.A(n_5345),
.B(n_958),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_5347),
.Y(n_5349)
);

NAND2xp5_ASAP7_75t_L g5350 ( 
.A(n_5349),
.B(n_5343),
.Y(n_5350)
);

AOI22xp5_ASAP7_75t_L g5351 ( 
.A1(n_5350),
.A2(n_5346),
.B1(n_5348),
.B2(n_5344),
.Y(n_5351)
);

AOI22x1_ASAP7_75t_L g5352 ( 
.A1(n_5351),
.A2(n_961),
.B1(n_959),
.B2(n_960),
.Y(n_5352)
);

OAI322xp33_ASAP7_75t_L g5353 ( 
.A1(n_5352),
.A2(n_969),
.A3(n_967),
.B1(n_964),
.B2(n_961),
.C1(n_962),
.C2(n_965),
.Y(n_5353)
);

XNOR2xp5_ASAP7_75t_L g5354 ( 
.A(n_5353),
.B(n_962),
.Y(n_5354)
);

NAND2x1_ASAP7_75t_L g5355 ( 
.A(n_5354),
.B(n_964),
.Y(n_5355)
);

AOI22xp33_ASAP7_75t_SL g5356 ( 
.A1(n_5355),
.A2(n_969),
.B1(n_965),
.B2(n_967),
.Y(n_5356)
);

OR2x6_ASAP7_75t_L g5357 ( 
.A(n_5356),
.B(n_970),
.Y(n_5357)
);

AOI21xp5_ASAP7_75t_L g5358 ( 
.A1(n_5357),
.A2(n_970),
.B(n_971),
.Y(n_5358)
);

AOI211xp5_ASAP7_75t_L g5359 ( 
.A1(n_5358),
.A2(n_973),
.B(n_971),
.C(n_972),
.Y(n_5359)
);


endmodule