module fake_jpeg_31043_n_381 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_381);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_381;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_9),
.B(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_20),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_27),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_29),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_67),
.Y(n_124)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_68),
.Y(n_106)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_74),
.Y(n_96)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_41),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_23),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_76),
.B(n_79),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_27),
.B(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_30),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_23),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

BUFx12f_ASAP7_75t_SL g83 ( 
.A(n_29),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_83),
.Y(n_86)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_92),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_102),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_113),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_32),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_70),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_34),
.B1(n_29),
.B2(n_35),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_34),
.B(n_35),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_68),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_70),
.Y(n_142)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_57),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_132),
.Y(n_181)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_86),
.A2(n_63),
.B1(n_73),
.B2(n_78),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_139),
.B1(n_56),
.B2(n_60),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_86),
.A2(n_82),
.B1(n_64),
.B2(n_45),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_154),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_155),
.B1(n_97),
.B2(n_108),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_32),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_148),
.B(n_150),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_94),
.B(n_37),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_28),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_65),
.B1(n_55),
.B2(n_46),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_34),
.B(n_44),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_71),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_111),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_88),
.B(n_43),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_50),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_142),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_175),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_115),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_183),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_169),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_51),
.B1(n_48),
.B2(n_37),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_136),
.B(n_150),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_114),
.B1(n_108),
.B2(n_112),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_177),
.A2(n_163),
.B1(n_169),
.B2(n_165),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_146),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_131),
.B(n_90),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_165),
.A2(n_152),
.B1(n_148),
.B2(n_149),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_185),
.A2(n_192),
.B1(n_172),
.B2(n_167),
.Y(n_222)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_186),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_193),
.B1(n_203),
.B2(n_204),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_188),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_125),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_189),
.B(n_194),
.Y(n_206)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_182),
.B(n_125),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_198),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_165),
.A2(n_145),
.B1(n_134),
.B2(n_157),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_132),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_199),
.B(n_166),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_140),
.B1(n_135),
.B2(n_136),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_201),
.A2(n_170),
.B1(n_180),
.B2(n_174),
.Y(n_209)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_174),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_155),
.B1(n_181),
.B2(n_160),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_181),
.A2(n_135),
.B1(n_114),
.B2(n_129),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_191),
.B(n_160),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_205),
.B(n_133),
.Y(n_236)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_222),
.B1(n_196),
.B2(n_147),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_203),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_218),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_162),
.B1(n_180),
.B2(n_179),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_214),
.A2(n_224),
.B1(n_200),
.B2(n_198),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_162),
.C(n_179),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_128),
.C(n_126),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_162),
.B(n_167),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_202),
.B(n_186),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_189),
.B(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_195),
.B(n_144),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_226),
.Y(n_245)
);

AO22x1_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_157),
.B1(n_171),
.B2(n_151),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_200),
.Y(n_233)
);

AOI32xp33_ASAP7_75t_L g223 ( 
.A1(n_193),
.A2(n_172),
.A3(n_123),
.B1(n_103),
.B2(n_138),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_186),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_133),
.B1(n_126),
.B2(n_128),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_43),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_199),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_229),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_184),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_235),
.B(n_221),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_190),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_241),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_233),
.Y(n_248)
);

AND2x6_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_184),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_103),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_247),
.B1(n_212),
.B2(n_219),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_127),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_243),
.C(n_244),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_188),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_127),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_208),
.A2(n_188),
.B1(n_196),
.B2(n_107),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_228),
.B(n_211),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_258),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_256),
.A2(n_235),
.B1(n_233),
.B2(n_246),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_211),
.Y(n_257)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_240),
.B(n_28),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_216),
.C(n_222),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_267),
.C(n_232),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_221),
.B1(n_224),
.B2(n_212),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_263),
.B1(n_93),
.B2(n_107),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_262),
.B(n_94),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_219),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_266),
.B(n_237),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_217),
.C(n_138),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_255),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_273),
.B(n_264),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_230),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_285),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_252),
.A2(n_233),
.B1(n_217),
.B2(n_40),
.Y(n_277)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_278),
.Y(n_306)
);

AOI22x1_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_112),
.B1(n_48),
.B2(n_104),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_279),
.A2(n_280),
.B1(n_104),
.B2(n_101),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_260),
.A2(n_40),
.B(n_17),
.Y(n_282)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_249),
.A2(n_25),
.B1(n_49),
.B2(n_50),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_94),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_284),
.B(n_288),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_47),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_101),
.B1(n_93),
.B2(n_36),
.Y(n_308)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_294),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_267),
.C(n_248),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_301),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_274),
.B(n_248),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_297),
.Y(n_321)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_259),
.C(n_264),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_288),
.B(n_261),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_304),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_308),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_47),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_285),
.B(n_47),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_278),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_268),
.A2(n_25),
.B1(n_49),
.B2(n_46),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_309),
.A2(n_275),
.B1(n_289),
.B2(n_280),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_317),
.B1(n_326),
.B2(n_300),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_286),
.C(n_281),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_315),
.B(n_320),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_291),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_303),
.A2(n_279),
.B1(n_25),
.B2(n_46),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_290),
.A2(n_47),
.B(n_110),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_318),
.A2(n_292),
.B(n_61),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_23),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_325),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_302),
.Y(n_320)
);

NOR4xp25_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_16),
.C(n_21),
.D(n_19),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_323),
.B(n_21),
.Y(n_328)
);

INVx13_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_324),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_23),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_300),
.A2(n_44),
.B1(n_39),
.B2(n_17),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_334),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_310),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_331),
.B(n_336),
.Y(n_340)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_332),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_333),
.A2(n_337),
.B1(n_338),
.B2(n_51),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_315),
.B(n_299),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_62),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_316),
.A2(n_297),
.B1(n_291),
.B2(n_305),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_314),
.A2(n_19),
.B1(n_1),
.B2(n_2),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_327),
.A2(n_312),
.B(n_324),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_339),
.A2(n_7),
.B(n_8),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_330),
.Y(n_341)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_341),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_331),
.A2(n_314),
.B(n_319),
.Y(n_342)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_342),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_329),
.A2(n_313),
.B1(n_325),
.B2(n_95),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_344),
.B(n_52),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_329),
.A2(n_95),
.B1(n_44),
.B2(n_39),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_345),
.B(n_350),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_346),
.B(n_347),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_336),
.B(n_0),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_332),
.A2(n_0),
.B(n_1),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_349),
.A2(n_4),
.B(n_6),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_341),
.B(n_3),
.Y(n_351)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_351),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_356),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_355),
.B(n_358),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_4),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_343),
.B(n_4),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_357),
.B(n_7),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_360),
.B(n_340),
.C(n_344),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_362),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_363),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_359),
.B(n_8),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_366),
.A2(n_10),
.B(n_12),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_8),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_367),
.B(n_351),
.C(n_353),
.Y(n_369)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_369),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_59),
.C(n_11),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_371),
.A2(n_366),
.B(n_364),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_372),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_375),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_374),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_368),
.C(n_373),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_378),
.A2(n_376),
.B(n_365),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_370),
.C(n_12),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_13),
.Y(n_381)
);


endmodule