module fake_jpeg_22115_n_55 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_55);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_55;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_27),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_26),
.B(n_1),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_30),
.B1(n_29),
.B2(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_17),
.B(n_4),
.Y(n_41)
);

AND2x6_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_40),
.B(n_3),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_48),
.B1(n_7),
.B2(n_9),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_40),
.B(n_8),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_43),
.B1(n_46),
.B2(n_10),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B(n_25),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_11),
.B(n_13),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_14),
.B(n_16),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_18),
.C(n_19),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_55)
);


endmodule