module fake_jpeg_6301_n_190 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_1),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_36),
.Y(n_57)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_2),
.C(n_4),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_2),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_2),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_28),
.B1(n_24),
.B2(n_17),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_44),
.Y(n_66)
);

CKINVDCx9p33_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_30),
.Y(n_76)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2x1_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_16),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_67),
.B(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_58),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_61),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_21),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_21),
.B1(n_29),
.B2(n_27),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_27),
.B1(n_25),
.B2(n_22),
.Y(n_92)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_65),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

OR2x4_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_28),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_69),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_31),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_34),
.B(n_30),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_76),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_80),
.Y(n_97)
);

BUFx4f_ASAP7_75t_SL g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_15),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_38),
.B1(n_28),
.B2(n_24),
.Y(n_84)
);

AO21x2_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_105),
.B(n_58),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_93),
.B(n_89),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_99),
.Y(n_127)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_91),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_106),
.B1(n_63),
.B2(n_52),
.Y(n_119)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_57),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_25),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_66),
.Y(n_107)
);

AO22x1_ASAP7_75t_L g105 ( 
.A1(n_55),
.A2(n_23),
.B1(n_22),
.B2(n_5),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_62),
.B1(n_71),
.B2(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_114),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_61),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_109),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_78),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_78),
.C(n_71),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_123),
.C(n_94),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_23),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_112),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_59),
.Y(n_112)
);

OR2x2_ASAP7_75t_SL g113 ( 
.A(n_105),
.B(n_6),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_113),
.A2(n_118),
.B1(n_125),
.B2(n_91),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_105),
.A3(n_98),
.B1(n_88),
.B2(n_97),
.C1(n_104),
.C2(n_101),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_59),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_124),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_100),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_7),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_94),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_82),
.C(n_86),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_88),
.A2(n_70),
.B(n_63),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_134),
.C(n_119),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_139),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_96),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_85),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_141),
.Y(n_150)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_111),
.B(n_108),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_95),
.B1(n_65),
.B2(n_96),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_146),
.B(n_149),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_109),
.B(n_113),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_116),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_152),
.C(n_130),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_117),
.B(n_111),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_155),
.B(n_129),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_132),
.A2(n_121),
.B(n_115),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_162),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_165),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_129),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_167),
.C(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_137),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_150),
.C(n_146),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_156),
.B1(n_143),
.B2(n_151),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_161),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_175),
.C(n_167),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_172),
.A2(n_158),
.B(n_156),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_164),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_179),
.C(n_170),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g178 ( 
.A(n_173),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_178),
.B(n_180),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_171),
.B(n_165),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_183),
.C(n_170),
.Y(n_185)
);

AO21x1_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_149),
.B(n_135),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_173),
.A3(n_120),
.B1(n_9),
.B2(n_10),
.C1(n_7),
.C2(n_8),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_187),
.C(n_8),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_13),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_133),
.B1(n_9),
.B2(n_10),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_189),
.Y(n_190)
);


endmodule