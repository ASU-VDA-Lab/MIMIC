module fake_jpeg_6957_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NAND2x1_ASAP7_75t_SL g24 ( 
.A(n_11),
.B(n_1),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_20),
.C(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_30),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_24),
.B1(n_15),
.B2(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_13),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_36),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_24),
.B1(n_15),
.B2(n_14),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_16),
.B1(n_19),
.B2(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_41),
.B1(n_40),
.B2(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_20),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g41 ( 
.A1(n_26),
.A2(n_22),
.A3(n_20),
.B1(n_23),
.B2(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_44),
.Y(n_51)
);

CKINVDCx10_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

AND2x6_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_23),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_49),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_57),
.Y(n_62)
);

MAJx2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_29),
.C(n_10),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_56),
.C(n_9),
.Y(n_61)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_29),
.C(n_11),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_46),
.B(n_43),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_61),
.B(n_58),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_11),
.C(n_18),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

AO221x1_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_63),
.B1(n_62),
.B2(n_54),
.C(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_67),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_58),
.C(n_5),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_6),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_4),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_6),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_72),
.B(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_7),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_9),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_8),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_75),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_8),
.Y(n_79)
);


endmodule