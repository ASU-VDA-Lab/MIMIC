module fake_netlist_5_1038_n_111 (n_8, n_10, n_4, n_5, n_7, n_0, n_12, n_9, n_14, n_2, n_16, n_13, n_3, n_11, n_17, n_15, n_6, n_1, n_111);

input n_8;
input n_10;
input n_4;
input n_5;
input n_7;
input n_0;
input n_12;
input n_9;
input n_14;
input n_2;
input n_16;
input n_13;
input n_3;
input n_11;
input n_17;
input n_15;
input n_6;
input n_1;

output n_111;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_108;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_18;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_19;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_109;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVxp67_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_0),
.Y(n_32)
);

CKINVDCx8_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

OA21x2_ASAP7_75t_L g39 ( 
.A1(n_20),
.A2(n_1),
.B(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

AND2x4_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_8),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

AND2x4_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_24),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_25),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

AND2x6_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_R g55 ( 
.A(n_45),
.B(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_R g59 ( 
.A(n_45),
.B(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_44),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_44),
.B1(n_51),
.B2(n_18),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_40),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_51),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_48),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_39),
.B1(n_53),
.B2(n_30),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_43),
.B(n_55),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

AOI211x1_ASAP7_75t_L g77 ( 
.A1(n_75),
.A2(n_32),
.B(n_63),
.C(n_38),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_70),
.B1(n_61),
.B2(n_64),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_74),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_48),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_73),
.Y(n_84)
);

OAI31xp33_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_70),
.A3(n_35),
.B(n_34),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_34),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_72),
.Y(n_88)
);

NOR2x1p5_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_52),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_71),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_72),
.B(n_84),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_72),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_86),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_88),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_88),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_92),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_33),
.B1(n_35),
.B2(n_89),
.Y(n_98)
);

OAI211xp5_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_33),
.B(n_39),
.C(n_49),
.Y(n_99)
);

OAI211xp5_ASAP7_75t_SL g100 ( 
.A1(n_96),
.A2(n_35),
.B(n_3),
.C(n_4),
.Y(n_100)
);

BUFx8_ASAP7_75t_SL g101 ( 
.A(n_98),
.Y(n_101)
);

OAI221xp5_ASAP7_75t_SL g102 ( 
.A1(n_97),
.A2(n_2),
.B1(n_4),
.B2(n_49),
.C(n_39),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_49),
.B(n_39),
.Y(n_103)
);

AO221x1_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_37),
.B1(n_57),
.B2(n_50),
.C(n_15),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_103),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_100),
.C(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_107),
.Y(n_108)
);

NOR2x1p5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_105),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_53),
.B1(n_65),
.B2(n_57),
.Y(n_110)
);

O2A1O1Ixp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_17),
.B(n_65),
.C(n_53),
.Y(n_111)
);


endmodule