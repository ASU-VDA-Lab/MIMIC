module fake_jpeg_19050_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp67_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_43),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_51),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_16),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_30),
.B1(n_22),
.B2(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_32),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_33),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_57),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_41),
.C(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_25),
.B1(n_42),
.B2(n_20),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_25),
.B1(n_42),
.B2(n_20),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_64),
.B1(n_74),
.B2(n_75),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_20),
.B1(n_35),
.B2(n_30),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_44),
.C(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_73),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_23),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_77),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_43),
.B1(n_23),
.B2(n_28),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_27),
.B1(n_33),
.B2(n_31),
.Y(n_121)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_83),
.Y(n_102)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_41),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_47),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_90),
.Y(n_105)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_89),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_55),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_53),
.B1(n_43),
.B2(n_55),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_121),
.B1(n_68),
.B2(n_60),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_119),
.C(n_17),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_47),
.B1(n_54),
.B2(n_39),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_70),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_21),
.B1(n_28),
.B2(n_16),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_69),
.B1(n_83),
.B2(n_80),
.Y(n_130)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_16),
.B(n_39),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_32),
.B(n_18),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_17),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_19),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_58),
.C(n_17),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_32),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_74),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_122),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_123),
.A2(n_133),
.B1(n_135),
.B2(n_146),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_124),
.A2(n_139),
.B(n_142),
.Y(n_180)
);

AOI32xp33_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_65),
.A3(n_82),
.B1(n_77),
.B2(n_72),
.Y(n_125)
);

XOR2x2_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_109),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_71),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_147),
.B1(n_149),
.B2(n_98),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_131),
.B(n_134),
.Y(n_181)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_66),
.B1(n_69),
.B2(n_73),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_96),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_72),
.B1(n_78),
.B2(n_91),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_136),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_138),
.B(n_140),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_32),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_17),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_107),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_32),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_143),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_39),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_148),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_106),
.B(n_109),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_99),
.A2(n_33),
.B1(n_31),
.B2(n_27),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_95),
.A2(n_33),
.B1(n_31),
.B2(n_27),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_95),
.A2(n_31),
.B1(n_27),
.B2(n_18),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_127),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_154),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_158),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_157),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_101),
.CI(n_115),
.CON(n_158),
.SN(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_98),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_166),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_105),
.C(n_113),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_171),
.C(n_17),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_164),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_117),
.B(n_116),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_165),
.A2(n_174),
.B(n_175),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_112),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_168),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_112),
.B1(n_117),
.B2(n_106),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_182),
.B1(n_166),
.B2(n_176),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_116),
.C(n_106),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_114),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_176),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_142),
.A2(n_92),
.B1(n_108),
.B2(n_109),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_143),
.B(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_143),
.B(n_123),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_180),
.B(n_182),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_189),
.A2(n_195),
.B1(n_202),
.B2(n_212),
.Y(n_233)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_149),
.B(n_147),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_196),
.Y(n_222)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_200),
.Y(n_215)
);

AO22x2_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_137),
.B1(n_94),
.B2(n_92),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_181),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_153),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_198),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_132),
.CI(n_18),
.CON(n_198),
.SN(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_103),
.C(n_94),
.Y(n_200)
);

OAI22x1_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_94),
.B1(n_108),
.B2(n_2),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_0),
.B(n_1),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_8),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_211),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_1),
.Y(n_207)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_1),
.B(n_2),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_151),
.B(n_171),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_179),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_213),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_8),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_214),
.B(n_150),
.Y(n_226)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_216),
.B(n_227),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_209),
.A2(n_178),
.B1(n_156),
.B2(n_173),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_221),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_234),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_158),
.B(n_163),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_220),
.B(n_236),
.Y(n_259)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_150),
.B(n_178),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_157),
.B1(n_177),
.B2(n_4),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_186),
.A2(n_3),
.B(n_4),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_199),
.B(n_10),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_237),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_184),
.B(n_10),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_238),
.B(n_211),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_253),
.Y(n_263)
);

NOR2x1_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_200),
.C(n_194),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_243),
.C(n_255),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_184),
.C(n_198),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_205),
.CI(n_198),
.CON(n_245),
.SN(n_245)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_247),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_223),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_217),
.B(n_193),
.CI(n_192),
.CON(n_250),
.SN(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_187),
.C(n_207),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_252),
.A2(n_259),
.B(n_195),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_229),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_187),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_257),
.B(n_188),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_217),
.B(n_222),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_190),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_227),
.C(n_221),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_261),
.B(n_262),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_231),
.C(n_233),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_190),
.C(n_189),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_277),
.C(n_261),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_276),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_246),
.B(n_239),
.Y(n_269)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_244),
.B(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_228),
.B(n_230),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_248),
.B(n_185),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_216),
.B1(n_234),
.B2(n_191),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_273),
.A2(n_249),
.B1(n_251),
.B2(n_256),
.Y(n_279)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_241),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_252),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_275),
.B(n_245),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_255),
.B(n_195),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_191),
.C(n_185),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_276),
.B1(n_265),
.B2(n_277),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_287),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_288),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_254),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_285),
.B(n_289),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_240),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_247),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_291),
.C(n_292),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_195),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_204),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_283),
.A2(n_266),
.B1(n_267),
.B2(n_264),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_296),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_271),
.B(n_204),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_298),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_271),
.B(n_6),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_14),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_5),
.C(n_6),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_301),
.C(n_11),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_7),
.C(n_8),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_11),
.B(n_12),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_302),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_304),
.A2(n_292),
.B1(n_278),
.B2(n_289),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_312),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_278),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_307),
.A2(n_300),
.B(n_294),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_308),
.B(n_311),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_12),
.B(n_13),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_308),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_295),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_316),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_299),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_319),
.Y(n_321)
);

AOI31xp33_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_305),
.A3(n_309),
.B(n_307),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_325),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_317),
.C(n_321),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_294),
.B(n_15),
.Y(n_328)
);


endmodule