module fake_ariane_2609_n_385 (n_83, n_8, n_56, n_60, n_64, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_112, n_45, n_11, n_52, n_73, n_77, n_15, n_93, n_23, n_61, n_108, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_385);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_112;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_93;
input n_23;
input n_61;
input n_108;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_385;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_119;
wire n_124;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_172;
wire n_347;
wire n_183;
wire n_373;
wire n_299;
wire n_133;
wire n_205;
wire n_341;
wire n_245;
wire n_319;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_117;
wire n_139;
wire n_130;
wire n_349;
wire n_346;
wire n_214;
wire n_348;
wire n_379;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_327;
wire n_372;
wire n_377;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_272;
wire n_339;
wire n_167;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_143;
wire n_152;
wire n_120;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_331;
wire n_320;
wire n_267;
wire n_335;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_247;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_248;
wire n_301;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_303;
wire n_168;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_141;
wire n_314;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_333;
wire n_376;
wire n_221;
wire n_321;
wire n_361;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_371;
wire n_199;
wire n_217;
wire n_178;
wire n_308;
wire n_201;
wire n_343;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_249;
wire n_212;
wire n_123;
wire n_355;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_135;
wire n_171;
wire n_384;
wire n_182;
wire n_316;
wire n_196;
wire n_125;
wire n_254;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_216;
wire n_223;
wire n_288;
wire n_179;
wire n_195;
wire n_213;
wire n_304;
wire n_306;
wire n_313;
wire n_203;
wire n_378;
wire n_150;
wire n_375;
wire n_324;
wire n_337;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_342;
wire n_246;
wire n_159;
wire n_358;
wire n_131;
wire n_263;
wire n_360;
wire n_229;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_118;
wire n_121;
wire n_353;
wire n_241;
wire n_357;
wire n_191;
wire n_382;
wire n_211;
wire n_322;
wire n_251;
wire n_351;
wire n_359;
wire n_155;
wire n_127;

BUFx3_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_5),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_3),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_13),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_34),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_3),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_37),
.Y(n_125)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_26),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_71),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_5),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_19),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_20),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_72),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_28),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_86),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_25),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_75),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_48),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_66),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_7),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_87),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_33),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_105),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_35),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_53),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_111),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_45),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_62),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_39),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_10),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_0),
.B(n_52),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_108),
.B(n_69),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_83),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_38),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_15),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_1),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_67),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_2),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_6),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_63),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_80),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_0),
.Y(n_179)
);

BUFx8_ASAP7_75t_SL g180 ( 
.A(n_120),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

CKINVDCx11_ASAP7_75t_R g187 ( 
.A(n_153),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_128),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_132),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_4),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_119),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_123),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_197),
.A2(n_126),
.B1(n_147),
.B2(n_175),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_187),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_126),
.B1(n_124),
.B2(n_172),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_179),
.B(n_159),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_154),
.B1(n_176),
.B2(n_131),
.Y(n_211)
);

NOR2x1p5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_127),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_159),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_196),
.B(n_166),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_160),
.B1(n_143),
.B2(n_171),
.Y(n_218)
);

OR2x6_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_138),
.Y(n_219)
);

AND2x6_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_194),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

NAND2x1p5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_133),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_191),
.B(n_170),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_136),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_R g227 ( 
.A(n_206),
.B(n_145),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_157),
.B1(n_146),
.B2(n_173),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_198),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_198),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_137),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_140),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_156),
.B1(n_150),
.B2(n_155),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_207),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_SL g244 ( 
.A1(n_207),
.A2(n_167),
.B(n_164),
.C(n_163),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_134),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_217),
.A2(n_162),
.B1(n_165),
.B2(n_169),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_151),
.B(n_139),
.C(n_141),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_223),
.B(n_144),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_209),
.A2(n_168),
.B1(n_148),
.B2(n_149),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_177),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_158),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_132),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_224),
.B(n_180),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

AND2x6_ASAP7_75t_SL g258 ( 
.A(n_218),
.B(n_180),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_211),
.A2(n_132),
.B1(n_7),
.B2(n_8),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

AOI21x1_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_202),
.B(n_203),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_SL g262 ( 
.A1(n_245),
.A2(n_220),
.B(n_205),
.C(n_132),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_233),
.B(n_242),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_227),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_246),
.A2(n_218),
.B1(n_200),
.B2(n_219),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_219),
.B(n_210),
.Y(n_266)
);

O2A1O1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_220),
.B(n_8),
.C(n_6),
.Y(n_267)
);

OAI21x1_ASAP7_75t_L g268 ( 
.A1(n_248),
.A2(n_220),
.B(n_11),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_210),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_210),
.B(n_12),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_9),
.B(n_14),
.Y(n_271)
);

NOR3xp33_ASAP7_75t_L g272 ( 
.A(n_233),
.B(n_210),
.C(n_17),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_232),
.A2(n_116),
.B(n_18),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_228),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_242),
.B(n_16),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_21),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_235),
.B(n_22),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_23),
.B(n_24),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_259),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_229),
.B(n_31),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_252),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_251),
.Y(n_283)
);

AOI21xp33_ASAP7_75t_L g284 ( 
.A1(n_243),
.A2(n_240),
.B(n_250),
.Y(n_284)
);

A2O1A1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_259),
.A2(n_32),
.B(n_36),
.C(n_40),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_230),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_286)
);

OA22x2_ASAP7_75t_L g287 ( 
.A1(n_239),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_287)
);

AOI22x1_ASAP7_75t_L g288 ( 
.A1(n_237),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_280),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_283),
.B1(n_265),
.B2(n_284),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_240),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_237),
.Y(n_294)
);

AOI31xp67_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_241),
.A3(n_238),
.B(n_255),
.Y(n_295)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_247),
.C(n_255),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g297 ( 
.A1(n_261),
.A2(n_236),
.B(n_57),
.Y(n_297)
);

AO32x2_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_56),
.A3(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_298)
);

AO32x2_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_61),
.A3(n_64),
.B1(n_68),
.B2(n_76),
.Y(n_299)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_276),
.B(n_256),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_114),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_271),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_273),
.A2(n_77),
.B(n_78),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_262),
.A2(n_81),
.B(n_89),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_273),
.B(n_90),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_285),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_296),
.A2(n_279),
.B(n_278),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_260),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_290),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_296),
.A2(n_278),
.B(n_270),
.Y(n_315)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_288),
.B(n_272),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_110),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_293),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

OA21x2_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_92),
.B(n_94),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_309),
.A2(n_295),
.B(n_308),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_302),
.Y(n_322)
);

AO21x2_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_297),
.B(n_309),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_319),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_293),
.B1(n_300),
.B2(n_305),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_322),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_312),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_299),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_304),
.Y(n_331)
);

OR2x6_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_306),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_325),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_313),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_326),
.Y(n_336)
);

AND2x4_ASAP7_75t_SL g337 ( 
.A(n_331),
.B(n_306),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_331),
.A2(n_311),
.B1(n_299),
.B2(n_321),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_299),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_332),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_298),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_328),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_298),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_336),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_339),
.Y(n_347)
);

AND2x4_ASAP7_75t_SL g348 ( 
.A(n_341),
.B(n_332),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_343),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_333),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_334),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_329),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_335),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_342),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_344),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_329),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_351),
.B(n_335),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_355),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_349),
.Y(n_359)
);

AND2x2_ASAP7_75t_SL g360 ( 
.A(n_348),
.B(n_338),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_341),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_347),
.Y(n_362)
);

NAND4xp25_ASAP7_75t_L g363 ( 
.A(n_359),
.B(n_338),
.C(n_345),
.D(n_346),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_362),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_353),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_359),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_364),
.Y(n_367)
);

AOI221xp5_ASAP7_75t_L g368 ( 
.A1(n_367),
.A2(n_363),
.B1(n_311),
.B2(n_315),
.C(n_355),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_366),
.B(n_352),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_369),
.Y(n_370)
);

OAI21xp33_ASAP7_75t_SL g371 ( 
.A1(n_368),
.A2(n_360),
.B(n_358),
.Y(n_371)
);

AOI322xp5_ASAP7_75t_L g372 ( 
.A1(n_371),
.A2(n_354),
.A3(n_356),
.B1(n_298),
.B2(n_315),
.C1(n_341),
.C2(n_323),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_370),
.B(n_337),
.Y(n_373)
);

NOR3xp33_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_307),
.C(n_361),
.Y(n_374)
);

NOR2x1p5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_372),
.Y(n_375)
);

NAND2xp33_ASAP7_75t_SL g376 ( 
.A(n_375),
.B(n_341),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_376),
.A2(n_332),
.B1(n_323),
.B2(n_348),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_377),
.Y(n_378)
);

AO22x2_ASAP7_75t_L g379 ( 
.A1(n_377),
.A2(n_316),
.B1(n_320),
.B2(n_323),
.Y(n_379)
);

OAI21x1_ASAP7_75t_L g380 ( 
.A1(n_378),
.A2(n_316),
.B(n_320),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_379),
.A2(n_306),
.B1(n_98),
.B2(n_99),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_381),
.A2(n_380),
.B(n_100),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_381),
.B(n_95),
.Y(n_383)
);

OA21x2_ASAP7_75t_L g384 ( 
.A1(n_382),
.A2(n_104),
.B(n_106),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_384),
.A2(n_383),
.B1(n_107),
.B2(n_109),
.Y(n_385)
);


endmodule