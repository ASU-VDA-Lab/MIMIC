module real_aes_9551_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1873;
wire n_1313;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1845;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1872;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_351;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1914;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_733;
wire n_402;
wire n_1404;
wire n_1856;
wire n_658;
wire n_676;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_1102;
wire n_661;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_727;
wire n_1802;
wire n_397;
wire n_1056;
wire n_1083;
wire n_1592;
wire n_1605;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_1457;
wire n_719;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1176;
wire n_640;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1823;
wire n_1547;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1868;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_729;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g377 ( .A1(n_0), .A2(n_168), .B1(n_378), .B2(n_389), .C(n_396), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_0), .A2(n_340), .B1(n_520), .B2(n_523), .C(n_527), .Y(n_519) );
OA22x2_ASAP7_75t_L g1172 ( .A1(n_1), .A2(n_1173), .B1(n_1229), .B2(n_1230), .Y(n_1172) );
INVxp67_ASAP7_75t_SL g1230 ( .A(n_1), .Y(n_1230) );
AOI22xp5_ASAP7_75t_L g1610 ( .A1(n_2), .A2(n_331), .B1(n_1585), .B2(n_1589), .Y(n_1610) );
CKINVDCx5p33_ASAP7_75t_R g1043 ( .A(n_3), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_4), .Y(n_1044) );
INVxp33_ASAP7_75t_L g1330 ( .A(n_5), .Y(n_1330) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_5), .A2(n_93), .B1(n_919), .B2(n_1384), .Y(n_1392) );
AOI221xp5_ASAP7_75t_L g1031 ( .A1(n_6), .A2(n_90), .B1(n_839), .B2(n_1032), .C(n_1034), .Y(n_1031) );
INVx1_ASAP7_75t_L g1051 ( .A(n_6), .Y(n_1051) );
AOI22xp33_ASAP7_75t_SL g916 ( .A1(n_7), .A2(n_152), .B1(n_917), .B2(n_919), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_7), .A2(n_57), .B1(n_835), .B2(n_949), .Y(n_948) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_8), .A2(n_260), .B1(n_728), .B2(n_730), .C(n_731), .Y(n_727) );
INVx1_ASAP7_75t_L g788 ( .A(n_8), .Y(n_788) );
INVx1_ASAP7_75t_L g1421 ( .A(n_9), .Y(n_1421) );
OAI22xp5_ASAP7_75t_L g1467 ( .A1(n_10), .A2(n_61), .B1(n_1132), .B2(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g1485 ( .A(n_10), .Y(n_1485) );
XNOR2x2_ASAP7_75t_L g909 ( .A(n_11), .B(n_910), .Y(n_909) );
CKINVDCx5p33_ASAP7_75t_R g675 ( .A(n_12), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g1611 ( .A1(n_13), .A2(n_282), .B1(n_1556), .B2(n_1602), .Y(n_1611) );
AOI22xp33_ASAP7_75t_SL g921 ( .A1(n_14), .A2(n_57), .B1(n_922), .B2(n_923), .Y(n_921) );
AOI21xp33_ASAP7_75t_L g951 ( .A1(n_14), .A2(n_546), .B(n_952), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_15), .A2(n_235), .B1(n_1176), .B2(n_1177), .Y(n_1175) );
CKINVDCx5p33_ASAP7_75t_R g1225 ( .A(n_15), .Y(n_1225) );
CKINVDCx5p33_ASAP7_75t_R g1137 ( .A(n_16), .Y(n_1137) );
INVxp67_ASAP7_75t_L g587 ( .A(n_17), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_17), .A2(n_59), .B1(n_629), .B2(n_630), .C(n_631), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g1411 ( .A1(n_18), .A2(n_286), .B1(n_858), .B2(n_1407), .Y(n_1411) );
INVxp67_ASAP7_75t_SL g1446 ( .A(n_18), .Y(n_1446) );
CKINVDCx16_ASAP7_75t_R g1627 ( .A(n_19), .Y(n_1627) );
INVxp33_ASAP7_75t_L g1332 ( .A(n_20), .Y(n_1332) );
AOI22xp33_ASAP7_75t_L g1391 ( .A1(n_20), .A2(n_200), .B1(n_1292), .B2(n_1386), .Y(n_1391) );
OAI221xp5_ASAP7_75t_L g1084 ( .A1(n_21), .A2(n_66), .B1(n_1085), .B2(n_1087), .C(n_1088), .Y(n_1084) );
INVx1_ASAP7_75t_L g1117 ( .A(n_21), .Y(n_1117) );
INVx1_ASAP7_75t_L g939 ( .A(n_22), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_22), .A2(n_293), .B1(n_949), .B2(n_952), .Y(n_956) );
AOI221xp5_ASAP7_75t_L g1452 ( .A1(n_23), .A2(n_334), .B1(n_874), .B2(n_1453), .C(n_1455), .Y(n_1452) );
INVx1_ASAP7_75t_L g1477 ( .A(n_23), .Y(n_1477) );
CKINVDCx5p33_ASAP7_75t_R g1254 ( .A(n_24), .Y(n_1254) );
XNOR2xp5_ASAP7_75t_L g1797 ( .A(n_25), .B(n_1798), .Y(n_1797) );
OAI22xp5_ASAP7_75t_L g1510 ( .A1(n_26), .A2(n_329), .B1(n_682), .B2(n_1511), .Y(n_1510) );
INVxp67_ASAP7_75t_SL g1548 ( .A(n_26), .Y(n_1548) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_27), .A2(n_342), .B1(n_624), .B2(n_683), .Y(n_726) );
INVx1_ASAP7_75t_L g760 ( .A(n_27), .Y(n_760) );
OAI221xp5_ASAP7_75t_L g581 ( .A1(n_28), .A2(n_121), .B1(n_582), .B2(n_583), .C(n_584), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_28), .A2(n_121), .B1(n_624), .B2(n_625), .Y(n_623) );
INVxp67_ASAP7_75t_SL g809 ( .A(n_29), .Y(n_809) );
AOI221xp5_ASAP7_75t_L g831 ( .A1(n_29), .A2(n_323), .B1(n_520), .B2(n_631), .C(n_829), .Y(n_831) );
AOI221xp5_ASAP7_75t_L g1039 ( .A1(n_30), .A2(n_225), .B1(n_630), .B2(n_631), .C(n_1040), .Y(n_1039) );
INVx1_ASAP7_75t_L g1063 ( .A(n_30), .Y(n_1063) );
CKINVDCx5p33_ASAP7_75t_R g644 ( .A(n_31), .Y(n_644) );
OAI211xp5_ASAP7_75t_SL g1404 ( .A1(n_32), .A2(n_565), .B(n_1405), .C(n_1414), .Y(n_1404) );
AOI221xp5_ASAP7_75t_L g1439 ( .A1(n_32), .A2(n_188), .B1(n_923), .B2(n_1440), .C(n_1442), .Y(n_1439) );
INVx1_ASAP7_75t_L g1103 ( .A(n_33), .Y(n_1103) );
INVx1_ASAP7_75t_L g350 ( .A(n_34), .Y(n_350) );
INVx1_ASAP7_75t_L g739 ( .A(n_35), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_35), .A2(n_308), .B1(n_778), .B2(n_780), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g1298 ( .A(n_36), .Y(n_1298) );
AOI22xp5_ASAP7_75t_L g1606 ( .A1(n_37), .A2(n_156), .B1(n_1585), .B2(n_1589), .Y(n_1606) );
INVx1_ASAP7_75t_L g647 ( .A(n_38), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_38), .A2(n_179), .B1(n_686), .B2(n_688), .C(n_690), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g1181 ( .A1(n_39), .A2(n_67), .B1(n_411), .B2(n_421), .C(n_980), .Y(n_1181) );
OAI222xp33_ASAP7_75t_L g1209 ( .A1(n_39), .A2(n_67), .B1(n_220), .B2(n_502), .C1(n_507), .C2(n_876), .Y(n_1209) );
AOI22xp33_ASAP7_75t_L g1591 ( .A1(n_40), .A2(n_216), .B1(n_1554), .B2(n_1562), .Y(n_1591) );
AOI21xp33_ASAP7_75t_L g1146 ( .A1(n_41), .A2(n_702), .B(n_1147), .Y(n_1146) );
AOI221xp5_ASAP7_75t_L g1167 ( .A1(n_41), .A2(n_83), .B1(n_380), .B2(n_438), .C(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1515 ( .A(n_42), .Y(n_1515) );
OAI221xp5_ASAP7_75t_L g1531 ( .A1(n_42), .A2(n_288), .B1(n_378), .B2(n_1532), .C(n_1533), .Y(n_1531) );
INVx1_ASAP7_75t_L g1862 ( .A(n_43), .Y(n_1862) );
AOI22xp33_ASAP7_75t_L g1899 ( .A1(n_43), .A2(n_213), .B1(n_769), .B2(n_1900), .Y(n_1899) );
AOI22xp33_ASAP7_75t_L g1895 ( .A1(n_44), .A2(n_147), .B1(n_769), .B2(n_917), .Y(n_1895) );
AOI22xp33_ASAP7_75t_L g1903 ( .A1(n_44), .A2(n_147), .B1(n_550), .B2(n_1257), .Y(n_1903) );
AOI22xp33_ASAP7_75t_SL g1406 ( .A1(n_45), .A2(n_101), .B1(n_634), .B2(n_1407), .Y(n_1406) );
AOI22xp33_ASAP7_75t_SL g1427 ( .A1(n_45), .A2(n_174), .B1(n_773), .B2(n_1428), .Y(n_1427) );
INVx1_ASAP7_75t_L g750 ( .A(n_46), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_46), .A2(n_316), .B1(n_773), .B2(n_775), .Y(n_774) );
AOI221xp5_ASAP7_75t_L g1412 ( .A1(n_47), .A2(n_196), .B1(n_618), .B2(n_634), .C(n_1413), .Y(n_1412) );
OAI21xp33_ASAP7_75t_SL g1425 ( .A1(n_47), .A2(n_1177), .B(n_1426), .Y(n_1425) );
OAI222xp33_ASAP7_75t_L g868 ( .A1(n_48), .A2(n_172), .B1(n_265), .B2(n_869), .C1(n_871), .C2(n_873), .Y(n_868) );
AOI221xp5_ASAP7_75t_L g903 ( .A1(n_48), .A2(n_172), .B1(n_904), .B2(n_906), .C(n_907), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g1600 ( .A1(n_49), .A2(n_125), .B1(n_1585), .B2(n_1589), .Y(n_1600) );
AO221x2_ASAP7_75t_L g1612 ( .A1(n_50), .A2(n_243), .B1(n_1556), .B2(n_1602), .C(n_1613), .Y(n_1612) );
CKINVDCx16_ASAP7_75t_R g1501 ( .A(n_51), .Y(n_1501) );
CKINVDCx5p33_ASAP7_75t_R g914 ( .A(n_52), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g1465 ( .A(n_53), .Y(n_1465) );
AOI22xp5_ASAP7_75t_SL g1595 ( .A1(n_54), .A2(n_232), .B1(n_1556), .B2(n_1562), .Y(n_1595) );
INVxp67_ASAP7_75t_SL g808 ( .A(n_55), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_55), .A2(n_207), .B1(n_621), .B2(n_833), .Y(n_832) );
OAI221xp5_ASAP7_75t_L g410 ( .A1(n_56), .A2(n_108), .B1(n_411), .B2(n_420), .C(n_425), .Y(n_410) );
OAI221xp5_ASAP7_75t_SL g501 ( .A1(n_56), .A2(n_108), .B1(n_502), .B2(n_507), .C(n_512), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g1191 ( .A(n_58), .Y(n_1191) );
INVxp33_ASAP7_75t_L g598 ( .A(n_59), .Y(n_598) );
INVxp67_ASAP7_75t_L g968 ( .A(n_60), .Y(n_968) );
INVx1_ASAP7_75t_L g1487 ( .A(n_61), .Y(n_1487) );
CKINVDCx14_ASAP7_75t_R g1572 ( .A(n_62), .Y(n_1572) );
AOI22xp33_ASAP7_75t_L g1524 ( .A1(n_63), .A2(n_201), .B1(n_549), .B2(n_1513), .Y(n_1524) );
AOI22xp33_ASAP7_75t_L g1540 ( .A1(n_63), .A2(n_201), .B1(n_778), .B2(n_1428), .Y(n_1540) );
OAI221xp5_ASAP7_75t_L g1139 ( .A1(n_64), .A2(n_138), .B1(n_1135), .B2(n_1140), .C(n_1141), .Y(n_1139) );
INVx1_ASAP7_75t_L g1171 ( .A(n_64), .Y(n_1171) );
INVxp67_ASAP7_75t_L g992 ( .A(n_65), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_65), .A2(n_98), .B1(n_838), .B2(n_1017), .Y(n_1016) );
AOI221xp5_ASAP7_75t_L g1114 ( .A1(n_66), .A2(n_202), .B1(n_895), .B2(n_1115), .C(n_1116), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1893 ( .A1(n_68), .A2(n_195), .B1(n_895), .B2(n_1894), .Y(n_1893) );
AOI22xp33_ASAP7_75t_L g1902 ( .A1(n_68), .A2(n_195), .B1(n_621), .B2(n_872), .Y(n_1902) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_69), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g1189 ( .A(n_70), .Y(n_1189) );
AOI21xp33_ASAP7_75t_L g1809 ( .A1(n_71), .A2(n_618), .B(n_735), .Y(n_1809) );
INVxp33_ASAP7_75t_L g1831 ( .A(n_71), .Y(n_1831) );
OAI22xp33_ASAP7_75t_L g1037 ( .A1(n_72), .A2(n_208), .B1(n_845), .B2(n_1012), .Y(n_1037) );
OAI221xp5_ASAP7_75t_L g1055 ( .A1(n_72), .A2(n_208), .B1(n_421), .B2(n_584), .C(n_1056), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1584 ( .A1(n_73), .A2(n_205), .B1(n_1585), .B2(n_1588), .Y(n_1584) );
INVx1_ASAP7_75t_L g997 ( .A(n_74), .Y(n_997) );
AOI22x1_ASAP7_75t_L g1401 ( .A1(n_75), .A2(n_1402), .B1(n_1447), .B2(n_1448), .Y(n_1401) );
INVxp67_ASAP7_75t_L g1447 ( .A(n_75), .Y(n_1447) );
XNOR2x2_ASAP7_75t_L g1449 ( .A(n_76), .B(n_1450), .Y(n_1449) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_77), .A2(n_261), .B1(n_1255), .B2(n_1371), .Y(n_1370) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_77), .A2(n_261), .B1(n_919), .B2(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1863 ( .A(n_78), .Y(n_1863) );
AOI22xp33_ASAP7_75t_L g1897 ( .A1(n_78), .A2(n_167), .B1(n_895), .B2(n_1898), .Y(n_1897) );
CKINVDCx20_ASAP7_75t_R g1803 ( .A(n_79), .Y(n_1803) );
CKINVDCx5p33_ASAP7_75t_R g936 ( .A(n_80), .Y(n_936) );
INVxp33_ASAP7_75t_L g580 ( .A(n_81), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_81), .A2(n_343), .B1(n_620), .B2(n_621), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_82), .A2(n_175), .B1(n_438), .B2(n_926), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g962 ( .A1(n_82), .A2(n_175), .B1(n_963), .B2(n_964), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_83), .A2(n_230), .B1(n_708), .B2(n_949), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_84), .A2(n_176), .B1(n_730), .B2(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1124 ( .A(n_84), .Y(n_1124) );
INVxp33_ASAP7_75t_SL g1528 ( .A(n_85), .Y(n_1528) );
AOI22xp33_ASAP7_75t_L g1544 ( .A1(n_85), .A2(n_327), .B1(n_1428), .B2(n_1542), .Y(n_1544) );
OAI221xp5_ASAP7_75t_L g649 ( .A1(n_86), .A2(n_157), .B1(n_411), .B2(n_583), .C(n_650), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_86), .A2(n_157), .B1(n_682), .B2(n_683), .Y(n_681) );
CKINVDCx14_ASAP7_75t_R g1614 ( .A(n_87), .Y(n_1614) );
INVx1_ASAP7_75t_L g846 ( .A(n_88), .Y(n_846) );
INVx1_ASAP7_75t_L g386 ( .A(n_89), .Y(n_386) );
OR2x2_ASAP7_75t_L g418 ( .A(n_89), .B(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_L g431 ( .A(n_89), .Y(n_431) );
BUFx2_ASAP7_75t_L g479 ( .A(n_89), .Y(n_479) );
INVx1_ASAP7_75t_L g1053 ( .A(n_90), .Y(n_1053) );
AOI221xp5_ASAP7_75t_L g1293 ( .A1(n_91), .A2(n_291), .B1(n_400), .B2(n_429), .C(n_919), .Y(n_1293) );
INVx1_ASAP7_75t_L g1316 ( .A(n_91), .Y(n_1316) );
AOI22xp33_ASAP7_75t_SL g927 ( .A1(n_92), .A2(n_106), .B1(n_917), .B2(n_919), .Y(n_927) );
INVx1_ASAP7_75t_L g961 ( .A(n_92), .Y(n_961) );
INVxp67_ASAP7_75t_L g1337 ( .A(n_93), .Y(n_1337) );
CKINVDCx5p33_ASAP7_75t_R g1800 ( .A(n_94), .Y(n_1800) );
AOI221xp5_ASAP7_75t_L g1812 ( .A1(n_95), .A2(n_223), .B1(n_1813), .B2(n_1815), .C(n_1818), .Y(n_1812) );
INVxp67_ASAP7_75t_SL g1839 ( .A(n_95), .Y(n_1839) );
AOI221xp5_ASAP7_75t_SL g1095 ( .A1(n_96), .A2(n_103), .B1(n_550), .B2(n_618), .C(n_855), .Y(n_1095) );
INVx1_ASAP7_75t_L g1112 ( .A(n_96), .Y(n_1112) );
INVxp33_ASAP7_75t_L g1363 ( .A(n_97), .Y(n_1363) );
AOI22xp33_ASAP7_75t_L g1375 ( .A1(n_97), .A2(n_295), .B1(n_617), .B2(n_1371), .Y(n_1375) );
INVxp33_ASAP7_75t_L g983 ( .A(n_98), .Y(n_983) );
INVx1_ASAP7_75t_L g1090 ( .A(n_99), .Y(n_1090) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_100), .A2(n_638), .B1(n_714), .B2(n_715), .Y(n_637) );
INVx1_ASAP7_75t_L g714 ( .A(n_100), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_101), .A2(n_115), .B1(n_779), .B2(n_1430), .Y(n_1429) );
INVx1_ASAP7_75t_L g455 ( .A(n_102), .Y(n_455) );
INVx1_ASAP7_75t_L g1111 ( .A(n_103), .Y(n_1111) );
XOR2x2_ASAP7_75t_L g1127 ( .A(n_104), .B(n_1128), .Y(n_1127) );
CKINVDCx5p33_ASAP7_75t_R g1303 ( .A(n_105), .Y(n_1303) );
NOR2xp33_ASAP7_75t_L g942 ( .A(n_106), .B(n_560), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g1178 ( .A1(n_107), .A2(n_220), .B1(n_476), .B2(n_1179), .Y(n_1178) );
CKINVDCx5p33_ASAP7_75t_R g1223 ( .A(n_107), .Y(n_1223) );
INVxp33_ASAP7_75t_L g1356 ( .A(n_109), .Y(n_1356) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_109), .A2(n_272), .B1(n_860), .B2(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1004 ( .A(n_110), .Y(n_1004) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_111), .Y(n_491) );
INVxp67_ASAP7_75t_L g978 ( .A(n_112), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_112), .A2(n_145), .B1(n_730), .B2(n_872), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_113), .A2(n_255), .B1(n_622), .B2(n_952), .Y(n_1154) );
OAI211xp5_ASAP7_75t_L g1156 ( .A1(n_113), .A2(n_1157), .B(n_1158), .C(n_1160), .Y(n_1156) );
INVx1_ASAP7_75t_L g1249 ( .A(n_114), .Y(n_1249) );
AOI221xp5_ASAP7_75t_L g1280 ( .A1(n_114), .A2(n_133), .B1(n_380), .B2(n_923), .C(n_1281), .Y(n_1280) );
AOI221xp5_ASAP7_75t_L g1409 ( .A1(n_115), .A2(n_174), .B1(n_520), .B2(n_741), .C(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g1020 ( .A(n_116), .Y(n_1020) );
OAI22xp33_ASAP7_75t_SL g1469 ( .A1(n_117), .A2(n_151), .B1(n_732), .B2(n_1133), .Y(n_1469) );
INVx1_ASAP7_75t_L g1488 ( .A(n_117), .Y(n_1488) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_118), .Y(n_1030) );
AOI221xp5_ASAP7_75t_L g1099 ( .A1(n_119), .A2(n_184), .B1(n_520), .B2(n_629), .C(n_631), .Y(n_1099) );
AOI221xp5_ASAP7_75t_L g1119 ( .A1(n_119), .A2(n_176), .B1(n_1120), .B2(n_1121), .C(n_1123), .Y(n_1119) );
XNOR2x1_ASAP7_75t_L g571 ( .A(n_120), .B(n_572), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g1462 ( .A(n_122), .Y(n_1462) );
CKINVDCx5p33_ASAP7_75t_R g674 ( .A(n_123), .Y(n_674) );
OAI222xp33_ASAP7_75t_L g875 ( .A1(n_124), .A2(n_192), .B1(n_324), .B2(n_845), .C1(n_876), .C2(n_877), .Y(n_875) );
INVx1_ASAP7_75t_L g888 ( .A(n_124), .Y(n_888) );
AOI221xp5_ASAP7_75t_L g740 ( .A1(n_126), .A2(n_300), .B1(n_546), .B2(n_741), .C(n_744), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_126), .A2(n_214), .B1(n_673), .B2(n_773), .Y(n_772) );
OAI22xp33_ASAP7_75t_L g1134 ( .A1(n_127), .A2(n_304), .B1(n_515), .B2(n_1135), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_127), .A2(n_183), .B1(n_767), .B2(n_781), .Y(n_1166) );
INVx1_ASAP7_75t_L g1884 ( .A(n_128), .Y(n_1884) );
AOI22xp33_ASAP7_75t_SL g1908 ( .A1(n_128), .A2(n_297), .B1(n_1101), .B2(n_1257), .Y(n_1908) );
INVxp67_ASAP7_75t_L g977 ( .A(n_129), .Y(n_977) );
AOI221xp5_ASAP7_75t_L g1009 ( .A1(n_129), .A2(n_189), .B1(n_617), .B2(n_618), .C(n_735), .Y(n_1009) );
AOI21xp5_ASAP7_75t_L g1155 ( .A1(n_130), .A2(n_838), .B(n_839), .Y(n_1155) );
INVx1_ASAP7_75t_L g1161 ( .A(n_130), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_131), .A2(n_183), .B1(n_1132), .B2(n_1133), .Y(n_1131) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_131), .A2(n_304), .B1(n_407), .B2(n_922), .Y(n_1165) );
CKINVDCx5p33_ASAP7_75t_R g1027 ( .A(n_132), .Y(n_1027) );
INVx1_ASAP7_75t_L g1269 ( .A(n_133), .Y(n_1269) );
OAI221xp5_ASAP7_75t_L g802 ( .A1(n_134), .A2(n_170), .B1(n_422), .B2(n_582), .C(n_584), .Y(n_802) );
OAI22xp33_ASAP7_75t_L g842 ( .A1(n_134), .A2(n_170), .B1(n_843), .B2(n_845), .Y(n_842) );
AOI221xp5_ASAP7_75t_L g1522 ( .A1(n_135), .A2(n_296), .B1(n_629), .B2(n_1410), .C(n_1523), .Y(n_1522) );
AOI22xp33_ASAP7_75t_L g1541 ( .A1(n_135), .A2(n_296), .B1(n_1542), .B2(n_1543), .Y(n_1541) );
CKINVDCx5p33_ASAP7_75t_R g1144 ( .A(n_136), .Y(n_1144) );
OAI221xp5_ASAP7_75t_L g979 ( .A1(n_137), .A2(n_178), .B1(n_411), .B2(n_421), .C(n_980), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g1011 ( .A1(n_137), .A2(n_178), .B1(n_625), .B2(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1159 ( .A(n_138), .Y(n_1159) );
INVx1_ASAP7_75t_L g1093 ( .A(n_139), .Y(n_1093) );
AOI22xp5_ASAP7_75t_SL g1594 ( .A1(n_140), .A2(n_162), .B1(n_1585), .B2(n_1589), .Y(n_1594) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_141), .A2(n_294), .B1(n_546), .B2(n_630), .C(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g902 ( .A(n_141), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g1194 ( .A(n_142), .Y(n_1194) );
INVx1_ASAP7_75t_L g374 ( .A(n_143), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_144), .Y(n_678) );
INVxp67_ASAP7_75t_L g973 ( .A(n_145), .Y(n_973) );
INVx1_ASAP7_75t_L g1339 ( .A(n_146), .Y(n_1339) );
OAI22xp5_ASAP7_75t_L g1349 ( .A1(n_146), .A2(n_281), .B1(n_1350), .B2(n_1352), .Y(n_1349) );
INVx1_ASAP7_75t_L g603 ( .A(n_148), .Y(n_603) );
INVxp33_ASAP7_75t_SL g1527 ( .A(n_149), .Y(n_1527) );
AOI22xp33_ASAP7_75t_L g1545 ( .A1(n_149), .A2(n_277), .B1(n_778), .B2(n_1543), .Y(n_1545) );
INVx1_ASAP7_75t_L g1560 ( .A(n_150), .Y(n_1560) );
INVx1_ASAP7_75t_L g1483 ( .A(n_151), .Y(n_1483) );
INVx1_ASAP7_75t_L g945 ( .A(n_152), .Y(n_945) );
INVx1_ASAP7_75t_L g1877 ( .A(n_153), .Y(n_1877) );
AOI22xp33_ASAP7_75t_L g1909 ( .A1(n_153), .A2(n_194), .B1(n_621), .B2(n_1910), .Y(n_1909) );
INVx1_ASAP7_75t_L g458 ( .A(n_154), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g1624 ( .A(n_155), .Y(n_1624) );
INVx1_ASAP7_75t_L g607 ( .A(n_158), .Y(n_607) );
INVx1_ASAP7_75t_L g1558 ( .A(n_159), .Y(n_1558) );
NAND2xp5_ASAP7_75t_L g1577 ( .A(n_159), .B(n_1571), .Y(n_1577) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_160), .A2(n_237), .B1(n_688), .B2(n_1097), .Y(n_1096) );
OAI221xp5_ASAP7_75t_L g1108 ( .A1(n_160), .A2(n_237), .B1(n_437), .B2(n_1109), .C(n_1110), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_161), .A2(n_214), .B1(n_523), .B2(n_747), .Y(n_746) );
AOI22xp33_ASAP7_75t_SL g766 ( .A1(n_161), .A2(n_300), .B1(n_767), .B2(n_769), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_163), .A2(n_697), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g787 ( .A(n_163), .Y(n_787) );
INVx2_ASAP7_75t_L g362 ( .A(n_164), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g1245 ( .A(n_165), .Y(n_1245) );
OAI22x1_ASAP7_75t_SL g1326 ( .A1(n_166), .A2(n_1327), .B1(n_1393), .B2(n_1394), .Y(n_1326) );
INVx1_ASAP7_75t_L g1393 ( .A(n_166), .Y(n_1393) );
INVx1_ASAP7_75t_L g1866 ( .A(n_167), .Y(n_1866) );
INVx1_ASAP7_75t_L g514 ( .A(n_168), .Y(n_514) );
BUFx3_ASAP7_75t_L g488 ( .A(n_169), .Y(n_488) );
INVx1_ASAP7_75t_L g518 ( .A(n_169), .Y(n_518) );
INVx1_ASAP7_75t_L g1415 ( .A(n_171), .Y(n_1415) );
INVx1_ASAP7_75t_L g653 ( .A(n_173), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_173), .A2(n_280), .B1(n_551), .B2(n_707), .Y(n_706) );
INVxp33_ASAP7_75t_L g800 ( .A(n_177), .Y(n_800) );
AOI221xp5_ASAP7_75t_L g837 ( .A1(n_177), .A2(n_219), .B1(n_630), .B2(n_838), .C(n_839), .Y(n_837) );
INVx1_ASAP7_75t_L g642 ( .A(n_179), .Y(n_642) );
CKINVDCx5p33_ASAP7_75t_R g1461 ( .A(n_180), .Y(n_1461) );
OAI221xp5_ASAP7_75t_L g1867 ( .A1(n_181), .A2(n_239), .B1(n_1868), .B2(n_1871), .C(n_1872), .Y(n_1867) );
INVx1_ASAP7_75t_L g1880 ( .A(n_181), .Y(n_1880) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_182), .A2(n_309), .B1(n_922), .B2(n_1292), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_182), .A2(n_309), .B1(n_1036), .B2(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1125 ( .A(n_184), .Y(n_1125) );
INVxp67_ASAP7_75t_L g433 ( .A(n_185), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_185), .A2(n_315), .B1(n_549), .B2(n_551), .Y(n_548) );
OAI221xp5_ASAP7_75t_SL g1804 ( .A1(n_186), .A2(n_330), .B1(n_843), .B2(n_1511), .C(n_1805), .Y(n_1804) );
OAI221xp5_ASAP7_75t_L g1833 ( .A1(n_186), .A2(n_330), .B1(n_411), .B2(n_422), .C(n_650), .Y(n_1833) );
INVx1_ASAP7_75t_L g403 ( .A(n_187), .Y(n_403) );
INVxp67_ASAP7_75t_SL g1416 ( .A(n_188), .Y(n_1416) );
INVxp67_ASAP7_75t_L g974 ( .A(n_189), .Y(n_974) );
INVx1_ASAP7_75t_L g1091 ( .A(n_190), .Y(n_1091) );
CKINVDCx5p33_ASAP7_75t_R g1192 ( .A(n_191), .Y(n_1192) );
INVx1_ASAP7_75t_L g882 ( .A(n_192), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_193), .A2(n_284), .B1(n_747), .B2(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g887 ( .A(n_193), .Y(n_887) );
INVx1_ASAP7_75t_L g1878 ( .A(n_194), .Y(n_1878) );
INVxp33_ASAP7_75t_SL g1435 ( .A(n_196), .Y(n_1435) );
INVxp67_ASAP7_75t_L g596 ( .A(n_197), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_197), .A2(n_254), .B1(n_621), .B2(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g1824 ( .A(n_198), .Y(n_1824) );
INVx1_ASAP7_75t_L g483 ( .A(n_199), .Y(n_483) );
INVx1_ASAP7_75t_L g531 ( .A(n_199), .Y(n_531) );
INVxp33_ASAP7_75t_L g1335 ( .A(n_200), .Y(n_1335) );
INVx1_ASAP7_75t_L g1089 ( .A(n_202), .Y(n_1089) );
INVxp33_ASAP7_75t_SL g797 ( .A(n_203), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_203), .A2(n_209), .B1(n_629), .B2(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g1258 ( .A(n_204), .Y(n_1258) );
OAI221xp5_ASAP7_75t_L g1286 ( .A1(n_204), .A2(n_228), .B1(n_1287), .B2(n_1289), .C(n_1290), .Y(n_1286) );
CKINVDCx20_ASAP7_75t_R g1565 ( .A(n_206), .Y(n_1565) );
INVx1_ASAP7_75t_L g815 ( .A(n_207), .Y(n_815) );
INVxp33_ASAP7_75t_SL g801 ( .A(n_209), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g1151 ( .A(n_210), .Y(n_1151) );
AOI221xp5_ASAP7_75t_L g1459 ( .A1(n_211), .A2(n_307), .B1(n_702), .B2(n_1036), .C(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1492 ( .A(n_211), .Y(n_1492) );
INVx1_ASAP7_75t_L g600 ( .A(n_212), .Y(n_600) );
INVx1_ASAP7_75t_L g1873 ( .A(n_213), .Y(n_1873) );
INVx1_ASAP7_75t_L g790 ( .A(n_215), .Y(n_790) );
AOI221xp5_ASAP7_75t_L g854 ( .A1(n_217), .A2(n_301), .B1(n_550), .B2(n_618), .C(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g885 ( .A(n_217), .Y(n_885) );
CKINVDCx14_ASAP7_75t_R g1615 ( .A(n_218), .Y(n_1615) );
INVxp33_ASAP7_75t_L g798 ( .A(n_219), .Y(n_798) );
INVx1_ASAP7_75t_L g611 ( .A(n_221), .Y(n_611) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_222), .Y(n_913) );
INVx1_ASAP7_75t_L g1837 ( .A(n_223), .Y(n_1837) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_224), .A2(n_231), .B1(n_741), .B2(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1049 ( .A(n_224), .Y(n_1049) );
INVx1_ASAP7_75t_L g1065 ( .A(n_225), .Y(n_1065) );
INVxp67_ASAP7_75t_L g989 ( .A(n_226), .Y(n_989) );
AOI221xp5_ASAP7_75t_L g1014 ( .A1(n_226), .A2(n_238), .B1(n_539), .B2(n_705), .C(n_1015), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1820 ( .A1(n_227), .A2(n_290), .B1(n_874), .B2(n_1821), .Y(n_1820) );
INVx1_ASAP7_75t_L g1836 ( .A(n_227), .Y(n_1836) );
INVx1_ASAP7_75t_L g1263 ( .A(n_228), .Y(n_1263) );
CKINVDCx5p33_ASAP7_75t_R g1865 ( .A(n_229), .Y(n_1865) );
INVx1_ASAP7_75t_L g1169 ( .A(n_230), .Y(n_1169) );
INVx1_ASAP7_75t_L g1054 ( .A(n_231), .Y(n_1054) );
XNOR2xp5_ASAP7_75t_L g1021 ( .A(n_232), .B(n_1022), .Y(n_1021) );
OAI211xp5_ASAP7_75t_SL g1417 ( .A1(n_233), .A2(n_1418), .B(n_1419), .C(n_1423), .Y(n_1417) );
INVx1_ASAP7_75t_L g1444 ( .A(n_233), .Y(n_1444) );
INVx1_ASAP7_75t_L g940 ( .A(n_234), .Y(n_940) );
OAI211xp5_ASAP7_75t_L g959 ( .A1(n_234), .A2(n_876), .B(n_960), .C(n_965), .Y(n_959) );
CKINVDCx5p33_ASAP7_75t_R g1221 ( .A(n_235), .Y(n_1221) );
CKINVDCx5p33_ASAP7_75t_R g1195 ( .A(n_236), .Y(n_1195) );
INVxp33_ASAP7_75t_L g986 ( .A(n_238), .Y(n_986) );
INVx1_ASAP7_75t_L g1881 ( .A(n_239), .Y(n_1881) );
AOI22xp33_ASAP7_75t_L g1808 ( .A1(n_240), .A2(n_250), .B1(n_539), .B2(n_622), .Y(n_1808) );
INVxp33_ASAP7_75t_L g1832 ( .A(n_240), .Y(n_1832) );
INVx1_ASAP7_75t_L g661 ( .A(n_241), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_241), .A2(n_258), .B1(n_702), .B2(n_704), .C(n_705), .Y(n_701) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_242), .Y(n_613) );
XNOR2x1_ASAP7_75t_L g850 ( .A(n_243), .B(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g456 ( .A(n_244), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g1623 ( .A(n_245), .Y(n_1623) );
BUFx3_ASAP7_75t_L g490 ( .A(n_246), .Y(n_490) );
INVx1_ASAP7_75t_L g498 ( .A(n_246), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g1187 ( .A(n_247), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g1457 ( .A(n_248), .Y(n_1457) );
AO221x2_ASAP7_75t_L g1553 ( .A1(n_249), .A2(n_317), .B1(n_1554), .B2(n_1561), .C(n_1564), .Y(n_1553) );
INVxp33_ASAP7_75t_L g1828 ( .A(n_250), .Y(n_1828) );
AOI22xp5_ASAP7_75t_L g1601 ( .A1(n_251), .A2(n_252), .B1(n_1556), .B2(n_1602), .Y(n_1601) );
AOI22xp5_ASAP7_75t_L g1851 ( .A1(n_251), .A2(n_1852), .B1(n_1856), .B2(n_1914), .Y(n_1851) );
AO22x2_ASAP7_75t_L g1857 ( .A1(n_251), .A2(n_1858), .B1(n_1912), .B2(n_1913), .Y(n_1857) );
INVxp67_ASAP7_75t_L g1912 ( .A(n_251), .Y(n_1912) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_253), .Y(n_358) );
AND2x2_ASAP7_75t_L g387 ( .A(n_253), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_253), .B(n_321), .Y(n_419) );
INVx1_ASAP7_75t_L g470 ( .A(n_253), .Y(n_470) );
INVxp67_ASAP7_75t_L g591 ( .A(n_254), .Y(n_591) );
INVx1_ASAP7_75t_L g1162 ( .A(n_255), .Y(n_1162) );
AOI21xp5_ASAP7_75t_L g1516 ( .A1(n_256), .A2(n_1517), .B(n_1518), .Y(n_1516) );
INVx1_ASAP7_75t_L g1535 ( .A(n_256), .Y(n_1535) );
OAI332xp33_ASAP7_75t_L g1182 ( .A1(n_257), .A2(n_428), .A3(n_466), .B1(n_1183), .B2(n_1186), .B3(n_1190), .C1(n_1193), .C2(n_1196), .Y(n_1182) );
INVx1_ASAP7_75t_L g1227 ( .A(n_257), .Y(n_1227) );
INVx1_ASAP7_75t_L g656 ( .A(n_258), .Y(n_656) );
INVx2_ASAP7_75t_L g485 ( .A(n_259), .Y(n_485) );
OR2x2_ASAP7_75t_L g500 ( .A(n_259), .B(n_483), .Y(n_500) );
INVx1_ASAP7_75t_L g784 ( .A(n_260), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g1185 ( .A(n_262), .Y(n_1185) );
INVx1_ASAP7_75t_L g995 ( .A(n_263), .Y(n_995) );
INVxp67_ASAP7_75t_L g440 ( .A(n_264), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_264), .A2(n_314), .B1(n_538), .B2(n_540), .C(n_545), .Y(n_537) );
INVx1_ASAP7_75t_L g908 ( .A(n_265), .Y(n_908) );
CKINVDCx16_ASAP7_75t_R g1080 ( .A(n_266), .Y(n_1080) );
INVx1_ASAP7_75t_L g817 ( .A(n_267), .Y(n_817) );
INVx1_ASAP7_75t_L g751 ( .A(n_268), .Y(n_751) );
INVxp67_ASAP7_75t_SL g1420 ( .A(n_269), .Y(n_1420) );
OAI211xp5_ASAP7_75t_SL g1431 ( .A1(n_269), .A2(n_448), .B(n_984), .C(n_1432), .Y(n_1431) );
INVx1_ASAP7_75t_L g1308 ( .A(n_270), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_270), .A2(n_302), .B1(n_1319), .B2(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1811 ( .A(n_271), .Y(n_1811) );
INVxp67_ASAP7_75t_L g1360 ( .A(n_272), .Y(n_1360) );
INVx1_ASAP7_75t_L g1334 ( .A(n_273), .Y(n_1334) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_274), .A2(n_298), .B1(n_621), .B2(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g900 ( .A(n_274), .Y(n_900) );
AOI22xp5_ASAP7_75t_SL g1607 ( .A1(n_275), .A2(n_278), .B1(n_1556), .B2(n_1562), .Y(n_1607) );
INVx1_ASAP7_75t_L g461 ( .A(n_276), .Y(n_461) );
INVxp67_ASAP7_75t_SL g1521 ( .A(n_277), .Y(n_1521) );
XNOR2xp5_ASAP7_75t_L g1235 ( .A(n_278), .B(n_1236), .Y(n_1235) );
AOI221xp5_ASAP7_75t_L g1512 ( .A1(n_279), .A2(n_288), .B1(n_629), .B2(n_1513), .C(n_1514), .Y(n_1512) );
INVxp33_ASAP7_75t_L g1534 ( .A(n_279), .Y(n_1534) );
INVx1_ASAP7_75t_L g665 ( .A(n_280), .Y(n_665) );
INVx1_ASAP7_75t_L g1340 ( .A(n_281), .Y(n_1340) );
INVx1_ASAP7_75t_L g931 ( .A(n_283), .Y(n_931) );
AOI21xp5_ASAP7_75t_L g957 ( .A1(n_283), .A2(n_529), .B(n_708), .Y(n_957) );
INVx1_ASAP7_75t_L g884 ( .A(n_284), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g646 ( .A(n_285), .Y(n_646) );
INVxp33_ASAP7_75t_L g1436 ( .A(n_286), .Y(n_1436) );
AOI22xp33_ASAP7_75t_L g1372 ( .A1(n_287), .A2(n_306), .B1(n_1373), .B2(n_1374), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g1385 ( .A1(n_287), .A2(n_306), .B1(n_1386), .B2(n_1387), .Y(n_1385) );
CKINVDCx5p33_ASAP7_75t_R g1456 ( .A(n_289), .Y(n_1456) );
INVx1_ASAP7_75t_L g1842 ( .A(n_290), .Y(n_1842) );
INVx1_ASAP7_75t_L g1317 ( .A(n_291), .Y(n_1317) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_292), .Y(n_668) );
INVx1_ASAP7_75t_L g935 ( .A(n_293), .Y(n_935) );
AOI221xp5_ASAP7_75t_L g894 ( .A1(n_294), .A2(n_298), .B1(n_895), .B2(n_897), .C(n_899), .Y(n_894) );
INVxp67_ASAP7_75t_L g1343 ( .A(n_295), .Y(n_1343) );
INVx1_ASAP7_75t_L g1887 ( .A(n_297), .Y(n_1887) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_299), .A2(n_332), .B1(n_634), .B2(n_841), .Y(n_1041) );
INVx1_ASAP7_75t_L g1067 ( .A(n_299), .Y(n_1067) );
INVx1_ASAP7_75t_L g893 ( .A(n_301), .Y(n_893) );
INVx1_ASAP7_75t_L g1306 ( .A(n_302), .Y(n_1306) );
CKINVDCx5p33_ASAP7_75t_R g867 ( .A(n_303), .Y(n_867) );
INVx1_ASAP7_75t_L g1003 ( .A(n_305), .Y(n_1003) );
INVx1_ASAP7_75t_L g1494 ( .A(n_307), .Y(n_1494) );
INVx1_ASAP7_75t_L g749 ( .A(n_308), .Y(n_749) );
INVx1_ASAP7_75t_L g1806 ( .A(n_310), .Y(n_1806) );
INVx1_ASAP7_75t_L g792 ( .A(n_311), .Y(n_792) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_312), .Y(n_352) );
AND3x2_ASAP7_75t_L g1559 ( .A(n_312), .B(n_350), .C(n_1560), .Y(n_1559) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_312), .B(n_350), .Y(n_1569) );
INVx2_ASAP7_75t_L g363 ( .A(n_313), .Y(n_363) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_314), .Y(n_447) );
INVxp33_ASAP7_75t_SL g436 ( .A(n_315), .Y(n_436) );
INVx1_ASAP7_75t_L g725 ( .A(n_316), .Y(n_725) );
CKINVDCx5p33_ASAP7_75t_R g1184 ( .A(n_318), .Y(n_1184) );
INVx1_ASAP7_75t_L g820 ( .A(n_319), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g1473 ( .A(n_320), .Y(n_1473) );
INVx1_ASAP7_75t_L g365 ( .A(n_321), .Y(n_365) );
INVx2_ASAP7_75t_L g388 ( .A(n_321), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g1472 ( .A(n_322), .Y(n_1472) );
INVxp67_ASAP7_75t_SL g814 ( .A(n_323), .Y(n_814) );
INVx1_ASAP7_75t_L g881 ( .A(n_324), .Y(n_881) );
INVxp33_ASAP7_75t_L g579 ( .A(n_325), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_325), .A2(n_326), .B1(n_550), .B2(n_617), .C(n_618), .Y(n_616) );
INVxp33_ASAP7_75t_L g577 ( .A(n_326), .Y(n_577) );
INVxp67_ASAP7_75t_SL g1507 ( .A(n_327), .Y(n_1507) );
INVx1_ASAP7_75t_L g818 ( .A(n_328), .Y(n_818) );
INVxp67_ASAP7_75t_SL g1547 ( .A(n_329), .Y(n_1547) );
INVx1_ASAP7_75t_L g1060 ( .A(n_332), .Y(n_1060) );
INVx1_ASAP7_75t_L g1422 ( .A(n_333), .Y(n_1422) );
INVx1_ASAP7_75t_L g1480 ( .A(n_334), .Y(n_1480) );
CKINVDCx5p33_ASAP7_75t_R g1504 ( .A(n_335), .Y(n_1504) );
CKINVDCx5p33_ASAP7_75t_R g1028 ( .A(n_336), .Y(n_1028) );
INVx1_ASAP7_75t_L g1266 ( .A(n_337), .Y(n_1266) );
AOI21xp5_ASAP7_75t_L g1284 ( .A1(n_337), .A2(n_917), .B(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g1823 ( .A(n_338), .Y(n_1823) );
INVx1_ASAP7_75t_L g821 ( .A(n_339), .Y(n_821) );
INVxp33_ASAP7_75t_SL g397 ( .A(n_340), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_341), .Y(n_733) );
INVx1_ASAP7_75t_L g756 ( .A(n_342), .Y(n_756) );
INVxp33_ASAP7_75t_L g576 ( .A(n_343), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_366), .B(n_1550), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_353), .Y(n_347) );
AND2x4_ASAP7_75t_L g1855 ( .A(n_348), .B(n_354), .Y(n_1855) );
NOR2xp33_ASAP7_75t_SL g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_SL g1850 ( .A(n_349), .Y(n_1850) );
NAND2xp5_ASAP7_75t_L g1919 ( .A(n_349), .B(n_351), .Y(n_1919) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g1849 ( .A(n_351), .B(n_1850), .Y(n_1849) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_359), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g1366 ( .A(n_356), .B(n_479), .Y(n_1366) );
OR2x6_ASAP7_75t_L g1890 ( .A(n_356), .B(n_479), .Y(n_1890) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g765 ( .A(n_357), .B(n_365), .Y(n_765) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g429 ( .A(n_358), .B(n_430), .Y(n_429) );
INVx8_ASAP7_75t_L g1362 ( .A(n_359), .Y(n_1362) );
OR2x6_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
INVx1_ASAP7_75t_L g435 ( .A(n_360), .Y(n_435) );
OR2x2_ASAP7_75t_L g476 ( .A(n_360), .B(n_418), .Y(n_476) );
INVx2_ASAP7_75t_SL g595 ( .A(n_360), .Y(n_595) );
INVx2_ASAP7_75t_SL g606 ( .A(n_360), .Y(n_606) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_360), .Y(n_667) );
BUFx2_ASAP7_75t_L g901 ( .A(n_360), .Y(n_901) );
OAI22xp33_ASAP7_75t_L g907 ( .A1(n_360), .A2(n_450), .B1(n_867), .B2(n_908), .Y(n_907) );
OAI22xp5_ASAP7_75t_L g1168 ( .A1(n_360), .A2(n_450), .B1(n_1144), .B2(n_1169), .Y(n_1168) );
OR2x6_ASAP7_75t_L g1365 ( .A(n_360), .B(n_1355), .Y(n_1365) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx2_ASAP7_75t_L g382 ( .A(n_362), .Y(n_382) );
INVx1_ASAP7_75t_L g394 ( .A(n_362), .Y(n_394) );
AND2x2_ASAP7_75t_L g402 ( .A(n_362), .B(n_363), .Y(n_402) );
AND2x4_ASAP7_75t_L g409 ( .A(n_362), .B(n_395), .Y(n_409) );
INVx1_ASAP7_75t_L g453 ( .A(n_362), .Y(n_453) );
INVx1_ASAP7_75t_L g384 ( .A(n_363), .Y(n_384) );
INVx2_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
INVx1_ASAP7_75t_L g416 ( .A(n_363), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_363), .B(n_382), .Y(n_446) );
INVx1_ASAP7_75t_L g452 ( .A(n_363), .Y(n_452) );
AND2x4_ASAP7_75t_L g1351 ( .A(n_364), .B(n_416), .Y(n_1351) );
INVx2_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g1352 ( .A(n_365), .B(n_759), .Y(n_1352) );
OAI22xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_1072), .B2(n_1073), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_716), .B2(n_1071), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
XNOR2x1_ASAP7_75t_L g371 ( .A(n_372), .B(n_570), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
XNOR2x1_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_471), .Y(n_375) );
NOR3xp33_ASAP7_75t_SL g376 ( .A(n_377), .B(n_410), .C(n_426), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_379), .A2(n_399), .B1(n_579), .B2(n_580), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_379), .A2(n_399), .B1(n_1053), .B2(n_1054), .Y(n_1052) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_385), .Y(n_379) );
AND2x2_ASAP7_75t_L g648 ( .A(n_380), .B(n_385), .Y(n_648) );
AND2x2_ASAP7_75t_L g789 ( .A(n_380), .B(n_385), .Y(n_789) );
AND2x2_ASAP7_75t_L g934 ( .A(n_380), .B(n_385), .Y(n_934) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_380), .B(n_385), .Y(n_1437) );
INVx2_ASAP7_75t_SL g1441 ( .A(n_380), .Y(n_1441) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_L g773 ( .A(n_381), .Y(n_773) );
INVx1_ASAP7_75t_L g896 ( .A(n_381), .Y(n_896) );
INVx1_ASAP7_75t_L g905 ( .A(n_381), .Y(n_905) );
BUFx6f_ASAP7_75t_L g922 ( .A(n_381), .Y(n_922) );
BUFx6f_ASAP7_75t_L g926 ( .A(n_381), .Y(n_926) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_381), .B(n_387), .Y(n_1307) );
AND2x4_ASAP7_75t_L g1354 ( .A(n_381), .B(n_1355), .Y(n_1354) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g424 ( .A(n_382), .Y(n_424) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x6_ASAP7_75t_L g391 ( .A(n_385), .B(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g399 ( .A(n_385), .B(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g406 ( .A(n_385), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g891 ( .A(n_385), .B(n_892), .Y(n_891) );
AND2x2_ASAP7_75t_L g938 ( .A(n_385), .B(n_602), .Y(n_938) );
AND2x2_ASAP7_75t_L g975 ( .A(n_385), .B(n_781), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_385), .A2(n_782), .B1(n_1108), .B2(n_1114), .Y(n_1107) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g467 ( .A(n_386), .Y(n_467) );
INVx2_ASAP7_75t_L g1301 ( .A(n_387), .Y(n_1301) );
AND2x4_ASAP7_75t_L g1304 ( .A(n_387), .B(n_768), .Y(n_1304) );
INVx1_ASAP7_75t_L g430 ( .A(n_388), .Y(n_430) );
INVx1_ASAP7_75t_L g469 ( .A(n_388), .Y(n_469) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g1533 ( .A1(n_390), .A2(n_643), .B1(n_1534), .B2(n_1535), .Y(n_1533) );
BUFx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_391), .A2(n_406), .B1(n_576), .B2(n_577), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_391), .A2(n_642), .B1(n_643), .B2(n_644), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_391), .A2(n_733), .B1(n_784), .B2(n_785), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_391), .A2(n_785), .B1(n_797), .B2(n_798), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_391), .A2(n_789), .B1(n_884), .B2(n_885), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_391), .A2(n_934), .B1(n_935), .B2(n_936), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_391), .A2(n_1049), .B1(n_1050), .B2(n_1051), .Y(n_1048) );
INVx1_ASAP7_75t_SL g1177 ( .A(n_391), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1491 ( .A1(n_391), .A2(n_406), .B1(n_1461), .B2(n_1492), .Y(n_1491) );
AOI22xp33_ASAP7_75t_L g1827 ( .A1(n_391), .A2(n_1806), .B1(n_1828), .B2(n_1829), .Y(n_1827) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_392), .B(n_417), .Y(n_425) );
BUFx2_ASAP7_75t_L g1430 ( .A(n_392), .Y(n_1430) );
BUFx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx2_ASAP7_75t_L g762 ( .A(n_393), .Y(n_762) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_393), .Y(n_771) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_393), .Y(n_781) );
INVx1_ASAP7_75t_L g920 ( .A(n_393), .Y(n_920) );
BUFx3_ASAP7_75t_L g1302 ( .A(n_393), .Y(n_1302) );
AND2x4_ASAP7_75t_L g1346 ( .A(n_393), .B(n_1347), .Y(n_1346) );
AND2x4_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B1(n_403), .B2(n_404), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g1474 ( .A1(n_398), .A2(n_1462), .B(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1532 ( .A(n_398), .Y(n_1532) );
BUFx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_399), .A2(n_646), .B1(n_647), .B2(n_648), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_399), .A2(n_787), .B1(n_788), .B2(n_789), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_399), .A2(n_789), .B1(n_800), .B2(n_801), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_399), .B(n_931), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g1434 ( .A1(n_399), .A2(n_1435), .B1(n_1436), .B2(n_1437), .Y(n_1434) );
AOI22xp33_ASAP7_75t_L g1830 ( .A1(n_399), .A2(n_1437), .B1(n_1831), .B2(n_1832), .Y(n_1830) );
INVx2_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g779 ( .A(n_401), .Y(n_779) );
INVx2_ASAP7_75t_SL g892 ( .A(n_401), .Y(n_892) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx6f_ASAP7_75t_L g768 ( .A(n_402), .Y(n_768) );
OAI221xp5_ASAP7_75t_L g512 ( .A1(n_403), .A2(n_513), .B1(n_514), .B2(n_515), .C(n_519), .Y(n_512) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_L g643 ( .A(n_406), .Y(n_643) );
BUFx2_ASAP7_75t_L g785 ( .A(n_406), .Y(n_785) );
BUFx2_ASAP7_75t_L g1050 ( .A(n_406), .Y(n_1050) );
BUFx2_ASAP7_75t_L g1829 ( .A(n_406), .Y(n_1829) );
BUFx3_ASAP7_75t_L g673 ( .A(n_407), .Y(n_673) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g602 ( .A(n_408), .Y(n_602) );
BUFx6f_ASAP7_75t_L g924 ( .A(n_408), .Y(n_924) );
INVx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_409), .Y(n_438) );
INVx1_ASAP7_75t_L g1001 ( .A(n_409), .Y(n_1001) );
INVx1_ASAP7_75t_L g1359 ( .A(n_409), .Y(n_1359) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g582 ( .A(n_412), .Y(n_582) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_413), .Y(n_1056) );
NAND2x1_ASAP7_75t_SL g413 ( .A(n_414), .B(n_417), .Y(n_413) );
NAND2x1p5_ASAP7_75t_L g1287 ( .A(n_414), .B(n_1288), .Y(n_1287) );
AOI22xp33_ASAP7_75t_L g1432 ( .A1(n_414), .A2(n_423), .B1(n_1421), .B2(n_1422), .Y(n_1432) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_416), .Y(n_755) );
NAND2x1p5_ASAP7_75t_L g422 ( .A(n_417), .B(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g754 ( .A(n_417), .B(n_755), .Y(n_754) );
AND2x4_ASAP7_75t_L g757 ( .A(n_417), .B(n_758), .Y(n_757) );
AND2x4_ASAP7_75t_L g761 ( .A(n_417), .B(n_762), .Y(n_761) );
AOI32xp33_ASAP7_75t_L g1426 ( .A1(n_417), .A2(n_1382), .A3(n_1427), .B1(n_1429), .B2(n_1431), .Y(n_1426) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g1279 ( .A(n_419), .Y(n_1279) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx4f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx4f_ASAP7_75t_L g583 ( .A(n_422), .Y(n_583) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x6_ASAP7_75t_L g1289 ( .A(n_424), .B(n_1278), .Y(n_1289) );
BUFx2_ASAP7_75t_L g584 ( .A(n_425), .Y(n_584) );
BUFx2_ASAP7_75t_L g650 ( .A(n_425), .Y(n_650) );
BUFx3_ASAP7_75t_L g980 ( .A(n_425), .Y(n_980) );
OAI33xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_432), .A3(n_439), .B1(n_454), .B2(n_457), .B3(n_462), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI33xp33_ASAP7_75t_L g585 ( .A1(n_428), .A2(n_464), .A3(n_586), .B1(n_593), .B2(n_599), .B3(n_604), .Y(n_585) );
OAI33xp33_ASAP7_75t_L g651 ( .A1(n_428), .A2(n_464), .A3(n_652), .B1(n_657), .B2(n_666), .B3(n_671), .Y(n_651) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_428), .Y(n_804) );
OAI33xp33_ASAP7_75t_L g981 ( .A1(n_428), .A2(n_982), .A3(n_988), .B1(n_994), .B2(n_1002), .B3(n_1005), .Y(n_981) );
OAI33xp33_ASAP7_75t_L g1057 ( .A1(n_428), .A2(n_464), .A3(n_1058), .B1(n_1064), .B2(n_1069), .B3(n_1070), .Y(n_1057) );
OAI33xp33_ASAP7_75t_L g1475 ( .A1(n_428), .A2(n_1476), .A3(n_1479), .B1(n_1481), .B2(n_1486), .B3(n_1489), .Y(n_1475) );
OAI33xp33_ASAP7_75t_L g1834 ( .A1(n_428), .A2(n_464), .A3(n_1835), .B1(n_1838), .B2(n_1843), .B3(n_1845), .Y(n_1834) );
OR2x6_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g1355 ( .A(n_430), .Y(n_1355) );
BUFx2_ASAP7_75t_L g569 ( .A(n_431), .Y(n_569) );
INVx2_ASAP7_75t_L g713 ( .A(n_431), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_436), .B2(n_437), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g457 ( .A1(n_434), .A2(n_458), .B1(n_459), .B2(n_461), .Y(n_457) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g1188 ( .A(n_435), .Y(n_1188) );
INVx1_ASAP7_75t_L g1443 ( .A(n_435), .Y(n_1443) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_437), .A2(n_441), .B1(n_455), .B2(n_456), .Y(n_454) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx4_ASAP7_75t_L g592 ( .A(n_438), .Y(n_592) );
INVx2_ASAP7_75t_SL g1122 ( .A(n_438), .Y(n_1122) );
BUFx3_ASAP7_75t_L g1841 ( .A(n_438), .Y(n_1841) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_447), .B2(n_448), .Y(n_439) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g1183 ( .A1(n_443), .A2(n_592), .B1(n_1184), .B2(n_1185), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1843 ( .A1(n_443), .A2(n_1803), .B1(n_1824), .B2(n_1844), .Y(n_1843) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g996 ( .A(n_444), .Y(n_996) );
INVx2_ASAP7_75t_L g1109 ( .A(n_444), .Y(n_1109) );
INVx2_ASAP7_75t_SL g1482 ( .A(n_444), .Y(n_1482) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g590 ( .A(n_445), .Y(n_590) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g660 ( .A(n_446), .Y(n_660) );
INVx1_ASAP7_75t_L g813 ( .A(n_446), .Y(n_813) );
OAI22xp33_ASAP7_75t_L g819 ( .A1(n_448), .A2(n_806), .B1(n_820), .B2(n_821), .Y(n_819) );
OAI22xp5_ASAP7_75t_SL g1002 ( .A1(n_448), .A2(n_594), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1070 ( .A1(n_448), .A2(n_1027), .B1(n_1043), .B2(n_1059), .Y(n_1070) );
OAI22xp5_ASAP7_75t_SL g1193 ( .A1(n_448), .A2(n_667), .B1(n_1194), .B2(n_1195), .Y(n_1193) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g597 ( .A(n_449), .Y(n_597) );
INVx2_ASAP7_75t_L g1445 ( .A(n_449), .Y(n_1445) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx3_ASAP7_75t_L g460 ( .A(n_450), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_450), .A2(n_900), .B1(n_901), .B2(n_902), .Y(n_899) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
AND2x2_ASAP7_75t_L g610 ( .A(n_452), .B(n_453), .Y(n_610) );
INVx1_ASAP7_75t_L g759 ( .A(n_453), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_455), .A2(n_494), .B(n_501), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_456), .A2(n_458), .B1(n_559), .B2(n_564), .Y(n_558) );
BUFx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g1186 ( .A1(n_460), .A2(n_1187), .B1(n_1188), .B2(n_1189), .Y(n_1186) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_461), .A2(n_533), .B1(n_537), .B2(n_548), .C(n_553), .Y(n_532) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI33xp33_ASAP7_75t_L g1537 ( .A1(n_463), .A2(n_1538), .A3(n_1540), .B1(n_1541), .B2(n_1544), .B3(n_1545), .Y(n_1537) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OAI33xp33_ASAP7_75t_L g803 ( .A1(n_464), .A2(n_804), .A3(n_805), .B1(n_810), .B2(n_816), .B3(n_819), .Y(n_803) );
CKINVDCx8_ASAP7_75t_R g464 ( .A(n_465), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g1896 ( .A(n_465), .B(n_1897), .C(n_1899), .Y(n_1896) );
INVx5_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx6_ASAP7_75t_L g782 ( .A(n_466), .Y(n_782) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx2_ASAP7_75t_L g929 ( .A(n_468), .Y(n_929) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g1348 ( .A(n_469), .Y(n_1348) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_491), .B(n_492), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI21xp33_ASAP7_75t_SL g612 ( .A1(n_474), .A2(n_613), .B(n_614), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_474), .A2(n_722), .B1(n_723), .B2(n_751), .Y(n_721) );
AOI21xp33_ASAP7_75t_SL g1799 ( .A1(n_474), .A2(n_1800), .B(n_1801), .Y(n_1799) );
INVx5_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g677 ( .A(n_475), .Y(n_677) );
INVx1_ASAP7_75t_L g847 ( .A(n_475), .Y(n_847) );
INVx2_ASAP7_75t_SL g1019 ( .A(n_475), .Y(n_1019) );
INVx2_ASAP7_75t_L g1045 ( .A(n_475), .Y(n_1045) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx2_ASAP7_75t_L g889 ( .A(n_476), .Y(n_889) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
AND2x4_ASAP7_75t_L g1321 ( .A(n_479), .B(n_530), .Y(n_1321) );
AND2x4_ASAP7_75t_L g1911 ( .A(n_479), .B(n_530), .Y(n_1911) );
INVx2_ASAP7_75t_L g876 ( .A(n_480), .Y(n_876) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_486), .Y(n_480) );
AND2x4_ASAP7_75t_L g503 ( .A(n_481), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g508 ( .A(n_481), .Y(n_508) );
AND2x4_ASAP7_75t_L g626 ( .A(n_481), .B(n_510), .Y(n_626) );
AND2x2_ASAP7_75t_L g684 ( .A(n_481), .B(n_510), .Y(n_684) );
AND2x4_ASAP7_75t_L g844 ( .A(n_481), .B(n_504), .Y(n_844) );
BUFx2_ASAP7_75t_L g865 ( .A(n_481), .Y(n_865) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_481), .B(n_510), .Y(n_1092) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x4_ASAP7_75t_L g530 ( .A(n_484), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g547 ( .A(n_485), .B(n_531), .Y(n_547) );
INVx1_ASAP7_75t_L g1243 ( .A(n_485), .Y(n_1243) );
HB1xp67_ASAP7_75t_L g1248 ( .A(n_485), .Y(n_1248) );
INVx1_ASAP7_75t_L g1252 ( .A(n_485), .Y(n_1252) );
INVx6_ASAP7_75t_L g526 ( .A(n_486), .Y(n_526) );
BUFx2_ASAP7_75t_L g838 ( .A(n_486), .Y(n_838) );
INVx2_ASAP7_75t_L g1033 ( .A(n_486), .Y(n_1033) );
AND2x4_ASAP7_75t_L g1246 ( .A(n_486), .B(n_1247), .Y(n_1246) );
AND2x4_ASAP7_75t_L g486 ( .A(n_487), .B(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g511 ( .A(n_487), .Y(n_511) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g497 ( .A(n_488), .B(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g522 ( .A(n_488), .B(n_490), .Y(n_522) );
INVx1_ASAP7_75t_L g506 ( .A(n_489), .Y(n_506) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x4_ASAP7_75t_L g517 ( .A(n_490), .B(n_518), .Y(n_517) );
AOI31xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_532), .A3(n_558), .B(n_567), .Y(n_492) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_495), .A2(n_600), .B1(n_616), .B2(n_619), .C(n_623), .Y(n_615) );
AOI211xp5_ASAP7_75t_L g680 ( .A1(n_495), .A2(n_670), .B(n_681), .C(n_685), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_495), .A2(n_559), .B1(n_749), .B2(n_750), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g1414 ( .A1(n_495), .A2(n_559), .B1(n_1415), .B2(n_1416), .Y(n_1414) );
INVx1_ASAP7_75t_L g1509 ( .A(n_495), .Y(n_1509) );
AOI21xp5_ASAP7_75t_L g1802 ( .A1(n_495), .A2(n_1803), .B(n_1804), .Y(n_1802) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_499), .Y(n_495) );
INVx2_ASAP7_75t_SL g513 ( .A(n_496), .Y(n_513) );
INVx1_ASAP7_75t_L g687 ( .A(n_496), .Y(n_687) );
BUFx3_ASAP7_75t_L g1097 ( .A(n_496), .Y(n_1097) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_497), .Y(n_539) );
BUFx2_ASAP7_75t_L g629 ( .A(n_497), .Y(n_629) );
INVx2_ASAP7_75t_SL g703 ( .A(n_497), .Y(n_703) );
BUFx6f_ASAP7_75t_L g743 ( .A(n_497), .Y(n_743) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_497), .Y(n_829) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_497), .Y(n_860) );
BUFx2_ASAP7_75t_L g872 ( .A(n_497), .Y(n_872) );
BUFx3_ASAP7_75t_L g952 ( .A(n_497), .Y(n_952) );
AND2x6_ASAP7_75t_L g1270 ( .A(n_497), .B(n_1242), .Y(n_1270) );
INVx1_ASAP7_75t_L g563 ( .A(n_498), .Y(n_563) );
AND2x4_ASAP7_75t_L g536 ( .A(n_499), .B(n_521), .Y(n_536) );
AND2x2_ASAP7_75t_L g828 ( .A(n_499), .B(n_829), .Y(n_828) );
AOI221xp5_ASAP7_75t_L g866 ( .A1(n_499), .A2(n_559), .B1(n_867), .B2(n_868), .C(n_875), .Y(n_866) );
A2O1A1Ixp33_ASAP7_75t_L g960 ( .A1(n_499), .A2(n_617), .B(n_961), .C(n_962), .Y(n_960) );
AOI222xp33_ASAP7_75t_L g1083 ( .A1(n_499), .A2(n_503), .B1(n_1084), .B2(n_1091), .C1(n_1092), .C2(n_1093), .Y(n_1083) );
OAI21xp5_ASAP7_75t_L g1130 ( .A1(n_499), .A2(n_1131), .B(n_1134), .Y(n_1130) );
OAI21xp33_ASAP7_75t_L g1466 ( .A1(n_499), .A2(n_1467), .B(n_1469), .Y(n_1466) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g560 ( .A(n_500), .B(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g565 ( .A(n_500), .B(n_566), .Y(n_565) );
A2O1A1Ixp33_ASAP7_75t_SL g1198 ( .A1(n_500), .A2(n_1199), .B(n_1203), .C(n_1208), .Y(n_1198) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_SL g624 ( .A(n_503), .Y(n_624) );
INVx1_ASAP7_75t_L g682 ( .A(n_503), .Y(n_682) );
AOI222xp33_ASAP7_75t_L g1419 ( .A1(n_503), .A2(n_684), .B1(n_1102), .B2(n_1420), .C1(n_1421), .C2(n_1422), .Y(n_1419) );
INVxp67_ASAP7_75t_L g1140 ( .A(n_504), .Y(n_1140) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g1262 ( .A(n_506), .Y(n_1262) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
INVx1_ASAP7_75t_SL g556 ( .A(n_508), .Y(n_556) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g1141 ( .A(n_510), .Y(n_1141) );
BUFx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x6_ASAP7_75t_L g1264 ( .A(n_511), .B(n_1243), .Y(n_1264) );
INVx1_ASAP7_75t_L g620 ( .A(n_513), .Y(n_620) );
INVx1_ASAP7_75t_L g747 ( .A(n_515), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g1220 ( .A1(n_515), .A2(n_1221), .B1(n_1222), .B2(n_1223), .Y(n_1220) );
INVx1_ASAP7_75t_L g1513 ( .A(n_515), .Y(n_1513) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g552 ( .A(n_516), .Y(n_552) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_516), .Y(n_874) );
BUFx6f_ASAP7_75t_L g1017 ( .A(n_516), .Y(n_1017) );
AND2x6_ASAP7_75t_L g1250 ( .A(n_516), .B(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1378 ( .A(n_516), .Y(n_1378) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g566 ( .A(n_517), .Y(n_566) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_517), .Y(n_622) );
INVx1_ASAP7_75t_L g689 ( .A(n_517), .Y(n_689) );
INVx1_ASAP7_75t_L g1202 ( .A(n_517), .Y(n_1202) );
INVx1_ASAP7_75t_L g562 ( .A(n_518), .Y(n_562) );
BUFx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx4f_ASAP7_75t_L g617 ( .A(n_521), .Y(n_617) );
INVx2_ASAP7_75t_SL g856 ( .A(n_521), .Y(n_856) );
AND2x4_ASAP7_75t_L g864 ( .A(n_521), .B(n_865), .Y(n_864) );
BUFx6f_ASAP7_75t_L g1207 ( .A(n_521), .Y(n_1207) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_522), .Y(n_544) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_525), .Y(n_550) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_526), .Y(n_635) );
INVx1_ASAP7_75t_L g708 ( .A(n_526), .Y(n_708) );
INVx2_ASAP7_75t_L g735 ( .A(n_526), .Y(n_735) );
INVx2_ASAP7_75t_SL g835 ( .A(n_526), .Y(n_835) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_526), .Y(n_863) );
INVx1_ASAP7_75t_L g1101 ( .A(n_526), .Y(n_1101) );
INVx2_ASAP7_75t_L g1268 ( .A(n_526), .Y(n_1268) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OAI221xp5_ASAP7_75t_L g1460 ( .A1(n_528), .A2(n_694), .B1(n_1135), .B2(n_1461), .C(n_1462), .Y(n_1460) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_530), .Y(n_618) );
INVx2_ASAP7_75t_L g697 ( .A(n_530), .Y(n_697) );
INVx1_ASAP7_75t_L g839 ( .A(n_530), .Y(n_839) );
INVx1_ASAP7_75t_L g1272 ( .A(n_531), .Y(n_1272) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_535), .A2(n_555), .B1(n_611), .B2(n_628), .C(n_633), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g1810 ( .A1(n_535), .A2(n_555), .B1(n_1811), .B2(n_1812), .C(n_1820), .Y(n_1810) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g700 ( .A(n_536), .Y(n_700) );
INVx2_ASAP7_75t_SL g738 ( .A(n_536), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g1013 ( .A1(n_536), .A2(n_864), .B1(n_1004), .B2(n_1014), .C(n_1016), .Y(n_1013) );
INVx1_ASAP7_75t_L g1418 ( .A(n_536), .Y(n_1418) );
BUFx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g729 ( .A(n_539), .Y(n_729) );
BUFx3_ASAP7_75t_L g858 ( .A(n_539), .Y(n_858) );
INVx1_ASAP7_75t_L g963 ( .A(n_539), .Y(n_963) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g704 ( .A(n_541), .Y(n_704) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g1257 ( .A(n_543), .Y(n_1257) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_544), .Y(n_557) );
BUFx6f_ASAP7_75t_L g1015 ( .A(n_544), .Y(n_1015) );
AND2x4_ASAP7_75t_L g1240 ( .A(n_544), .B(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1817 ( .A(n_544), .Y(n_1817) );
BUFx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g1819 ( .A(n_546), .Y(n_1819) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
BUFx3_ASAP7_75t_L g632 ( .A(n_547), .Y(n_632) );
INVx1_ASAP7_75t_L g705 ( .A(n_547), .Y(n_705) );
INVx2_ASAP7_75t_L g1149 ( .A(n_547), .Y(n_1149) );
INVx1_ASAP7_75t_L g1906 ( .A(n_547), .Y(n_1906) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_555), .A2(n_675), .B1(n_699), .B2(n_701), .C(n_706), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_555), .A2(n_737), .B1(n_739), .B2(n_740), .C(n_746), .Y(n_736) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_555), .A2(n_737), .B1(n_821), .B2(n_831), .C(n_832), .Y(n_830) );
AOI21xp33_ASAP7_75t_L g1094 ( .A1(n_555), .A2(n_1095), .B(n_1096), .Y(n_1094) );
INVx1_ASAP7_75t_L g1208 ( .A(n_555), .Y(n_1208) );
INVx1_ASAP7_75t_L g1423 ( .A(n_555), .Y(n_1423) );
HB1xp67_ASAP7_75t_L g1525 ( .A(n_555), .Y(n_1525) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_557), .Y(n_630) );
INVx1_ASAP7_75t_L g745 ( .A(n_557), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g1088 ( .A1(n_557), .A2(n_829), .B1(n_1089), .B2(n_1090), .Y(n_1088) );
OAI21xp33_ASAP7_75t_L g1872 ( .A1(n_557), .A2(n_1241), .B(n_1873), .Y(n_1872) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_559), .A2(n_564), .B1(n_603), .B2(n_607), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_559), .A2(n_564), .B1(n_668), .B2(n_674), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_559), .A2(n_817), .B1(n_820), .B2(n_826), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g1018 ( .A1(n_559), .A2(n_564), .B1(n_997), .B2(n_1003), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_559), .A2(n_828), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1526 ( .A1(n_559), .A2(n_564), .B1(n_1527), .B2(n_1528), .Y(n_1526) );
AOI22xp33_ASAP7_75t_L g1822 ( .A1(n_559), .A2(n_564), .B1(n_1823), .B2(n_1824), .Y(n_1822) );
INVx6_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g695 ( .A(n_561), .Y(n_695) );
INVx2_ASAP7_75t_L g1086 ( .A(n_561), .Y(n_1086) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g693 ( .A(n_562), .B(n_563), .Y(n_693) );
AOI211xp5_ASAP7_75t_L g724 ( .A1(n_564), .A2(n_725), .B(n_726), .C(n_727), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g836 ( .A1(n_564), .A2(n_818), .B1(n_837), .B2(n_840), .C(n_842), .Y(n_836) );
AOI221xp5_ASAP7_75t_L g1029 ( .A1(n_564), .A2(n_1030), .B1(n_1031), .B2(n_1035), .C(n_1037), .Y(n_1029) );
INVx4_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g841 ( .A(n_566), .Y(n_841) );
INVx2_ASAP7_75t_L g950 ( .A(n_566), .Y(n_950) );
AOI31xp33_ASAP7_75t_L g614 ( .A1(n_567), .A2(n_615), .A3(n_627), .B(n_636), .Y(n_614) );
INVx5_ASAP7_75t_L g823 ( .A(n_567), .Y(n_823) );
AOI221x1_ASAP7_75t_SL g1236 ( .A1(n_567), .A2(n_1237), .B1(n_1271), .B2(n_1273), .C(n_1311), .Y(n_1236) );
BUFx8_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g1024 ( .A(n_568), .Y(n_1024) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx2_ASAP7_75t_L g722 ( .A(n_569), .Y(n_722) );
AND2x4_ASAP7_75t_L g1271 ( .A(n_569), .B(n_1272), .Y(n_1271) );
XOR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_637), .Y(n_570) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_612), .Y(n_572) );
NOR3xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_581), .C(n_585), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_578), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B1(n_591), .B2(n_592), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_588), .A2(n_600), .B1(n_601), .B2(n_603), .Y(n_599) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g1066 ( .A(n_589), .Y(n_1066) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx2_ASAP7_75t_L g669 ( .A(n_590), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_592), .A2(n_811), .B1(n_814), .B2(n_815), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_592), .A2(n_669), .B1(n_817), .B2(n_818), .Y(n_816) );
INVx2_ASAP7_75t_L g1428 ( .A(n_592), .Y(n_1428) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_596), .B1(n_597), .B2(n_598), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g906 ( .A(n_601), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_601), .A2(n_658), .B1(n_1191), .B2(n_1192), .Y(n_1190) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g664 ( .A(n_602), .Y(n_664) );
INVx2_ASAP7_75t_L g776 ( .A(n_602), .Y(n_776) );
INVx2_ASAP7_75t_L g898 ( .A(n_602), .Y(n_898) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_607), .B1(n_608), .B2(n_611), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g652 ( .A1(n_605), .A2(n_653), .B1(n_654), .B2(n_656), .Y(n_652) );
INVx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g805 ( .A1(n_608), .A2(n_806), .B1(n_808), .B2(n_809), .Y(n_805) );
OAI22xp33_ASAP7_75t_L g1845 ( .A1(n_608), .A2(n_1811), .B1(n_1823), .B2(n_1846), .Y(n_1845) );
BUFx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g655 ( .A(n_609), .Y(n_655) );
OAI22xp33_ASAP7_75t_L g1116 ( .A1(n_609), .A2(n_667), .B1(n_1090), .B2(n_1117), .Y(n_1116) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_609), .A2(n_667), .B1(n_1124), .B2(n_1125), .Y(n_1123) );
INVx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g987 ( .A(n_610), .Y(n_987) );
BUFx2_ASAP7_75t_L g1062 ( .A(n_610), .Y(n_1062) );
INVx2_ASAP7_75t_L g1277 ( .A(n_610), .Y(n_1277) );
INVx1_ASAP7_75t_L g1214 ( .A(n_621), .Y(n_1214) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx3_ASAP7_75t_L g1036 ( .A(n_622), .Y(n_1036) );
INVx1_ASAP7_75t_L g1408 ( .A(n_622), .Y(n_1408) );
INVx1_ASAP7_75t_L g1468 ( .A(n_622), .Y(n_1468) );
INVx2_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g845 ( .A(n_626), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_626), .A2(n_844), .B1(n_913), .B2(n_914), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g1470 ( .A1(n_626), .A2(n_1471), .B1(n_1472), .B2(n_1473), .Y(n_1470) );
HB1xp67_ASAP7_75t_L g1523 ( .A(n_630), .Y(n_1523) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI221xp5_ASAP7_75t_L g1215 ( .A1(n_632), .A2(n_1184), .B1(n_1189), .B2(n_1216), .C(n_1218), .Y(n_1215) );
INVx1_ASAP7_75t_L g1410 ( .A(n_632), .Y(n_1410) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_634), .A2(n_1192), .B1(n_1194), .B2(n_1200), .Y(n_1199) );
INVx4_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g1138 ( .A(n_635), .Y(n_1138) );
INVx1_ASAP7_75t_L g715 ( .A(n_638), .Y(n_715) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_676), .Y(n_638) );
NOR3xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_649), .C(n_651), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_645), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_643), .A2(n_887), .B1(n_888), .B2(n_889), .Y(n_886) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_644), .A2(n_646), .B1(n_691), .B2(n_694), .C(n_696), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g671 ( .A1(n_654), .A2(n_672), .B1(n_674), .B2(n_675), .Y(n_671) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B1(n_662), .B2(n_665), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g1115 ( .A(n_664), .Y(n_1115) );
OAI22xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_669), .B2(n_670), .Y(n_666) );
INVx1_ASAP7_75t_L g807 ( .A(n_667), .Y(n_807) );
INVx1_ASAP7_75t_L g1847 ( .A(n_667), .Y(n_1847) );
CKINVDCx5p33_ASAP7_75t_R g672 ( .A(n_673), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B(n_679), .Y(n_676) );
AOI31xp33_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_698), .A3(n_709), .B(n_710), .Y(n_679) );
INVx2_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g730 ( .A(n_689), .Y(n_730) );
INVx1_ASAP7_75t_L g1374 ( .A(n_689), .Y(n_1374) );
OAI221xp5_ASAP7_75t_L g1455 ( .A1(n_691), .A2(n_742), .B1(n_1456), .B2(n_1457), .C(n_1458), .Y(n_1455) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_SL g732 ( .A(n_692), .Y(n_732) );
BUFx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g870 ( .A(n_693), .Y(n_870) );
BUFx4f_ASAP7_75t_L g947 ( .A(n_693), .Y(n_947) );
INVx2_ASAP7_75t_L g955 ( .A(n_693), .Y(n_955) );
INVx1_ASAP7_75t_L g1217 ( .A(n_693), .Y(n_1217) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
BUFx2_ASAP7_75t_L g1518 ( .A(n_697), .Y(n_1518) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g1040 ( .A(n_703), .Y(n_1040) );
INVx2_ASAP7_75t_L g1910 ( .A(n_703), .Y(n_1910) );
INVx1_ASAP7_75t_L g1458 ( .A(n_705), .Y(n_1458) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g1454 ( .A(n_708), .Y(n_1454) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g1006 ( .A1(n_711), .A2(n_1007), .B1(n_1019), .B2(n_1020), .Y(n_1006) );
OAI31xp33_ASAP7_75t_L g1197 ( .A1(n_711), .A2(n_1198), .A3(n_1209), .B(n_1210), .Y(n_1197) );
CKINVDCx8_ASAP7_75t_R g711 ( .A(n_712), .Y(n_711) );
BUFx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g764 ( .A(n_713), .B(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g928 ( .A(n_713), .B(n_929), .Y(n_928) );
INVx2_ASAP7_75t_L g1105 ( .A(n_713), .Y(n_1105) );
OR2x6_ASAP7_75t_L g1314 ( .A(n_713), .B(n_1149), .Y(n_1314) );
AND2x4_ASAP7_75t_L g1382 ( .A(n_713), .B(n_765), .Y(n_1382) );
OR2x2_ASAP7_75t_L g1905 ( .A(n_713), .B(n_1906), .Y(n_1905) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
HB1xp67_ASAP7_75t_L g1071 ( .A(n_717), .Y(n_1071) );
XNOR2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_848), .Y(n_717) );
XOR2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_791), .Y(n_718) );
XNOR2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_790), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_752), .Y(n_720) );
INVx2_ASAP7_75t_L g878 ( .A(n_722), .Y(n_878) );
OAI31xp33_ASAP7_75t_L g941 ( .A1(n_722), .A2(n_942), .A3(n_943), .B(n_959), .Y(n_941) );
OAI31xp33_ASAP7_75t_SL g1451 ( .A1(n_722), .A2(n_1452), .A3(n_1459), .B(n_1463), .Y(n_1451) );
NAND3xp33_ASAP7_75t_SL g723 ( .A(n_724), .B(n_736), .C(n_748), .Y(n_723) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI21xp5_ASAP7_75t_SL g731 ( .A1(n_732), .A2(n_733), .B(n_734), .Y(n_731) );
BUFx3_ASAP7_75t_L g1821 ( .A(n_735), .Y(n_1821) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g1042 ( .A(n_738), .Y(n_1042) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
BUFx3_ASAP7_75t_L g1219 ( .A(n_743), .Y(n_1219) );
A2O1A1Ixp33_ASAP7_75t_SL g1464 ( .A1(n_744), .A2(n_1138), .B(n_1142), .C(n_1465), .Y(n_1464) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AND4x1_ASAP7_75t_L g752 ( .A(n_753), .B(n_763), .C(n_783), .D(n_786), .Y(n_752) );
AOI221xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_756), .B1(n_757), .B2(n_760), .C(n_761), .Y(n_753) );
AOI221xp5_ASAP7_75t_L g880 ( .A1(n_754), .A2(n_757), .B1(n_761), .B2(n_881), .C(n_882), .Y(n_880) );
AOI221xp5_ASAP7_75t_L g912 ( .A1(n_754), .A2(n_757), .B1(n_761), .B2(n_913), .C(n_914), .Y(n_912) );
AOI221xp5_ASAP7_75t_L g1126 ( .A1(n_754), .A2(n_757), .B1(n_761), .B2(n_1091), .C(n_1093), .Y(n_1126) );
AOI21xp5_ASAP7_75t_L g1170 ( .A1(n_754), .A2(n_761), .B(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1499 ( .A(n_754), .Y(n_1499) );
AOI221xp5_ASAP7_75t_L g1546 ( .A1(n_754), .A2(n_757), .B1(n_761), .B2(n_1547), .C(n_1548), .Y(n_1546) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_757), .A2(n_889), .B1(n_1137), .B2(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1497 ( .A(n_757), .Y(n_1497) );
AND2x4_ASAP7_75t_L g1882 ( .A(n_758), .B(n_1883), .Y(n_1882) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g1495 ( .A1(n_761), .A2(n_1472), .B1(n_1473), .B2(n_1496), .C(n_1498), .Y(n_1495) );
INVx1_ASAP7_75t_L g1345 ( .A(n_762), .Y(n_1345) );
HB1xp67_ASAP7_75t_L g1543 ( .A(n_762), .Y(n_1543) );
AOI33xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_766), .A3(n_772), .B1(n_774), .B2(n_777), .B3(n_782), .Y(n_763) );
AOI222xp33_ASAP7_75t_L g890 ( .A1(n_764), .A2(n_782), .B1(n_891), .B2(n_893), .C1(n_894), .C2(n_903), .Y(n_890) );
AOI33xp33_ASAP7_75t_L g915 ( .A1(n_764), .A2(n_916), .A3(n_921), .B1(n_925), .B2(n_927), .B3(n_928), .Y(n_915) );
AOI22xp5_ASAP7_75t_L g1118 ( .A1(n_764), .A2(n_889), .B1(n_1103), .B2(n_1119), .Y(n_1118) );
AOI322xp5_ASAP7_75t_L g1164 ( .A1(n_764), .A2(n_782), .A3(n_975), .B1(n_1151), .B2(n_1165), .C1(n_1166), .C2(n_1167), .Y(n_1164) );
NAND3xp33_ASAP7_75t_L g1892 ( .A(n_764), .B(n_1893), .C(n_1895), .Y(n_1892) );
AOI22xp5_ASAP7_75t_L g1110 ( .A1(n_767), .A2(n_1111), .B1(n_1112), .B2(n_1113), .Y(n_1110) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx3_ASAP7_75t_L g918 ( .A(n_768), .Y(n_918) );
BUFx2_ASAP7_75t_L g1384 ( .A(n_768), .Y(n_1384) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g1113 ( .A(n_770), .Y(n_1113) );
INVx2_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
HB1xp67_ASAP7_75t_L g1542 ( .A(n_773), .Y(n_1542) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_776), .A2(n_1028), .B1(n_1030), .B2(n_1066), .Y(n_1069) );
INVx2_ASAP7_75t_SL g1894 ( .A(n_776), .Y(n_1894) );
BUFx3_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g1005 ( .A(n_782), .Y(n_1005) );
AOI33xp33_ASAP7_75t_L g1380 ( .A1(n_782), .A2(n_1381), .A3(n_1383), .B1(n_1385), .B2(n_1391), .B3(n_1392), .Y(n_1380) );
AOI22xp5_ASAP7_75t_L g1438 ( .A1(n_782), .A2(n_785), .B1(n_1439), .B2(n_1446), .Y(n_1438) );
INVx2_ASAP7_75t_L g1489 ( .A(n_782), .Y(n_1489) );
XNOR2x1_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
AND2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_822), .Y(n_793) );
NOR3xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_802), .C(n_803), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_799), .Y(n_795) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
BUFx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g1838 ( .A1(n_812), .A2(n_1839), .B1(n_1840), .B2(n_1842), .Y(n_1838) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g991 ( .A(n_813), .Y(n_991) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_824), .B1(n_846), .B2(n_847), .Y(n_822) );
OAI21xp33_ASAP7_75t_L g1403 ( .A1(n_823), .A2(n_1404), .B(n_1417), .Y(n_1403) );
INVx1_ASAP7_75t_SL g1529 ( .A(n_823), .Y(n_1529) );
NAND3xp33_ASAP7_75t_L g824 ( .A(n_825), .B(n_830), .C(n_836), .Y(n_824) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AOI221xp5_ASAP7_75t_L g1008 ( .A1(n_828), .A2(n_995), .B1(n_1009), .B2(n_1010), .C(n_1011), .Y(n_1008) );
INVx1_ASAP7_75t_L g1133 ( .A(n_829), .Y(n_1133) );
BUFx2_ASAP7_75t_L g1373 ( .A(n_829), .Y(n_1373) );
INVx1_ASAP7_75t_L g1814 ( .A(n_829), .Y(n_1814) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g1228 ( .A(n_839), .Y(n_1228) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_SL g877 ( .A(n_844), .Y(n_877) );
INVx4_ASAP7_75t_L g1012 ( .A(n_844), .Y(n_1012) );
AOI21xp5_ASAP7_75t_L g1503 ( .A1(n_847), .A2(n_1504), .B(n_1505), .Y(n_1503) );
XOR2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_966), .Y(n_848) );
XNOR2x1_ASAP7_75t_L g849 ( .A(n_850), .B(n_909), .Y(n_849) );
NOR2x1_ASAP7_75t_L g851 ( .A(n_852), .B(n_879), .Y(n_851) );
AOI21xp5_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_866), .B(n_878), .Y(n_852) );
AOI221xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_857), .B1(n_859), .B2(n_861), .C(n_864), .Y(n_853) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g1034 ( .A(n_856), .Y(n_1034) );
INVx1_ASAP7_75t_L g1413 ( .A(n_856), .Y(n_1413) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g958 ( .A(n_864), .Y(n_958) );
AOI221xp5_ASAP7_75t_L g1038 ( .A1(n_864), .A2(n_1039), .B1(n_1041), .B2(n_1042), .C(n_1043), .Y(n_1038) );
BUFx3_ASAP7_75t_L g1142 ( .A(n_865), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx2_ASAP7_75t_SL g873 ( .A(n_874), .Y(n_873) );
INVx2_ASAP7_75t_L g1102 ( .A(n_876), .Y(n_1102) );
AOI31xp33_ASAP7_75t_L g1801 ( .A1(n_878), .A2(n_1802), .A3(n_1810), .B(n_1822), .Y(n_1801) );
NAND4xp25_ASAP7_75t_L g879 ( .A(n_880), .B(n_883), .C(n_886), .D(n_890), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_889), .A2(n_938), .B1(n_939), .B2(n_940), .Y(n_937) );
AOI22xp33_ASAP7_75t_SL g1493 ( .A1(n_889), .A2(n_1437), .B1(n_1465), .B2(n_1494), .Y(n_1493) );
AOI22xp5_ASAP7_75t_L g976 ( .A1(n_891), .A2(n_934), .B1(n_977), .B2(n_978), .Y(n_976) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_891), .A2(n_938), .B1(n_1161), .B2(n_1162), .Y(n_1160) );
INVx1_ASAP7_75t_L g1196 ( .A(n_891), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_892), .B(n_1297), .Y(n_1296) );
BUFx2_ASAP7_75t_L g1900 ( .A(n_892), .Y(n_1900) );
INVx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g1068 ( .A(n_897), .Y(n_1068) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
HB1xp67_ASAP7_75t_L g1844 ( .A(n_898), .Y(n_1844) );
INVx2_ASAP7_75t_SL g985 ( .A(n_901), .Y(n_985) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g1120 ( .A(n_905), .Y(n_1120) );
INVx1_ASAP7_75t_L g993 ( .A(n_906), .Y(n_993) );
NAND3xp33_ASAP7_75t_L g910 ( .A(n_911), .B(n_932), .C(n_941), .Y(n_910) );
AND3x1_ASAP7_75t_L g911 ( .A(n_912), .B(n_915), .C(n_930), .Y(n_911) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx3_ASAP7_75t_L g1292 ( .A(n_924), .Y(n_1292) );
OAI22xp5_ASAP7_75t_L g1479 ( .A1(n_924), .A2(n_990), .B1(n_1457), .B2(n_1480), .Y(n_1479) );
INVx2_ASAP7_75t_L g1898 ( .A(n_924), .Y(n_1898) );
BUFx3_ASAP7_75t_L g1386 ( .A(n_926), .Y(n_1386) );
INVx2_ASAP7_75t_SL g1285 ( .A(n_929), .Y(n_1285) );
AND2x2_ASAP7_75t_L g932 ( .A(n_933), .B(n_937), .Y(n_932) );
INVx1_ASAP7_75t_L g1157 ( .A(n_934), .Y(n_1157) );
INVx1_ASAP7_75t_L g1176 ( .A(n_934), .Y(n_1176) );
OAI211xp5_ASAP7_75t_L g953 ( .A1(n_936), .A2(n_954), .B(n_956), .C(n_957), .Y(n_953) );
AOI22xp5_ASAP7_75t_L g972 ( .A1(n_938), .A2(n_973), .B1(n_974), .B2(n_975), .Y(n_972) );
INVx2_ASAP7_75t_L g1179 ( .A(n_938), .Y(n_1179) );
NAND3xp33_ASAP7_75t_L g943 ( .A(n_944), .B(n_953), .C(n_958), .Y(n_943) );
OAI211xp5_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_946), .B(n_948), .C(n_951), .Y(n_944) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx2_ASAP7_75t_SL g1135 ( .A(n_947), .Y(n_1135) );
INVx2_ASAP7_75t_L g1807 ( .A(n_947), .Y(n_1807) );
INVx1_ASAP7_75t_L g1087 ( .A(n_949), .Y(n_1087) );
BUFx2_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx2_ASAP7_75t_L g964 ( .A(n_950), .Y(n_964) );
INVx2_ASAP7_75t_SL g1205 ( .A(n_952), .Y(n_1205) );
BUFx3_ASAP7_75t_L g1319 ( .A(n_952), .Y(n_1319) );
OAI211xp5_ASAP7_75t_L g1143 ( .A1(n_954), .A2(n_1144), .B(n_1145), .C(n_1146), .Y(n_1143) );
BUFx3_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g1153 ( .A(n_955), .Y(n_1153) );
INVx1_ASAP7_75t_L g1324 ( .A(n_964), .Y(n_1324) );
XNOR2xp5_ASAP7_75t_L g966 ( .A(n_967), .B(n_1021), .Y(n_966) );
XNOR2x1_ASAP7_75t_L g967 ( .A(n_968), .B(n_969), .Y(n_967) );
AND2x2_ASAP7_75t_L g969 ( .A(n_970), .B(n_1006), .Y(n_969) );
NOR3xp33_ASAP7_75t_L g970 ( .A(n_971), .B(n_979), .C(n_981), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_972), .B(n_976), .Y(n_971) );
OAI22xp33_ASAP7_75t_L g982 ( .A1(n_983), .A2(n_984), .B1(n_986), .B2(n_987), .Y(n_982) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVx2_ASAP7_75t_SL g1059 ( .A(n_985), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_989), .A2(n_990), .B1(n_992), .B2(n_993), .Y(n_988) );
BUFx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
OAI22xp5_ASAP7_75t_SL g994 ( .A1(n_995), .A2(n_996), .B1(n_997), .B2(n_998), .Y(n_994) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
HB1xp67_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1001), .Y(n_1310) );
NAND3xp33_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1013), .C(n_1018), .Y(n_1007) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1012), .Y(n_1471) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1046), .Y(n_1022) );
AOI22xp5_ASAP7_75t_L g1023 ( .A1(n_1024), .A2(n_1025), .B1(n_1044), .B2(n_1045), .Y(n_1023) );
NAND3xp33_ASAP7_75t_SL g1025 ( .A(n_1026), .B(n_1029), .C(n_1038), .Y(n_1025) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
NOR3xp33_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1055), .C(n_1057), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1052), .Y(n_1047) );
OAI22xp33_ASAP7_75t_L g1058 ( .A1(n_1059), .A2(n_1060), .B1(n_1061), .B2(n_1063), .Y(n_1058) );
OAI22xp33_ASAP7_75t_L g1835 ( .A1(n_1061), .A2(n_1443), .B1(n_1836), .B2(n_1837), .Y(n_1835) );
INVx2_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_1065), .A2(n_1066), .B1(n_1067), .B2(n_1068), .Y(n_1064) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
XNOR2xp5_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1396), .Y(n_1073) );
XOR2xp5_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1232), .Y(n_1074) );
HB1xp67_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
OAI22x1_ASAP7_75t_L g1076 ( .A1(n_1077), .A2(n_1078), .B1(n_1172), .B2(n_1231), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
XNOR2x1_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1127), .Y(n_1078) );
XNOR2x1_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1081), .Y(n_1079) );
OR2x2_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1106), .Y(n_1081) );
AOI31xp33_ASAP7_75t_SL g1082 ( .A1(n_1083), .A2(n_1094), .A3(n_1098), .B(n_1104), .Y(n_1082) );
INVx2_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVx2_ASAP7_75t_L g1132 ( .A(n_1086), .Y(n_1132) );
HB1xp67_ASAP7_75t_L g1213 ( .A(n_1086), .Y(n_1213) );
INVx2_ASAP7_75t_L g1226 ( .A(n_1086), .Y(n_1226) );
INVx3_ASAP7_75t_L g1511 ( .A(n_1092), .Y(n_1511) );
INVxp67_ASAP7_75t_L g1222 ( .A(n_1097), .Y(n_1222) );
AOI22xp5_ASAP7_75t_L g1098 ( .A1(n_1099), .A2(n_1100), .B1(n_1102), .B2(n_1103), .Y(n_1098) );
BUFx2_ASAP7_75t_L g1371 ( .A(n_1101), .Y(n_1371) );
INVx2_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
AOI211xp5_ASAP7_75t_L g1128 ( .A1(n_1105), .A2(n_1129), .B(n_1156), .C(n_1163), .Y(n_1128) );
NAND3xp33_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1118), .C(n_1126), .Y(n_1106) );
INVxp67_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
NAND4xp25_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1136), .C(n_1143), .D(n_1150), .Y(n_1129) );
A2O1A1Ixp33_ASAP7_75t_L g1136 ( .A1(n_1137), .A2(n_1138), .B(n_1139), .C(n_1142), .Y(n_1136) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
OAI211xp5_ASAP7_75t_L g1150 ( .A1(n_1151), .A2(n_1152), .B(n_1154), .C(n_1155), .Y(n_1150) );
OAI221xp5_ASAP7_75t_L g1315 ( .A1(n_1152), .A2(n_1226), .B1(n_1316), .B2(n_1317), .C(n_1318), .Y(n_1315) );
OAI221xp5_ASAP7_75t_L g1322 ( .A1(n_1152), .A2(n_1212), .B1(n_1298), .B2(n_1303), .C(n_1323), .Y(n_1322) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1170), .Y(n_1163) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1172), .Y(n_1231) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1173), .Y(n_1229) );
NAND3xp33_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1180), .C(n_1197), .Y(n_1173) );
NOR2xp33_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1178), .Y(n_1174) );
NOR2xp33_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1182), .Y(n_1180) );
OAI22xp5_ASAP7_75t_L g1211 ( .A1(n_1185), .A2(n_1187), .B1(n_1212), .B2(n_1214), .Y(n_1211) );
OAI22xp33_ASAP7_75t_L g1476 ( .A1(n_1188), .A2(n_1456), .B1(n_1477), .B2(n_1478), .Y(n_1476) );
OAI22xp33_ASAP7_75t_L g1486 ( .A1(n_1188), .A2(n_1445), .B1(n_1487), .B2(n_1488), .Y(n_1486) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_1191), .A2(n_1195), .B1(n_1204), .B2(n_1206), .Y(n_1203) );
BUFx2_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
INVx2_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
BUFx2_ASAP7_75t_SL g1206 ( .A(n_1207), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g1338 ( .A(n_1207), .Y(n_1338) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_1211), .A2(n_1215), .B1(n_1220), .B2(n_1224), .Y(n_1210) );
OAI21xp5_ASAP7_75t_SL g1514 ( .A1(n_1212), .A2(n_1515), .B(n_1516), .Y(n_1514) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
OAI221xp5_ASAP7_75t_L g1224 ( .A1(n_1216), .A2(n_1225), .B1(n_1226), .B2(n_1227), .C(n_1228), .Y(n_1224) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1216), .Y(n_1517) );
BUFx2_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_1233), .A2(n_1234), .B1(n_1325), .B2(n_1395), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
NAND4xp25_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1244), .C(n_1253), .D(n_1265), .Y(n_1237) );
BUFx2_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
NAND4xp25_ASAP7_75t_L g1328 ( .A(n_1239), .B(n_1329), .C(n_1333), .D(n_1336), .Y(n_1328) );
INVx5_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_1245), .A2(n_1246), .B1(n_1249), .B2(n_1250), .Y(n_1244) );
AOI222xp33_ASAP7_75t_L g1294 ( .A1(n_1245), .A2(n_1295), .B1(n_1298), .B2(n_1299), .C1(n_1303), .C2(n_1304), .Y(n_1294) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_1246), .A2(n_1250), .B1(n_1334), .B2(n_1335), .Y(n_1333) );
AOI221xp5_ASAP7_75t_L g1864 ( .A1(n_1246), .A2(n_1270), .B1(n_1865), .B2(n_1866), .C(n_1867), .Y(n_1864) );
AND2x4_ASAP7_75t_L g1260 ( .A(n_1247), .B(n_1261), .Y(n_1260) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1860 ( .A1(n_1250), .A2(n_1861), .B1(n_1862), .B2(n_1863), .Y(n_1860) );
AND2x4_ASAP7_75t_L g1267 ( .A(n_1251), .B(n_1268), .Y(n_1267) );
AND2x4_ASAP7_75t_L g1861 ( .A(n_1251), .B(n_1268), .Y(n_1861) );
INVx1_ASAP7_75t_SL g1251 ( .A(n_1252), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1869 ( .A(n_1252), .B(n_1870), .Y(n_1869) );
AOI222xp33_ASAP7_75t_L g1253 ( .A1(n_1254), .A2(n_1255), .B1(n_1258), .B2(n_1259), .C1(n_1263), .C2(n_1264), .Y(n_1253) );
OAI21xp5_ASAP7_75t_SL g1281 ( .A1(n_1254), .A2(n_1282), .B(n_1284), .Y(n_1281) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
AOI222xp33_ASAP7_75t_L g1336 ( .A1(n_1259), .A2(n_1264), .B1(n_1337), .B2(n_1338), .C1(n_1339), .C2(n_1340), .Y(n_1336) );
BUFx4f_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
INVx1_ASAP7_75t_L g1870 ( .A(n_1262), .Y(n_1870) );
INVx3_ASAP7_75t_L g1871 ( .A(n_1264), .Y(n_1871) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_1266), .A2(n_1267), .B1(n_1269), .B2(n_1270), .Y(n_1265) );
HB1xp67_ASAP7_75t_L g1331 ( .A(n_1267), .Y(n_1331) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_1270), .A2(n_1330), .B1(n_1331), .B2(n_1332), .Y(n_1329) );
AO211x2_ASAP7_75t_L g1327 ( .A1(n_1271), .A2(n_1328), .B(n_1341), .C(n_1367), .Y(n_1327) );
BUFx6f_ASAP7_75t_L g1874 ( .A(n_1271), .Y(n_1874) );
NAND3xp33_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1294), .C(n_1305), .Y(n_1273) );
NOR3xp33_ASAP7_75t_SL g1274 ( .A(n_1275), .B(n_1280), .C(n_1286), .Y(n_1274) );
INVx2_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
OR2x6_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1278), .Y(n_1276) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1277), .Y(n_1283) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1278), .Y(n_1288) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1278), .Y(n_1297) );
INVx2_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1283), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1293), .Y(n_1290) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1292), .Y(n_1484) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
AND2x4_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1302), .Y(n_1299) );
AND2x4_ASAP7_75t_L g1309 ( .A(n_1300), .B(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
AOI22xp33_ASAP7_75t_L g1305 ( .A1(n_1306), .A2(n_1307), .B1(n_1308), .B2(n_1309), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g1311 ( .A1(n_1312), .A2(n_1315), .B1(n_1320), .B2(n_1322), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
INVx2_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
CKINVDCx5p33_ASAP7_75t_R g1369 ( .A(n_1314), .Y(n_1369) );
INVx4_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
BUFx4f_ASAP7_75t_L g1379 ( .A(n_1321), .Y(n_1379) );
HB1xp67_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
INVxp67_ASAP7_75t_SL g1395 ( .A(n_1326), .Y(n_1395) );
INVx2_ASAP7_75t_L g1394 ( .A(n_1327), .Y(n_1394) );
AOI22xp33_ASAP7_75t_SL g1361 ( .A1(n_1334), .A2(n_1362), .B1(n_1363), .B2(n_1364), .Y(n_1361) );
AOI31xp33_ASAP7_75t_L g1341 ( .A1(n_1342), .A2(n_1353), .A3(n_1361), .B(n_1366), .Y(n_1341) );
AOI211xp5_ASAP7_75t_L g1342 ( .A1(n_1343), .A2(n_1344), .B(n_1346), .C(n_1349), .Y(n_1342) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1885 ( .A(n_1345), .Y(n_1885) );
CKINVDCx11_ASAP7_75t_R g1888 ( .A(n_1346), .Y(n_1888) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVxp67_ASAP7_75t_L g1883 ( .A(n_1348), .Y(n_1883) );
INVx2_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
AOI222xp33_ASAP7_75t_L g1879 ( .A1(n_1351), .A2(n_1880), .B1(n_1881), .B2(n_1882), .C1(n_1884), .C2(n_1885), .Y(n_1879) );
AOI22xp33_ASAP7_75t_SL g1353 ( .A1(n_1354), .A2(n_1356), .B1(n_1357), .B2(n_1360), .Y(n_1353) );
AOI22xp33_ASAP7_75t_L g1876 ( .A1(n_1354), .A2(n_1357), .B1(n_1877), .B2(n_1878), .Y(n_1876) );
AND2x4_ASAP7_75t_L g1357 ( .A(n_1355), .B(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
HB1xp67_ASAP7_75t_L g1390 ( .A(n_1359), .Y(n_1390) );
AOI22xp33_ASAP7_75t_L g1886 ( .A1(n_1362), .A2(n_1364), .B1(n_1865), .B2(n_1887), .Y(n_1886) );
INVx4_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1380), .Y(n_1367) );
AOI33xp33_ASAP7_75t_L g1368 ( .A1(n_1369), .A2(n_1370), .A3(n_1372), .B1(n_1375), .B2(n_1376), .B3(n_1379), .Y(n_1368) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
BUFx3_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
INVx2_ASAP7_75t_L g1539 ( .A(n_1382), .Y(n_1539) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
HB1xp67_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
BUFx3_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
AOI22xp5_ASAP7_75t_L g1398 ( .A1(n_1399), .A2(n_1400), .B1(n_1500), .B2(n_1549), .Y(n_1398) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
XNOR2xp5_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1449), .Y(n_1400) );
INVx2_ASAP7_75t_SL g1448 ( .A(n_1402), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1403), .B(n_1424), .Y(n_1402) );
AOI22xp5_ASAP7_75t_L g1405 ( .A1(n_1406), .A2(n_1409), .B1(n_1411), .B2(n_1412), .Y(n_1405) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
OAI22xp33_ASAP7_75t_L g1442 ( .A1(n_1415), .A2(n_1443), .B1(n_1444), .B2(n_1445), .Y(n_1442) );
CKINVDCx5p33_ASAP7_75t_R g1520 ( .A(n_1418), .Y(n_1520) );
NOR2xp33_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1433), .Y(n_1424) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1438), .Y(n_1433) );
INVx3_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
NAND4xp25_ASAP7_75t_L g1450 ( .A(n_1451), .B(n_1474), .C(n_1490), .D(n_1495), .Y(n_1450) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
NAND3xp33_ASAP7_75t_SL g1463 ( .A(n_1464), .B(n_1466), .C(n_1470), .Y(n_1463) );
OAI22xp5_ASAP7_75t_L g1481 ( .A1(n_1482), .A2(n_1483), .B1(n_1484), .B2(n_1485), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1491), .B(n_1493), .Y(n_1490) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
INVx2_ASAP7_75t_SL g1549 ( .A(n_1500), .Y(n_1549) );
XNOR2x1_ASAP7_75t_L g1500 ( .A(n_1501), .B(n_1502), .Y(n_1500) );
OAI22xp5_ASAP7_75t_L g1625 ( .A1(n_1501), .A2(n_1555), .B1(n_1626), .B2(n_1627), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1502 ( .A(n_1503), .B(n_1530), .Y(n_1502) );
AOI31xp33_ASAP7_75t_L g1505 ( .A1(n_1506), .A2(n_1519), .A3(n_1526), .B(n_1529), .Y(n_1505) );
AOI211xp5_ASAP7_75t_SL g1506 ( .A1(n_1507), .A2(n_1508), .B(n_1510), .C(n_1512), .Y(n_1506) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
AOI221xp5_ASAP7_75t_L g1519 ( .A1(n_1520), .A2(n_1521), .B1(n_1522), .B2(n_1524), .C(n_1525), .Y(n_1519) );
NOR2xp33_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1536), .Y(n_1530) );
NAND2xp5_ASAP7_75t_SL g1536 ( .A(n_1537), .B(n_1546), .Y(n_1536) );
INVx2_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
OAI221xp5_ASAP7_75t_L g1550 ( .A1(n_1551), .A2(n_1795), .B1(n_1797), .B2(n_1848), .C(n_1851), .Y(n_1550) );
AOI211xp5_ASAP7_75t_L g1551 ( .A1(n_1552), .A2(n_1578), .B(n_1708), .C(n_1762), .Y(n_1551) );
OAI321xp33_ASAP7_75t_L g1708 ( .A1(n_1552), .A2(n_1640), .A3(n_1709), .B1(n_1715), .B2(n_1719), .C(n_1734), .Y(n_1708) );
INVx3_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
AOI211xp5_ASAP7_75t_L g1734 ( .A1(n_1553), .A2(n_1735), .B(n_1749), .C(n_1758), .Y(n_1734) );
NAND2xp5_ASAP7_75t_L g1755 ( .A(n_1553), .B(n_1756), .Y(n_1755) );
INVx3_ASAP7_75t_L g1770 ( .A(n_1553), .Y(n_1770) );
NAND3xp33_ASAP7_75t_L g1776 ( .A(n_1553), .B(n_1612), .C(n_1670), .Y(n_1776) );
AND2x2_ASAP7_75t_L g1788 ( .A(n_1553), .B(n_1789), .Y(n_1788) );
INVx2_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
INVx2_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
AND2x4_ASAP7_75t_L g1556 ( .A(n_1557), .B(n_1559), .Y(n_1556) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1557), .Y(n_1563) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1558), .B(n_1571), .Y(n_1570) );
AND2x4_ASAP7_75t_L g1562 ( .A(n_1559), .B(n_1563), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1559), .B(n_1563), .Y(n_1602) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1560), .Y(n_1571) );
INVx1_ASAP7_75t_L g1796 ( .A(n_1561), .Y(n_1796) );
BUFx3_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1562), .Y(n_1626) );
HB1xp67_ASAP7_75t_L g1918 ( .A(n_1563), .Y(n_1918) );
OAI22xp33_ASAP7_75t_L g1564 ( .A1(n_1565), .A2(n_1566), .B1(n_1572), .B2(n_1573), .Y(n_1564) );
BUFx3_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
OAI22xp5_ASAP7_75t_L g1622 ( .A1(n_1567), .A2(n_1574), .B1(n_1623), .B2(n_1624), .Y(n_1622) );
BUFx6f_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
OAI22xp5_ASAP7_75t_L g1613 ( .A1(n_1568), .A2(n_1576), .B1(n_1614), .B2(n_1615), .Y(n_1613) );
OR2x2_ASAP7_75t_L g1568 ( .A(n_1569), .B(n_1570), .Y(n_1568) );
OR2x2_ASAP7_75t_L g1576 ( .A(n_1569), .B(n_1577), .Y(n_1576) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1569), .Y(n_1587) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1570), .Y(n_1586) );
HB1xp67_ASAP7_75t_L g1917 ( .A(n_1571), .Y(n_1917) );
HB1xp67_ASAP7_75t_L g1573 ( .A(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1577), .Y(n_1590) );
NAND4xp25_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1658), .C(n_1671), .D(n_1693), .Y(n_1578) );
NOR3xp33_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1645), .C(n_1650), .Y(n_1579) );
OAI211xp5_ASAP7_75t_L g1580 ( .A1(n_1581), .A2(n_1596), .B(n_1616), .C(n_1637), .Y(n_1580) );
OAI221xp5_ASAP7_75t_L g1735 ( .A1(n_1581), .A2(n_1713), .B1(n_1736), .B2(n_1744), .C(n_1745), .Y(n_1735) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
NAND2xp5_ASAP7_75t_L g1673 ( .A(n_1582), .B(n_1674), .Y(n_1673) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_1583), .B(n_1592), .Y(n_1582) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1583), .Y(n_1618) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1583), .Y(n_1636) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1583), .Y(n_1655) );
OR2x2_ASAP7_75t_L g1668 ( .A(n_1583), .B(n_1593), .Y(n_1668) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_1584), .B(n_1591), .Y(n_1583) );
AND2x4_ASAP7_75t_L g1585 ( .A(n_1586), .B(n_1587), .Y(n_1585) );
AND2x4_ASAP7_75t_L g1589 ( .A(n_1587), .B(n_1590), .Y(n_1589) );
BUFx2_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
OR2x2_ASAP7_75t_L g1635 ( .A(n_1592), .B(n_1636), .Y(n_1635) );
AND2x4_ASAP7_75t_L g1640 ( .A(n_1592), .B(n_1620), .Y(n_1640) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1592), .B(n_1621), .Y(n_1703) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1592), .Y(n_1722) );
NOR2xp33_ASAP7_75t_L g1729 ( .A(n_1592), .B(n_1730), .Y(n_1729) );
AOI221xp5_ASAP7_75t_L g1778 ( .A1(n_1592), .A2(n_1779), .B1(n_1781), .B2(n_1783), .C(n_1784), .Y(n_1778) );
INVx3_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_1593), .B(n_1620), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1657 ( .A(n_1593), .B(n_1621), .Y(n_1657) );
AND2x2_ASAP7_75t_L g1684 ( .A(n_1593), .B(n_1655), .Y(n_1684) );
AOI322xp5_ASAP7_75t_L g1693 ( .A1(n_1593), .A2(n_1598), .A3(n_1694), .B1(n_1696), .B2(n_1699), .C1(n_1702), .C2(n_1704), .Y(n_1693) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1594), .B(n_1595), .Y(n_1593) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
AND2x2_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1603), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1665 ( .A(n_1598), .B(n_1643), .Y(n_1665) );
OR2x2_ASAP7_75t_L g1679 ( .A(n_1598), .B(n_1605), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1701 ( .A(n_1598), .B(n_1612), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1720 ( .A(n_1598), .B(n_1721), .Y(n_1720) );
NOR2xp33_ASAP7_75t_L g1739 ( .A(n_1598), .B(n_1609), .Y(n_1739) );
AND2x2_ASAP7_75t_L g1742 ( .A(n_1598), .B(n_1609), .Y(n_1742) );
AND2x2_ASAP7_75t_L g1756 ( .A(n_1598), .B(n_1644), .Y(n_1756) );
BUFx3_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
BUFx2_ASAP7_75t_L g1632 ( .A(n_1599), .Y(n_1632) );
INVxp67_ASAP7_75t_L g1642 ( .A(n_1599), .Y(n_1642) );
OR2x2_ASAP7_75t_L g1728 ( .A(n_1599), .B(n_1612), .Y(n_1728) );
AND2x2_ASAP7_75t_L g1766 ( .A(n_1599), .B(n_1629), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1600), .B(n_1601), .Y(n_1599) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1604), .B(n_1608), .Y(n_1603) );
NOR2xp33_ASAP7_75t_L g1649 ( .A(n_1604), .B(n_1630), .Y(n_1649) );
NAND2xp5_ASAP7_75t_L g1695 ( .A(n_1604), .B(n_1640), .Y(n_1695) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1604), .B(n_1629), .Y(n_1721) );
OAI21xp5_ASAP7_75t_SL g1749 ( .A1(n_1604), .A2(n_1750), .B(n_1757), .Y(n_1749) );
AND2x2_ASAP7_75t_L g1773 ( .A(n_1604), .B(n_1688), .Y(n_1773) );
INVx2_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1617 ( .A(n_1605), .B(n_1618), .Y(n_1617) );
AND2x2_ASAP7_75t_L g1631 ( .A(n_1605), .B(n_1632), .Y(n_1631) );
BUFx2_ASAP7_75t_L g1661 ( .A(n_1605), .Y(n_1661) );
INVx2_ASAP7_75t_L g1670 ( .A(n_1605), .Y(n_1670) );
NAND2xp5_ASAP7_75t_L g1700 ( .A(n_1605), .B(n_1701), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1605), .B(n_1608), .Y(n_1711) );
A2O1A1Ixp33_ASAP7_75t_L g1723 ( .A1(n_1605), .A2(n_1656), .B(n_1724), .C(n_1726), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1730 ( .A(n_1605), .B(n_1620), .Y(n_1730) );
NAND2xp5_ASAP7_75t_L g1768 ( .A(n_1605), .B(n_1703), .Y(n_1768) );
NAND2xp5_ASAP7_75t_L g1780 ( .A(n_1605), .B(n_1725), .Y(n_1780) );
AND2x2_ASAP7_75t_L g1605 ( .A(n_1606), .B(n_1607), .Y(n_1605) );
NAND2xp5_ASAP7_75t_L g1718 ( .A(n_1608), .B(n_1631), .Y(n_1718) );
AND2x2_ASAP7_75t_L g1608 ( .A(n_1609), .B(n_1612), .Y(n_1608) );
OR2x2_ASAP7_75t_L g1630 ( .A(n_1609), .B(n_1612), .Y(n_1630) );
AND2x2_ASAP7_75t_L g1643 ( .A(n_1609), .B(n_1644), .Y(n_1643) );
INVx2_ASAP7_75t_L g1682 ( .A(n_1609), .Y(n_1682) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1610), .B(n_1611), .Y(n_1609) );
AOI32xp33_ASAP7_75t_L g1616 ( .A1(n_1612), .A2(n_1617), .A3(n_1619), .B1(n_1628), .B2(n_1633), .Y(n_1616) );
INVx2_ASAP7_75t_SL g1644 ( .A(n_1612), .Y(n_1644) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_1612), .B(n_1682), .Y(n_1688) );
NAND2xp5_ASAP7_75t_L g1663 ( .A(n_1618), .B(n_1664), .Y(n_1663) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1618), .B(n_1703), .Y(n_1702) );
O2A1O1Ixp33_ASAP7_75t_L g1767 ( .A1(n_1618), .A2(n_1682), .B(n_1718), .C(n_1768), .Y(n_1767) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1619), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1732 ( .A(n_1619), .B(n_1733), .Y(n_1732) );
INVx2_ASAP7_75t_SL g1634 ( .A(n_1620), .Y(n_1634) );
HB1xp67_ASAP7_75t_L g1646 ( .A(n_1620), .Y(n_1646) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1620), .Y(n_1674) );
AOI21xp5_ASAP7_75t_L g1736 ( .A1(n_1620), .A2(n_1737), .B(n_1740), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1743 ( .A(n_1620), .B(n_1670), .Y(n_1743) );
NAND2xp5_ASAP7_75t_L g1782 ( .A(n_1620), .B(n_1692), .Y(n_1782) );
OAI32xp33_ASAP7_75t_L g1786 ( .A1(n_1620), .A2(n_1634), .A3(n_1687), .B1(n_1721), .B2(n_1725), .Y(n_1786) );
CKINVDCx5p33_ASAP7_75t_R g1620 ( .A(n_1621), .Y(n_1620) );
OR2x2_ASAP7_75t_L g1621 ( .A(n_1622), .B(n_1625), .Y(n_1621) );
AND2x2_ASAP7_75t_L g1783 ( .A(n_1628), .B(n_1634), .Y(n_1783) );
AND2x2_ASAP7_75t_L g1628 ( .A(n_1629), .B(n_1631), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1629), .B(n_1642), .Y(n_1675) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1630), .Y(n_1629) );
OR2x2_ASAP7_75t_L g1678 ( .A(n_1630), .B(n_1679), .Y(n_1678) );
AND2x2_ASAP7_75t_L g1687 ( .A(n_1631), .B(n_1688), .Y(n_1687) );
NOR2xp33_ASAP7_75t_L g1681 ( .A(n_1632), .B(n_1682), .Y(n_1681) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1632), .B(n_1688), .Y(n_1707) );
NOR2x1_ASAP7_75t_L g1748 ( .A(n_1632), .B(n_1644), .Y(n_1748) );
NOR2xp33_ASAP7_75t_L g1633 ( .A(n_1634), .B(n_1635), .Y(n_1633) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1634), .Y(n_1664) );
INVx2_ASAP7_75t_L g1717 ( .A(n_1634), .Y(n_1717) );
NOR2xp33_ASAP7_75t_L g1746 ( .A(n_1635), .B(n_1747), .Y(n_1746) );
OAI22xp5_ASAP7_75t_L g1777 ( .A1(n_1635), .A2(n_1663), .B1(n_1689), .B2(n_1741), .Y(n_1777) );
INVxp67_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
A2O1A1Ixp33_ASAP7_75t_L g1757 ( .A1(n_1638), .A2(n_1694), .B(n_1713), .C(n_1727), .Y(n_1757) );
NOR2xp33_ASAP7_75t_L g1638 ( .A(n_1639), .B(n_1641), .Y(n_1638) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
AOI22xp5_ASAP7_75t_L g1750 ( .A1(n_1640), .A2(n_1751), .B1(n_1753), .B2(n_1754), .Y(n_1750) );
AND2x2_ASAP7_75t_L g1760 ( .A(n_1640), .B(n_1692), .Y(n_1760) );
INVx2_ASAP7_75t_L g1733 ( .A(n_1641), .Y(n_1733) );
NAND2xp5_ASAP7_75t_L g1641 ( .A(n_1642), .B(n_1643), .Y(n_1641) );
AND2x2_ASAP7_75t_L g1648 ( .A(n_1642), .B(n_1649), .Y(n_1648) );
AND2x2_ASAP7_75t_L g1710 ( .A(n_1642), .B(n_1711), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1725 ( .A(n_1642), .B(n_1688), .Y(n_1725) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1643), .Y(n_1651) );
NOR2xp33_ASAP7_75t_L g1645 ( .A(n_1646), .B(n_1647), .Y(n_1645) );
A2O1A1Ixp33_ASAP7_75t_L g1771 ( .A1(n_1647), .A2(n_1652), .B(n_1772), .C(n_1774), .Y(n_1771) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
NOR2xp33_ASAP7_75t_L g1650 ( .A(n_1651), .B(n_1652), .Y(n_1650) );
OR2x2_ASAP7_75t_L g1689 ( .A(n_1651), .B(n_1679), .Y(n_1689) );
NAND2xp5_ASAP7_75t_L g1697 ( .A(n_1651), .B(n_1698), .Y(n_1697) );
OR2x2_ASAP7_75t_L g1652 ( .A(n_1653), .B(n_1656), .Y(n_1652) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1654), .Y(n_1789) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1655), .Y(n_1692) );
AOI21xp5_ASAP7_75t_L g1758 ( .A1(n_1656), .A2(n_1759), .B(n_1761), .Y(n_1758) );
CKINVDCx5p33_ASAP7_75t_R g1656 ( .A(n_1657), .Y(n_1656) );
NAND2xp5_ASAP7_75t_L g1660 ( .A(n_1657), .B(n_1661), .Y(n_1660) );
O2A1O1Ixp33_ASAP7_75t_L g1658 ( .A1(n_1659), .A2(n_1662), .B(n_1665), .C(n_1666), .Y(n_1658) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
INVx2_ASAP7_75t_L g1706 ( .A(n_1661), .Y(n_1706) );
NAND2xp5_ASAP7_75t_SL g1738 ( .A(n_1661), .B(n_1739), .Y(n_1738) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
OR2x2_ASAP7_75t_L g1792 ( .A(n_1664), .B(n_1780), .Y(n_1792) );
AND2x2_ASAP7_75t_L g1669 ( .A(n_1665), .B(n_1670), .Y(n_1669) );
NOR2xp33_ASAP7_75t_L g1752 ( .A(n_1665), .B(n_1725), .Y(n_1752) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1667), .B(n_1669), .Y(n_1666) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1668), .Y(n_1667) );
NAND2xp5_ASAP7_75t_L g1680 ( .A(n_1670), .B(n_1681), .Y(n_1680) );
NAND2xp5_ASAP7_75t_L g1785 ( .A(n_1670), .B(n_1703), .Y(n_1785) );
AOI211xp5_ASAP7_75t_L g1671 ( .A1(n_1672), .A2(n_1675), .B(n_1676), .C(n_1685), .Y(n_1671) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1673), .Y(n_1672) );
NAND2xp5_ASAP7_75t_L g1683 ( .A(n_1674), .B(n_1684), .Y(n_1683) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1674), .B(n_1692), .Y(n_1691) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1674), .Y(n_1714) );
OAI22xp5_ASAP7_75t_L g1676 ( .A1(n_1677), .A2(n_1678), .B1(n_1680), .B2(n_1683), .Y(n_1676) );
OAI31xp33_ASAP7_75t_L g1790 ( .A1(n_1684), .A2(n_1720), .A3(n_1791), .B(n_1793), .Y(n_1790) );
AOI21xp33_ASAP7_75t_L g1685 ( .A1(n_1686), .A2(n_1689), .B(n_1690), .Y(n_1685) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1688), .Y(n_1698) );
NOR2xp33_ASAP7_75t_L g1764 ( .A(n_1690), .B(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
INVx2_ASAP7_75t_L g1713 ( .A(n_1692), .Y(n_1713) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
NAND2xp5_ASAP7_75t_L g1705 ( .A(n_1706), .B(n_1707), .Y(n_1705) );
NAND2xp5_ASAP7_75t_L g1747 ( .A(n_1706), .B(n_1748), .Y(n_1747) );
NAND2xp5_ASAP7_75t_L g1794 ( .A(n_1707), .B(n_1717), .Y(n_1794) );
AOI21xp33_ASAP7_75t_SL g1709 ( .A1(n_1710), .A2(n_1712), .B(n_1714), .Y(n_1709) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1711), .Y(n_1744) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1713), .Y(n_1712) );
INVxp67_ASAP7_75t_SL g1715 ( .A(n_1716), .Y(n_1715) );
NAND2xp5_ASAP7_75t_L g1716 ( .A(n_1717), .B(n_1718), .Y(n_1716) );
AOI211xp5_ASAP7_75t_L g1719 ( .A1(n_1720), .A2(n_1722), .B(n_1723), .C(n_1731), .Y(n_1719) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1720), .Y(n_1761) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1722), .Y(n_1753) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
O2A1O1Ixp33_ASAP7_75t_L g1774 ( .A1(n_1725), .A2(n_1760), .B(n_1775), .C(n_1777), .Y(n_1774) );
NAND2xp5_ASAP7_75t_L g1726 ( .A(n_1727), .B(n_1729), .Y(n_1726) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
INVxp67_ASAP7_75t_L g1731 ( .A(n_1732), .Y(n_1731) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1738), .Y(n_1737) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
NAND2xp5_ASAP7_75t_L g1741 ( .A(n_1742), .B(n_1743), .Y(n_1741) );
O2A1O1Ixp33_ASAP7_75t_SL g1784 ( .A1(n_1742), .A2(n_1785), .B(n_1786), .C(n_1787), .Y(n_1784) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1752), .Y(n_1751) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
NAND3xp33_ASAP7_75t_L g1762 ( .A(n_1763), .B(n_1778), .C(n_1790), .Y(n_1762) );
O2A1O1Ixp33_ASAP7_75t_L g1763 ( .A1(n_1764), .A2(n_1767), .B(n_1769), .C(n_1771), .Y(n_1763) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
INVx2_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
INVx1_ASAP7_75t_L g1772 ( .A(n_1773), .Y(n_1772) );
INVx1_ASAP7_75t_L g1775 ( .A(n_1776), .Y(n_1775) );
INVx1_ASAP7_75t_L g1779 ( .A(n_1780), .Y(n_1779) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1782), .Y(n_1781) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1788), .Y(n_1787) );
INVxp67_ASAP7_75t_L g1791 ( .A(n_1792), .Y(n_1791) );
INVxp67_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
HB1xp67_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
AND2x2_ASAP7_75t_L g1798 ( .A(n_1799), .B(n_1825), .Y(n_1798) );
OAI211xp5_ASAP7_75t_L g1805 ( .A1(n_1806), .A2(n_1807), .B(n_1808), .C(n_1809), .Y(n_1805) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1814), .Y(n_1813) );
HB1xp67_ASAP7_75t_L g1815 ( .A(n_1816), .Y(n_1815) );
INVx1_ASAP7_75t_L g1816 ( .A(n_1817), .Y(n_1816) );
INVx1_ASAP7_75t_L g1818 ( .A(n_1819), .Y(n_1818) );
NOR3xp33_ASAP7_75t_SL g1825 ( .A(n_1826), .B(n_1833), .C(n_1834), .Y(n_1825) );
NAND2xp5_ASAP7_75t_L g1826 ( .A(n_1827), .B(n_1830), .Y(n_1826) );
INVx1_ASAP7_75t_L g1840 ( .A(n_1841), .Y(n_1840) );
INVx1_ASAP7_75t_L g1846 ( .A(n_1847), .Y(n_1846) );
CKINVDCx5p33_ASAP7_75t_R g1848 ( .A(n_1849), .Y(n_1848) );
A2O1A1Ixp33_ASAP7_75t_L g1915 ( .A1(n_1850), .A2(n_1916), .B(n_1918), .C(n_1919), .Y(n_1915) );
BUFx2_ASAP7_75t_L g1852 ( .A(n_1853), .Y(n_1852) );
INVx1_ASAP7_75t_L g1853 ( .A(n_1854), .Y(n_1853) );
INVx1_ASAP7_75t_L g1854 ( .A(n_1855), .Y(n_1854) );
HB1xp67_ASAP7_75t_L g1856 ( .A(n_1857), .Y(n_1856) );
INVx1_ASAP7_75t_L g1913 ( .A(n_1858), .Y(n_1913) );
AOI221x1_ASAP7_75t_L g1858 ( .A1(n_1859), .A2(n_1874), .B1(n_1875), .B2(n_1889), .C(n_1891), .Y(n_1858) );
NAND2xp5_ASAP7_75t_L g1859 ( .A(n_1860), .B(n_1864), .Y(n_1859) );
INVx1_ASAP7_75t_L g1868 ( .A(n_1869), .Y(n_1868) );
NAND4xp25_ASAP7_75t_SL g1875 ( .A(n_1876), .B(n_1879), .C(n_1886), .D(n_1888), .Y(n_1875) );
CKINVDCx16_ASAP7_75t_R g1889 ( .A(n_1890), .Y(n_1889) );
NAND4xp25_ASAP7_75t_L g1891 ( .A(n_1892), .B(n_1896), .C(n_1901), .D(n_1907), .Y(n_1891) );
NAND3xp33_ASAP7_75t_L g1901 ( .A(n_1902), .B(n_1903), .C(n_1904), .Y(n_1901) );
INVx3_ASAP7_75t_L g1904 ( .A(n_1905), .Y(n_1904) );
NAND3xp33_ASAP7_75t_L g1907 ( .A(n_1908), .B(n_1909), .C(n_1911), .Y(n_1907) );
HB1xp67_ASAP7_75t_L g1914 ( .A(n_1915), .Y(n_1914) );
INVx1_ASAP7_75t_L g1916 ( .A(n_1917), .Y(n_1916) );
endmodule