module fake_jpeg_21138_n_409 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_409);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_409;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_49),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_71),
.Y(n_105)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_56),
.Y(n_116)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_58),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_59),
.B(n_64),
.Y(n_143)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_25),
.B(n_0),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_66),
.A2(n_90),
.B(n_2),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx2_ASAP7_75t_SL g95 ( 
.A(n_68),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_69),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_20),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_70),
.B(n_84),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_28),
.B(n_33),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_75),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_15),
.Y(n_77)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_17),
.B(n_27),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_85),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_21),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_40),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_17),
.B(n_0),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_24),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_3),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_27),
.B1(n_44),
.B2(n_39),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_92),
.A2(n_129),
.B1(n_29),
.B2(n_36),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_96),
.A2(n_128),
.B(n_3),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_51),
.A2(n_40),
.B1(n_31),
.B2(n_39),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_98),
.A2(n_112),
.B1(n_68),
.B2(n_48),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_127),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_62),
.A2(n_40),
.B1(n_44),
.B2(n_42),
.Y(n_112)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g129 ( 
.A1(n_81),
.A2(n_42),
.B1(n_36),
.B2(n_35),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_133),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_132),
.B(n_50),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_75),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_77),
.Y(n_173)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_150),
.B(n_170),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_52),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_154),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_152),
.A2(n_155),
.B1(n_161),
.B2(n_166),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

BUFx4f_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_55),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_66),
.B1(n_60),
.B2(n_90),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_156),
.A2(n_122),
.B1(n_114),
.B2(n_117),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_104),
.A2(n_83),
.B1(n_68),
.B2(n_29),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_115),
.A2(n_83),
.B1(n_73),
.B2(n_86),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_112),
.A2(n_63),
.B1(n_32),
.B2(n_30),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_164),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_47),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_154),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_94),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_165),
.B(n_168),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_98),
.A2(n_35),
.B1(n_34),
.B2(n_32),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_79),
.B1(n_26),
.B2(n_34),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_143),
.B(n_30),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_125),
.A2(n_80),
.B1(n_89),
.B2(n_45),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_171),
.A2(n_188),
.B1(n_149),
.B2(n_146),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_172),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_178),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_121),
.B(n_56),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_136),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

BUFx8_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_101),
.B(n_26),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_119),
.B(n_56),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_67),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_103),
.B(n_99),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_140),
.A2(n_76),
.B1(n_72),
.B2(n_69),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_93),
.Y(n_189)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_190),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_193),
.A2(n_195),
.B(n_199),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_46),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_148),
.A2(n_141),
.B1(n_117),
.B2(n_123),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_103),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_124),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_209),
.B1(n_213),
.B2(n_175),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_163),
.A2(n_123),
.B(n_139),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_136),
.B(n_124),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_151),
.A2(n_135),
.B1(n_110),
.B2(n_106),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_218),
.A2(n_116),
.B1(n_189),
.B2(n_147),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_171),
.A2(n_175),
.B1(n_177),
.B2(n_179),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_221),
.A2(n_181),
.B1(n_190),
.B2(n_186),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_158),
.B(n_160),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_193),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_229),
.A2(n_232),
.B1(n_234),
.B2(n_238),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_164),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_247),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_204),
.A2(n_187),
.B1(n_183),
.B2(n_176),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_221),
.B1(n_224),
.B2(n_218),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_180),
.B1(n_157),
.B2(n_162),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_193),
.A2(n_148),
.B1(n_180),
.B2(n_157),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_169),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_236),
.B(n_239),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_172),
.B1(n_168),
.B2(n_165),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_237),
.A2(n_231),
.B1(n_202),
.B2(n_251),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_206),
.A2(n_174),
.B1(n_106),
.B2(n_110),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_192),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_240),
.B(n_251),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_201),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_249),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_242),
.A2(n_235),
.B(n_249),
.Y(n_281)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_3),
.C(n_4),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_4),
.B(n_5),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_196),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_194),
.A2(n_116),
.B1(n_169),
.B2(n_153),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_258),
.B1(n_234),
.B2(n_229),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_212),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_219),
.A2(n_224),
.B1(n_198),
.B2(n_215),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_191),
.C(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_200),
.Y(n_252)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_259),
.Y(n_276)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_255),
.Y(n_280)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_256),
.B(n_257),
.Y(n_289)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_208),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_199),
.B(n_147),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_198),
.B(n_147),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_260),
.A2(n_226),
.B(n_211),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_261),
.A2(n_270),
.B1(n_277),
.B2(n_283),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_263),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_219),
.B1(n_205),
.B2(n_213),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_236),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_242),
.A2(n_195),
.B1(n_214),
.B2(n_222),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_232),
.A2(n_195),
.B1(n_222),
.B2(n_216),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_227),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_253),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_250),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_255),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_281),
.A2(n_286),
.B(n_288),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_287),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_238),
.A2(n_216),
.B1(n_202),
.B2(n_223),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_246),
.B1(n_240),
.B2(n_231),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_249),
.A2(n_226),
.B(n_223),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_253),
.A2(n_211),
.B(n_228),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_292),
.B(n_283),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_293),
.A2(n_299),
.B1(n_300),
.B2(n_309),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_254),
.C(n_259),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_303),
.C(n_304),
.Y(n_319)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_296),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_237),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_297),
.B(n_298),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_254),
.B1(n_247),
.B2(n_252),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_269),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_301),
.B(n_302),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_230),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_256),
.C(n_243),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_203),
.C(n_257),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_272),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_310),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_265),
.A2(n_245),
.B1(n_228),
.B2(n_203),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_245),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_311),
.Y(n_324)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_312),
.A2(n_314),
.B1(n_268),
.B2(n_289),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_286),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_88),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_211),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_276),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_315),
.B(n_320),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_297),
.A2(n_271),
.B1(n_265),
.B2(n_266),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_316),
.A2(n_317),
.B1(n_325),
.B2(n_332),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_297),
.A2(n_271),
.B1(n_266),
.B2(n_282),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_281),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_288),
.C(n_274),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_323),
.B(n_326),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_308),
.A2(n_279),
.B1(n_273),
.B2(n_267),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_284),
.C(n_280),
.Y(n_326)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_328),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_329),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_287),
.C(n_211),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_330),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_308),
.A2(n_196),
.B1(n_5),
.B2(n_6),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_294),
.A2(n_196),
.B1(n_7),
.B2(n_9),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_334),
.A2(n_335),
.B1(n_309),
.B2(n_299),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_290),
.A2(n_4),
.B1(n_7),
.B2(n_9),
.Y(n_335)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_336),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_321),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_338),
.B(n_347),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_318),
.A2(n_301),
.B1(n_290),
.B2(n_298),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_340),
.A2(n_350),
.B1(n_293),
.B2(n_306),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_322),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_348),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_327),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_348),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_335),
.A2(n_307),
.B1(n_333),
.B2(n_325),
.Y(n_346)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_346),
.Y(n_366)
);

INVx6_ASAP7_75t_L g347 ( 
.A(n_334),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_324),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_352),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_329),
.A2(n_312),
.B1(n_296),
.B2(n_291),
.Y(n_350)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_331),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_317),
.Y(n_353)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_353),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_341),
.A2(n_316),
.B(n_306),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_355),
.A2(n_337),
.B(n_345),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_357),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_354),
.B(n_326),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_351),
.B(n_319),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_358),
.B(n_343),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_344),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_352),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_319),
.C(n_330),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_369),
.C(n_340),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_320),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g378 ( 
.A(n_363),
.B(n_367),
.C(n_347),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_315),
.Y(n_367)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_368),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_342),
.B(n_323),
.C(n_336),
.Y(n_369)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_370),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_378),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_372),
.B(n_379),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_355),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_337),
.C(n_349),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_380),
.C(n_356),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_365),
.B(n_305),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_375),
.B(n_366),
.Y(n_386)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_368),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_311),
.C(n_332),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_82),
.C(n_10),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_7),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_376),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_384),
.A2(n_387),
.B1(n_381),
.B2(n_382),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_363),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_385),
.B(n_386),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_374),
.A2(n_369),
.B1(n_364),
.B2(n_360),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_384),
.A2(n_377),
.B1(n_364),
.B2(n_361),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_392),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_388),
.A2(n_378),
.B1(n_361),
.B2(n_359),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_396),
.C(n_387),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_389),
.A2(n_359),
.B1(n_311),
.B2(n_97),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_394),
.B(n_383),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_395),
.A2(n_9),
.B(n_10),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_397),
.A2(n_396),
.B(n_390),
.Y(n_401)
);

NOR3xp33_ASAP7_75t_L g402 ( 
.A(n_399),
.B(n_395),
.C(n_394),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_400),
.B(n_385),
.C(n_12),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_401),
.A2(n_403),
.B(n_398),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_402),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_405),
.B(n_11),
.Y(n_406)
);

A2O1A1Ixp33_ASAP7_75t_L g407 ( 
.A1(n_406),
.A2(n_404),
.B(n_12),
.C(n_13),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_407),
.A2(n_11),
.B(n_404),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_11),
.Y(n_409)
);


endmodule