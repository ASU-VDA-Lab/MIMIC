module fake_ariane_3034_n_2061 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2061);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2061;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_212;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g208 ( 
.A(n_17),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_22),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_69),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_95),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_123),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_29),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_36),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_14),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_93),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_40),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_180),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_57),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_154),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_18),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_2),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_19),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_103),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_98),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_53),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_10),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_8),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_128),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_191),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_104),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_120),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_124),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_22),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_86),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_41),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_81),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_142),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_41),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_198),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_207),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_177),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_97),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_170),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_158),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_71),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_141),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_45),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_42),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_132),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_202),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_7),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_28),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_20),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_51),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_160),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_60),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_94),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_19),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_6),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_72),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_149),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_115),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_125),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_96),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_148),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_109),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_189),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_143),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_179),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_9),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_164),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_201),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_113),
.Y(n_281)
);

INVxp33_ASAP7_75t_SL g282 ( 
.A(n_10),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_1),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_31),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_182),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_138),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_21),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_52),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_134),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_20),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_129),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_181),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_54),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_167),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_60),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_192),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_206),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_161),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_51),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_30),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_64),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_150),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_77),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_25),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_47),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_13),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_89),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_147),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_63),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_48),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_38),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_186),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_25),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_5),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_13),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_122),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_18),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_45),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_12),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_57),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_28),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_63),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_90),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_187),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_99),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_0),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_88),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_65),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_34),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_49),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_146),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_46),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_33),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_70),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_169),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_157),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_155),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_14),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_81),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_61),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_64),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_75),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_84),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_26),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_204),
.Y(n_345)
);

INVx4_ASAP7_75t_R g346 ( 
.A(n_72),
.Y(n_346)
);

CKINVDCx11_ASAP7_75t_R g347 ( 
.A(n_117),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_140),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_116),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_197),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_86),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_190),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_106),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_172),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_61),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_153),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_17),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_32),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_92),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_77),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_11),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_108),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_184),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_46),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_183),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_193),
.B(n_119),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_136),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_114),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_130),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_165),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_131),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_156),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_31),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_80),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_121),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_79),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_101),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_44),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_162),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_151),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_40),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_139),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_185),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_196),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_133),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_24),
.Y(n_386)
);

BUFx8_ASAP7_75t_SL g387 ( 
.A(n_145),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_105),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_152),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_135),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_66),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_26),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_107),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_66),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_58),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_100),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_175),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_91),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_118),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_137),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_222),
.Y(n_401)
);

INVxp33_ASAP7_75t_SL g402 ( 
.A(n_339),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_391),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_254),
.Y(n_404)
);

INVxp33_ASAP7_75t_SL g405 ( 
.A(n_339),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_355),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_254),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_323),
.B(n_0),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_387),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_347),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_254),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_272),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_323),
.B(n_1),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_254),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_254),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_296),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_349),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_356),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_362),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_383),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_282),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_394),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_262),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_210),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_311),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_266),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_309),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_215),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_217),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_254),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_355),
.Y(n_431)
);

INVxp33_ASAP7_75t_SL g432 ( 
.A(n_220),
.Y(n_432)
);

BUFx6f_ASAP7_75t_SL g433 ( 
.A(n_307),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_352),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g435 ( 
.A(n_295),
.B(n_2),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_223),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_254),
.B(n_3),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_228),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_233),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_234),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_254),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_254),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_240),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_218),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_242),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_218),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_219),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_301),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_243),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_219),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_321),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_229),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_311),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_229),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_245),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_374),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_358),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_208),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_252),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_352),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_256),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_260),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_365),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_301),
.Y(n_464)
);

INVxp33_ASAP7_75t_SL g465 ( 
.A(n_267),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_230),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_230),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_365),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_250),
.B(n_3),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_250),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_307),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_251),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_307),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_251),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_208),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_400),
.B(n_253),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_253),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_268),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_255),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_307),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_255),
.B(n_4),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_273),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_222),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_273),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_283),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_275),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_287),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_275),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_209),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_276),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_301),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_276),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_300),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_271),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_281),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_209),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_281),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_374),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_289),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_289),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_303),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_271),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_292),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_292),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_297),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_297),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_353),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_304),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_491),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_408),
.B(n_301),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_491),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_491),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_491),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_404),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_404),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_413),
.B(n_301),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_407),
.Y(n_517)
);

AND3x2_ASAP7_75t_L g518 ( 
.A(n_406),
.B(n_431),
.C(n_456),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_401),
.B(n_295),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_407),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_448),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_448),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_411),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_476),
.B(n_308),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_411),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_414),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_464),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_414),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_415),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_415),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_430),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_430),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_401),
.B(n_444),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_464),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_441),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_433),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_442),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_444),
.B(n_290),
.Y(n_540)
);

OA21x2_ASAP7_75t_L g541 ( 
.A1(n_437),
.A2(n_316),
.B(n_308),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_446),
.B(n_290),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_446),
.B(n_329),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_447),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_447),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_450),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_450),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_433),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_452),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_452),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_454),
.B(n_329),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_454),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_466),
.B(n_316),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_466),
.B(n_335),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

BUFx8_ASAP7_75t_L g557 ( 
.A(n_433),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_467),
.B(n_335),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_470),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_433),
.B(n_434),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_470),
.B(n_336),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_472),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_472),
.B(n_336),
.Y(n_563)
);

OA21x2_ASAP7_75t_L g564 ( 
.A1(n_474),
.A2(n_354),
.B(n_348),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_474),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_477),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_477),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_501),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_479),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_498),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_479),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_482),
.B(n_257),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_401),
.B(n_333),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_482),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_484),
.B(n_333),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_434),
.B(n_392),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_484),
.B(n_348),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_468),
.B(n_392),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_486),
.B(n_338),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_486),
.B(n_354),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_488),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_488),
.B(n_359),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_490),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_490),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_425),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_492),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_492),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_460),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_495),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_423),
.A2(n_360),
.B1(n_225),
.B2(n_227),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_495),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_497),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_497),
.Y(n_593)
);

AND2x2_ASAP7_75t_R g594 ( 
.A(n_463),
.B(n_346),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_412),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_499),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_499),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_570),
.B(n_468),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_557),
.Y(n_599)
);

BUFx4f_ASAP7_75t_L g600 ( 
.A(n_541),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_537),
.Y(n_601)
);

NOR2x1p5_ASAP7_75t_L g602 ( 
.A(n_595),
.B(n_409),
.Y(n_602)
);

BUFx8_ASAP7_75t_SL g603 ( 
.A(n_534),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_560),
.B(n_424),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_569),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_537),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_585),
.B(n_432),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_569),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_538),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_569),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_585),
.B(n_465),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_560),
.B(n_428),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_568),
.B(n_429),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_L g614 ( 
.A(n_524),
.B(n_481),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_540),
.B(n_453),
.Y(n_615)
);

INVxp33_ASAP7_75t_L g616 ( 
.A(n_588),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_569),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_L g618 ( 
.A(n_524),
.B(n_421),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_576),
.A2(n_402),
.B1(n_405),
.B2(n_469),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_537),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_576),
.B(n_436),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_578),
.B(n_438),
.Y(n_622)
);

AND2x6_ASAP7_75t_L g623 ( 
.A(n_557),
.B(n_359),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_569),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_533),
.B(n_439),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_533),
.B(n_500),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_539),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_533),
.B(n_500),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_539),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_541),
.A2(n_435),
.B1(n_504),
.B2(n_503),
.Y(n_630)
);

BUFx10_ASAP7_75t_L g631 ( 
.A(n_533),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_578),
.B(n_440),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_569),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_570),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_569),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_510),
.A2(n_422),
.B1(n_435),
.B2(n_326),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_534),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_569),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_538),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_574),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_574),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_574),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_541),
.A2(n_504),
.B1(n_505),
.B2(n_503),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_588),
.B(n_416),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_539),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_540),
.B(n_505),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_520),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_588),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_520),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_557),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_510),
.B(n_443),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_533),
.B(n_458),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_557),
.B(n_445),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_594),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_557),
.B(n_449),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_574),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_516),
.A2(n_310),
.B1(n_314),
.B2(n_306),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_538),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_519),
.B(n_506),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_520),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_517),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_574),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_520),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_573),
.B(n_417),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_545),
.B(n_506),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_545),
.B(n_455),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_574),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_SL g668 ( 
.A(n_538),
.B(n_459),
.Y(n_668)
);

OAI22xp33_ASAP7_75t_L g669 ( 
.A1(n_554),
.A2(n_462),
.B1(n_478),
.B2(n_461),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_513),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_574),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_516),
.B(n_485),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_550),
.B(n_487),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_513),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_541),
.A2(n_564),
.B1(n_573),
.B2(n_519),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_550),
.B(n_327),
.C(n_392),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_513),
.Y(n_677)
);

INVxp67_ASAP7_75t_SL g678 ( 
.A(n_517),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_551),
.B(n_493),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_574),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_SL g681 ( 
.A(n_590),
.B(n_471),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_573),
.B(n_475),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_540),
.B(n_489),
.Y(n_683)
);

BUFx10_ASAP7_75t_L g684 ( 
.A(n_519),
.Y(n_684)
);

NAND3xp33_ASAP7_75t_L g685 ( 
.A(n_551),
.B(n_392),
.C(n_368),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_590),
.Y(n_686)
);

OR2x6_ASAP7_75t_L g687 ( 
.A(n_542),
.B(n_543),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_553),
.B(n_508),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_553),
.B(n_556),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_587),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_587),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_517),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_512),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_520),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_520),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_556),
.B(n_483),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_542),
.B(n_496),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_542),
.B(n_232),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_587),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_573),
.Y(n_700)
);

BUFx8_ASAP7_75t_SL g701 ( 
.A(n_573),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_554),
.B(n_213),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_559),
.B(n_494),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_559),
.B(n_507),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_520),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_566),
.B(n_502),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_587),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_587),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_512),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_566),
.B(n_331),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_520),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_587),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_517),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_555),
.B(n_213),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_567),
.B(n_403),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_567),
.B(n_392),
.C(n_368),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_512),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_512),
.Y(n_718)
);

INVxp33_ASAP7_75t_L g719 ( 
.A(n_543),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_587),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_571),
.B(n_473),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_512),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_552),
.A2(n_319),
.B1(n_320),
.B2(n_317),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_571),
.B(n_480),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_581),
.A2(n_330),
.B1(n_332),
.B2(n_322),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_587),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_541),
.A2(n_338),
.B1(n_364),
.B2(n_288),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_581),
.B(n_363),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_517),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_546),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_526),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_583),
.B(n_418),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_526),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_526),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_586),
.B(n_369),
.Y(n_735)
);

BUFx8_ASAP7_75t_SL g736 ( 
.A(n_594),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_526),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_552),
.B(n_232),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_526),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_564),
.A2(n_364),
.B1(n_284),
.B2(n_278),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_546),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_546),
.Y(n_742)
);

NAND2xp33_ASAP7_75t_SL g743 ( 
.A(n_538),
.B(n_334),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_526),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_SL g745 ( 
.A(n_549),
.B(n_586),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_673),
.B(n_688),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_607),
.B(n_591),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_L g748 ( 
.A(n_660),
.B(n_526),
.Y(n_748)
);

A2O1A1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_619),
.A2(n_548),
.B(n_547),
.C(n_555),
.Y(n_749)
);

INVx8_ASAP7_75t_L g750 ( 
.A(n_623),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_637),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_696),
.Y(n_752)
);

INVxp33_ASAP7_75t_L g753 ( 
.A(n_648),
.Y(n_753)
);

NOR2xp67_ASAP7_75t_L g754 ( 
.A(n_650),
.B(n_562),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_740),
.A2(n_727),
.B1(n_630),
.B2(n_687),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_631),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_601),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_611),
.B(n_591),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_689),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_646),
.B(n_593),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_600),
.B(n_514),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_621),
.B(n_419),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_693),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_687),
.A2(n_564),
.B1(n_593),
.B2(n_579),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_600),
.B(n_514),
.Y(n_765)
);

NAND2xp33_ASAP7_75t_SL g766 ( 
.A(n_602),
.B(n_549),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_599),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_709),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_622),
.B(n_420),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_717),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_646),
.B(n_562),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_632),
.B(n_426),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_717),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_631),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_600),
.B(n_515),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_631),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_661),
.B(n_515),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_718),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_687),
.A2(n_564),
.B1(n_579),
.B2(n_575),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_661),
.B(n_523),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_661),
.B(n_523),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_634),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_619),
.A2(n_561),
.B1(n_563),
.B2(n_558),
.Y(n_783)
);

NOR2xp67_ASAP7_75t_SL g784 ( 
.A(n_599),
.B(n_549),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_614),
.B(n_562),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_601),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_634),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_698),
.B(n_565),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_698),
.B(n_565),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_738),
.B(n_565),
.Y(n_790)
);

NAND2x1_ASAP7_75t_L g791 ( 
.A(n_609),
.B(n_549),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_692),
.B(n_525),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_651),
.A2(n_589),
.B1(n_592),
.B2(n_584),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_721),
.B(n_427),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_659),
.A2(n_687),
.B1(n_672),
.B2(n_679),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_601),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_738),
.B(n_584),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_718),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_687),
.B(n_575),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_692),
.B(n_525),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_598),
.B(n_575),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_606),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_722),
.Y(n_803)
);

OR2x6_ASAP7_75t_L g804 ( 
.A(n_659),
.B(n_579),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_703),
.B(n_451),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_666),
.B(n_584),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_678),
.A2(n_532),
.B(n_531),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_692),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_710),
.B(n_589),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_615),
.B(n_589),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_615),
.B(n_592),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_722),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_713),
.B(n_531),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_SL g814 ( 
.A(n_681),
.B(n_518),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_702),
.B(n_592),
.Y(n_815)
);

AO21x2_ASAP7_75t_L g816 ( 
.A1(n_730),
.A2(n_561),
.B(n_558),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_702),
.B(n_596),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_714),
.B(n_652),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_626),
.A2(n_532),
.B(n_548),
.C(n_547),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_714),
.B(n_596),
.Y(n_820)
);

NOR2x1p5_ASAP7_75t_L g821 ( 
.A(n_598),
.B(n_563),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_730),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_R g823 ( 
.A(n_668),
.B(n_457),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_704),
.B(n_518),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_606),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_SL g826 ( 
.A(n_732),
.B(n_549),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_731),
.A2(n_528),
.B(n_526),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_631),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_659),
.A2(n_580),
.B1(n_582),
.B2(n_577),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_606),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_645),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_652),
.B(n_597),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_713),
.B(n_528),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_706),
.B(n_577),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_652),
.B(n_597),
.Y(n_835)
);

OR2x6_ASAP7_75t_L g836 ( 
.A(n_659),
.B(n_580),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_628),
.B(n_597),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_713),
.B(n_528),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_719),
.B(n_613),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_683),
.B(n_547),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_683),
.B(n_547),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_697),
.B(n_548),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_741),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_697),
.B(n_682),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_645),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_682),
.B(n_659),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_618),
.B(n_548),
.C(n_341),
.Y(n_847)
);

OAI21xp5_ASAP7_75t_L g848 ( 
.A1(n_647),
.A2(n_564),
.B(n_511),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_682),
.B(n_528),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_682),
.B(n_528),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_665),
.B(n_528),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_741),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_636),
.A2(n_388),
.B1(n_372),
.B2(n_375),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_643),
.B(n_259),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_644),
.B(n_259),
.Y(n_855)
);

INVx8_ASAP7_75t_L g856 ( 
.A(n_623),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_742),
.Y(n_857)
);

NOR3xp33_ASAP7_75t_L g858 ( 
.A(n_669),
.B(n_264),
.C(n_261),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_729),
.B(n_684),
.Y(n_859)
);

AND2x2_ASAP7_75t_SL g860 ( 
.A(n_675),
.B(n_216),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_700),
.B(n_528),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_729),
.B(n_742),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_729),
.B(n_528),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_684),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_645),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_670),
.Y(n_866)
);

OAI221xp5_ASAP7_75t_L g867 ( 
.A1(n_723),
.A2(n_264),
.B1(n_328),
.B2(n_315),
.C(n_340),
.Y(n_867)
);

NAND2x1p5_ASAP7_75t_L g868 ( 
.A(n_599),
.B(n_653),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_644),
.B(n_261),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_670),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_620),
.B(n_529),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_674),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_620),
.B(n_529),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_684),
.B(n_529),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_627),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_627),
.B(n_529),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_629),
.B(n_529),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_674),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_629),
.B(n_529),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_684),
.B(n_728),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_677),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_735),
.B(n_623),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_664),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_715),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_677),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_605),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_660),
.B(n_529),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_604),
.A2(n_388),
.B1(n_372),
.B2(n_375),
.Y(n_888)
);

INVxp33_ASAP7_75t_L g889 ( 
.A(n_616),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_L g890 ( 
.A(n_660),
.B(n_529),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_724),
.B(n_625),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_623),
.B(n_530),
.Y(n_892)
);

OR2x2_ASAP7_75t_L g893 ( 
.A(n_664),
.B(n_278),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_SL g894 ( 
.A1(n_686),
.A2(n_313),
.B1(n_241),
.B2(n_232),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_623),
.B(n_530),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_701),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_612),
.A2(n_385),
.B1(n_390),
.B2(n_397),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_723),
.B(n_284),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_660),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_623),
.B(n_530),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_660),
.B(n_530),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_623),
.B(n_720),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_737),
.B(n_530),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_655),
.B(n_342),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_731),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_605),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_746),
.B(n_609),
.Y(n_907)
);

OR2x2_ASAP7_75t_L g908 ( 
.A(n_787),
.B(n_751),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_771),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_782),
.Y(n_910)
);

AOI21xp33_ASAP7_75t_L g911 ( 
.A1(n_772),
.A2(n_654),
.B(n_657),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_884),
.A2(n_752),
.B(n_749),
.C(n_747),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_761),
.A2(n_744),
.B(n_733),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_756),
.B(n_609),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_834),
.B(n_737),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_761),
.A2(n_649),
.B(n_647),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_758),
.B(n_737),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_875),
.Y(n_918)
);

CKINVDCx10_ASAP7_75t_R g919 ( 
.A(n_804),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_765),
.A2(n_744),
.B(n_733),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_811),
.B(n_737),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_818),
.A2(n_639),
.B1(n_658),
.B2(n_609),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_811),
.B(n_725),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_765),
.A2(n_775),
.B(n_903),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_775),
.A2(n_649),
.B(n_647),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_848),
.A2(n_663),
.B(n_649),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_795),
.A2(n_658),
.B1(n_639),
.B2(n_633),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_863),
.A2(n_658),
.B(n_639),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_807),
.A2(n_694),
.B(n_663),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_851),
.A2(n_658),
.B(n_639),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_762),
.B(n_603),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_899),
.A2(n_745),
.B(n_694),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_839),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_759),
.B(n_610),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_783),
.B(n_610),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_844),
.B(n_610),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_822),
.Y(n_937)
);

OAI321xp33_ASAP7_75t_L g938 ( 
.A1(n_867),
.A2(n_315),
.A3(n_318),
.B1(n_293),
.B2(n_340),
.C(n_299),
.Y(n_938)
);

INVx1_ASAP7_75t_SL g939 ( 
.A(n_889),
.Y(n_939)
);

BUFx2_ASAP7_75t_SL g940 ( 
.A(n_896),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_755),
.A2(n_635),
.B1(n_667),
.B2(n_633),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_827),
.A2(n_694),
.B(n_663),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_799),
.B(n_602),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_862),
.A2(n_705),
.B(n_695),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_880),
.A2(n_705),
.B(n_695),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_788),
.B(n_789),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_790),
.B(n_633),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_774),
.B(n_743),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_887),
.A2(n_705),
.B(n_695),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_767),
.Y(n_950)
);

AOI21xp33_ASAP7_75t_L g951 ( 
.A1(n_753),
.A2(n_676),
.B(n_617),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_829),
.A2(n_841),
.B(n_842),
.C(n_840),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_887),
.A2(n_901),
.B(n_806),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_797),
.B(n_633),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_777),
.A2(n_739),
.B(n_711),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_901),
.A2(n_739),
.B(n_711),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_776),
.A2(n_667),
.B1(n_708),
.B2(n_635),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_776),
.A2(n_667),
.B1(n_708),
.B2(n_635),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_871),
.A2(n_739),
.B(n_711),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_858),
.A2(n_667),
.B(n_708),
.C(n_726),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_777),
.A2(n_624),
.B(n_608),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_873),
.A2(n_640),
.B(n_638),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_785),
.A2(n_640),
.B(n_638),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_760),
.A2(n_318),
.B(n_328),
.C(n_305),
.Y(n_964)
);

INVx11_ASAP7_75t_L g965 ( 
.A(n_896),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_780),
.A2(n_792),
.B(n_781),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_767),
.Y(n_967)
);

INVx6_ASAP7_75t_L g968 ( 
.A(n_804),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_810),
.B(n_821),
.Y(n_969)
);

AOI21x1_ASAP7_75t_L g970 ( 
.A1(n_892),
.A2(n_642),
.B(n_641),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_799),
.B(n_804),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_875),
.Y(n_972)
);

NOR2x1p5_ASAP7_75t_L g973 ( 
.A(n_855),
.B(n_736),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_875),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_843),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_815),
.B(n_708),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_817),
.B(n_726),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_820),
.B(n_726),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_805),
.B(n_660),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_832),
.B(n_734),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_804),
.Y(n_981)
);

AOI21xp33_ASAP7_75t_L g982 ( 
.A1(n_753),
.A2(n_860),
.B(n_794),
.Y(n_982)
);

BUFx8_ASAP7_75t_L g983 ( 
.A(n_883),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_835),
.B(n_734),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_801),
.B(n_883),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_823),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_860),
.A2(n_676),
.B1(n_313),
.B2(n_241),
.Y(n_987)
);

AND2x2_ASAP7_75t_SL g988 ( 
.A(n_814),
.B(n_305),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_R g989 ( 
.A(n_766),
.B(n_641),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_779),
.B(n_734),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_809),
.B(n_854),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_854),
.B(n_734),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_891),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_869),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_846),
.B(n_734),
.Y(n_995)
);

OAI22xp33_ASAP7_75t_L g996 ( 
.A1(n_898),
.A2(n_386),
.B1(n_357),
.B2(n_361),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_823),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_836),
.A2(n_691),
.B1(n_642),
.B2(n_712),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_852),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_764),
.B(n_734),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_833),
.A2(n_662),
.B(n_656),
.Y(n_1001)
);

BUFx2_ASAP7_75t_SL g1002 ( 
.A(n_754),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_828),
.B(n_656),
.Y(n_1003)
);

AO21x1_ASAP7_75t_L g1004 ( 
.A1(n_882),
.A2(n_680),
.B(n_671),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_833),
.A2(n_680),
.B(n_671),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_838),
.A2(n_691),
.B(n_690),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_838),
.A2(n_699),
.B(n_690),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_780),
.A2(n_707),
.B(n_699),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_853),
.A2(n_716),
.B(n_685),
.C(n_398),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_889),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_748),
.A2(n_535),
.B(n_530),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_824),
.B(n_904),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_781),
.A2(n_800),
.B(n_813),
.C(n_792),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_893),
.B(n_343),
.Y(n_1014)
);

OAI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_836),
.A2(n_378),
.B1(n_344),
.B2(n_351),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_748),
.A2(n_535),
.B(n_530),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_849),
.B(n_850),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_800),
.A2(n_716),
.B(n_685),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_826),
.B(n_509),
.Y(n_1019)
);

CKINVDCx8_ASAP7_75t_R g1020 ( 
.A(n_836),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_836),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_813),
.A2(n_511),
.B(n_509),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_890),
.A2(n_874),
.B(n_876),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_857),
.Y(n_1024)
);

AOI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_861),
.A2(n_376),
.B(n_373),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_808),
.B(n_530),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_828),
.B(n_535),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_763),
.Y(n_1028)
);

OR2x6_ASAP7_75t_L g1029 ( 
.A(n_750),
.B(n_269),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_750),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_877),
.A2(n_544),
.B(n_535),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_750),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_864),
.B(n_535),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_837),
.B(n_535),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_888),
.B(n_535),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_819),
.A2(n_398),
.B(n_400),
.C(n_366),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_750),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_856),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_SL g1039 ( 
.A(n_868),
.B(n_381),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_897),
.B(n_535),
.Y(n_1040)
);

AO21x1_ASAP7_75t_L g1041 ( 
.A1(n_895),
.A2(n_224),
.B(n_216),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_879),
.A2(n_544),
.B(n_235),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_894),
.B(n_395),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_816),
.B(n_544),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_900),
.A2(n_522),
.B(n_521),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_890),
.A2(n_770),
.B(n_768),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_886),
.A2(n_572),
.B(n_235),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_816),
.B(n_544),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_856),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_906),
.A2(n_572),
.B(n_258),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_773),
.A2(n_544),
.B(n_258),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_778),
.A2(n_544),
.B(n_337),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_859),
.B(n_353),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_798),
.A2(n_812),
.B(n_803),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_757),
.B(n_544),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_874),
.A2(n_544),
.B(n_337),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_905),
.A2(n_389),
.B(n_224),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_866),
.Y(n_1058)
);

OR2x6_ASAP7_75t_L g1059 ( 
.A(n_856),
.B(n_868),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_847),
.B(n_211),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_870),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_872),
.B(n_878),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_881),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_757),
.B(n_521),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_881),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_786),
.B(n_521),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_786),
.B(n_522),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_796),
.A2(n_536),
.B(n_527),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_885),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_905),
.A2(n_389),
.B(n_536),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_793),
.A2(n_294),
.B1(n_291),
.B2(n_286),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_796),
.B(n_527),
.Y(n_1072)
);

BUFx4f_ASAP7_75t_L g1073 ( 
.A(n_856),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_902),
.B(n_212),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_802),
.B(n_221),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_802),
.B(n_4),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_825),
.A2(n_279),
.B(n_399),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_825),
.B(n_226),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_830),
.B(n_231),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_831),
.A2(n_277),
.B(n_396),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_831),
.B(n_572),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_845),
.A2(n_274),
.B(n_393),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_937),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1012),
.B(n_845),
.Y(n_1084)
);

INVx4_ASAP7_75t_L g1085 ( 
.A(n_965),
.Y(n_1085)
);

BUFx4f_ASAP7_75t_SL g1086 ( 
.A(n_983),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_912),
.A2(n_865),
.B(n_885),
.C(n_791),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_SL g1088 ( 
.A1(n_988),
.A2(n_280),
.B1(n_384),
.B2(n_382),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_993),
.B(n_865),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_933),
.B(n_784),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_908),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_915),
.A2(n_247),
.B(n_380),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1045),
.A2(n_214),
.B(n_572),
.Y(n_1093)
);

BUFx12f_ASAP7_75t_L g1094 ( 
.A(n_997),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1063),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_983),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_1014),
.A2(n_12),
.B(n_15),
.C(n_16),
.Y(n_1097)
);

O2A1O1Ixp5_ASAP7_75t_SL g1098 ( 
.A1(n_911),
.A2(n_982),
.B(n_1075),
.C(n_1025),
.Y(n_1098)
);

AOI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1041),
.A2(n_214),
.B(n_572),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_946),
.A2(n_244),
.B(n_379),
.Y(n_1100)
);

INVx5_ASAP7_75t_L g1101 ( 
.A(n_1059),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1065),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_910),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_969),
.B(n_16),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_909),
.A2(n_246),
.B1(n_239),
.B2(n_238),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1069),
.Y(n_1106)
);

O2A1O1Ixp5_ASAP7_75t_L g1107 ( 
.A1(n_948),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_1107)
);

O2A1O1Ixp5_ASAP7_75t_L g1108 ( 
.A1(n_907),
.A2(n_23),
.B(n_27),
.C(n_29),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1028),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_923),
.A2(n_237),
.B1(n_236),
.B2(n_248),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_994),
.B(n_27),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_985),
.B(n_30),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1017),
.A2(n_249),
.B1(n_377),
.B2(n_263),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_975),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_999),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_1073),
.B(n_265),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1024),
.Y(n_1117)
);

NAND3xp33_ASAP7_75t_L g1118 ( 
.A(n_931),
.B(n_312),
.C(n_270),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1010),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_971),
.B(n_32),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_930),
.A2(n_325),
.B(n_371),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_1030),
.Y(n_1122)
);

OAI22x1_ASAP7_75t_L g1123 ( 
.A1(n_973),
.A2(n_1043),
.B1(n_971),
.B2(n_981),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_939),
.B(n_35),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_919),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_981),
.B(n_35),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1034),
.A2(n_345),
.B(n_370),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_986),
.B(n_37),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1030),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_968),
.B(n_37),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_SL g1131 ( 
.A1(n_1020),
.A2(n_367),
.B1(n_350),
.B2(n_324),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_952),
.A2(n_302),
.B(n_298),
.C(n_285),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_922),
.A2(n_257),
.B(n_163),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_935),
.A2(n_257),
.B1(n_39),
.B2(n_42),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_917),
.A2(n_979),
.B1(n_998),
.B2(n_921),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_927),
.A2(n_928),
.B(n_1026),
.Y(n_1136)
);

OAI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_938),
.A2(n_257),
.B1(n_39),
.B2(n_43),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_SL g1138 ( 
.A(n_940),
.B(n_572),
.Y(n_1138)
);

O2A1O1Ixp5_ASAP7_75t_L g1139 ( 
.A1(n_1004),
.A2(n_38),
.B(n_43),
.C(n_44),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1015),
.B(n_214),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_966),
.B(n_1013),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_945),
.A2(n_257),
.B(n_171),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_995),
.B(n_989),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_987),
.A2(n_572),
.B1(n_257),
.B2(n_214),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1058),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1061),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_945),
.A2(n_159),
.B(n_102),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_992),
.Y(n_1148)
);

AOI21x1_ASAP7_75t_L g1149 ( 
.A1(n_970),
.A2(n_214),
.B(n_572),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_943),
.B(n_47),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_L g1151 ( 
.A1(n_1074),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1076),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_R g1153 ( 
.A(n_1073),
.B(n_205),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_953),
.A2(n_572),
.B(n_56),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_968),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_968),
.B(n_55),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1032),
.Y(n_1157)
);

CKINVDCx16_ASAP7_75t_R g1158 ( 
.A(n_1039),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_996),
.B(n_55),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1062),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_950),
.B(n_214),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_990),
.B(n_214),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_936),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_R g1164 ( 
.A(n_1032),
.B(n_200),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1021),
.B(n_62),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1059),
.B(n_62),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_964),
.A2(n_214),
.B(n_68),
.C(n_69),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_953),
.A2(n_67),
.B(n_68),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_950),
.B(n_67),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_962),
.A2(n_87),
.B(n_188),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_950),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_918),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1032),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_934),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_960),
.B(n_980),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_972),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_974),
.B(n_74),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_962),
.A2(n_111),
.B(n_178),
.Y(n_1178)
);

O2A1O1Ixp5_ASAP7_75t_L g1179 ( 
.A1(n_1036),
.A2(n_74),
.B(n_75),
.C(n_76),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1064),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_967),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1002),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1066),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1067),
.Y(n_1184)
);

NOR2x1_ASAP7_75t_L g1185 ( 
.A(n_967),
.B(n_199),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_967),
.B(n_78),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_976),
.A2(n_978),
.B1(n_977),
.B2(n_984),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_957),
.B(n_80),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1053),
.B(n_82),
.Y(n_1189)
);

CKINVDCx8_ASAP7_75t_R g1190 ( 
.A(n_1053),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1038),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1000),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1060),
.A2(n_83),
.B(n_85),
.C(n_112),
.Y(n_1193)
);

OAI21xp33_ASAP7_75t_L g1194 ( 
.A1(n_1071),
.A2(n_126),
.B(n_127),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_947),
.B(n_144),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_954),
.B(n_174),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_958),
.B(n_176),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_929),
.A2(n_924),
.B(n_926),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1059),
.Y(n_1199)
);

NAND2x1p5_ASAP7_75t_L g1200 ( 
.A(n_1038),
.B(n_1049),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_951),
.B(n_1079),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1078),
.B(n_1003),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1054),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_941),
.B(n_1033),
.Y(n_1204)
);

NOR3xp33_ASAP7_75t_L g1205 ( 
.A(n_1082),
.B(n_1077),
.C(n_1080),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1029),
.B(n_1048),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1029),
.A2(n_1054),
.B1(n_1044),
.B2(n_1081),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1038),
.Y(n_1208)
);

CKINVDCx16_ASAP7_75t_R g1209 ( 
.A(n_1029),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_1081),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1072),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1049),
.B(n_1037),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_SL g1213 ( 
.A1(n_1049),
.A2(n_1047),
.B1(n_1050),
.B2(n_1018),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_924),
.B(n_1027),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1055),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_959),
.A2(n_1023),
.B(n_963),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1046),
.A2(n_1056),
.B(n_1008),
.C(n_961),
.Y(n_1217)
);

AOI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1051),
.A2(n_1052),
.B(n_1057),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1046),
.A2(n_1019),
.B1(n_914),
.B2(n_955),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1022),
.B(n_959),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_944),
.B(n_1031),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1057),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1035),
.B(n_1040),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_932),
.A2(n_913),
.B(n_920),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1056),
.A2(n_1009),
.B(n_913),
.C(n_920),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_916),
.A2(n_925),
.B(n_942),
.C(n_1006),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1070),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1037),
.B(n_1016),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1001),
.B(n_1005),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1068),
.Y(n_1230)
);

NOR3xp33_ASAP7_75t_SL g1231 ( 
.A(n_1007),
.B(n_949),
.C(n_956),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1042),
.A2(n_1051),
.B1(n_1052),
.B2(n_949),
.Y(n_1232)
);

CKINVDCx11_ASAP7_75t_R g1233 ( 
.A(n_1094),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1160),
.B(n_956),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1091),
.B(n_1011),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1187),
.A2(n_1225),
.A3(n_1198),
.B(n_1221),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1093),
.A2(n_1224),
.B(n_1216),
.Y(n_1237)
);

AOI221x1_ASAP7_75t_L g1238 ( 
.A1(n_1168),
.A2(n_1194),
.B1(n_1134),
.B2(n_1205),
.C(n_1193),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1083),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_SL g1240 ( 
.A1(n_1084),
.A2(n_1135),
.B(n_1201),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1137),
.A2(n_1088),
.B1(n_1158),
.B2(n_1104),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1218),
.A2(n_1136),
.B(n_1232),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1148),
.B(n_1201),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1104),
.A2(n_1204),
.B(n_1097),
.C(n_1202),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1103),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1232),
.A2(n_1142),
.B(n_1099),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1226),
.A2(n_1149),
.B(n_1227),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1141),
.A2(n_1214),
.B(n_1196),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1148),
.B(n_1204),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1171),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1141),
.A2(n_1214),
.B(n_1195),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1192),
.B(n_1152),
.Y(n_1252)
);

AOI221xp5_ASAP7_75t_L g1253 ( 
.A1(n_1137),
.A2(n_1111),
.B1(n_1124),
.B2(n_1167),
.C(n_1110),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1210),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1181),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1206),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1220),
.A2(n_1175),
.B(n_1197),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1188),
.A2(n_1132),
.B(n_1150),
.C(n_1174),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1203),
.A2(n_1217),
.A3(n_1219),
.B(n_1229),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1119),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1119),
.B(n_1146),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1130),
.A2(n_1156),
.B1(n_1120),
.B2(n_1166),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1120),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1190),
.B(n_1128),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1162),
.A2(n_1228),
.B(n_1229),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1188),
.A2(n_1166),
.B1(n_1154),
.B2(n_1114),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1115),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1175),
.A2(n_1197),
.B(n_1133),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_SL g1269 ( 
.A1(n_1209),
.A2(n_1086),
.B1(n_1124),
.B2(n_1125),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1089),
.B(n_1112),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1130),
.A2(n_1156),
.B1(n_1126),
.B2(n_1131),
.Y(n_1271)
);

NAND3xp33_ASAP7_75t_SL g1272 ( 
.A(n_1090),
.B(n_1118),
.C(n_1182),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1192),
.B(n_1180),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1095),
.A2(n_1102),
.B1(n_1106),
.B2(n_1189),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1147),
.A2(n_1170),
.B(n_1178),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1098),
.A2(n_1207),
.B(n_1215),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1129),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1117),
.B(n_1155),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1085),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1183),
.B(n_1184),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1129),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1087),
.A2(n_1143),
.B(n_1213),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1207),
.A2(n_1143),
.B(n_1161),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1126),
.A2(n_1105),
.B1(n_1123),
.B2(n_1177),
.Y(n_1284)
);

AOI221x1_ASAP7_75t_L g1285 ( 
.A1(n_1223),
.A2(n_1177),
.B1(n_1165),
.B2(n_1169),
.C(n_1186),
.Y(n_1285)
);

INVxp67_ASAP7_75t_L g1286 ( 
.A(n_1096),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1127),
.A2(n_1100),
.B(n_1092),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1223),
.A2(n_1211),
.A3(n_1145),
.B(n_1172),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1179),
.A2(n_1139),
.B(n_1231),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1176),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1231),
.A2(n_1108),
.B(n_1151),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1140),
.A2(n_1107),
.B(n_1113),
.C(n_1121),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1086),
.B(n_1155),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1199),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1185),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1116),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1230),
.A2(n_1101),
.A3(n_1144),
.B(n_1164),
.Y(n_1297)
);

AOI221xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1230),
.A2(n_1191),
.B1(n_1208),
.B2(n_1129),
.C(n_1122),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_L g1299 ( 
.A(n_1138),
.B(n_1129),
.C(n_1208),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1230),
.A2(n_1212),
.B(n_1101),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1157),
.Y(n_1301)
);

A2O1A1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1157),
.A2(n_1173),
.B(n_1212),
.C(n_1101),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1230),
.Y(n_1303)
);

AOI221xp5_ASAP7_75t_L g1304 ( 
.A1(n_1116),
.A2(n_1153),
.B1(n_1164),
.B2(n_1191),
.C(n_1208),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1153),
.Y(n_1305)
);

AO32x2_ASAP7_75t_L g1306 ( 
.A1(n_1191),
.A2(n_1187),
.A3(n_1134),
.B1(n_1135),
.B2(n_1219),
.Y(n_1306)
);

BUFx2_ASAP7_75t_R g1307 ( 
.A(n_1200),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1200),
.A2(n_1191),
.B(n_1208),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1141),
.A2(n_1214),
.B(n_1204),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1216),
.A2(n_1198),
.B(n_1224),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1120),
.B(n_787),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1187),
.A2(n_1004),
.A3(n_1041),
.B(n_1044),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1094),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1086),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1093),
.A2(n_1224),
.B(n_1216),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1141),
.A2(n_1214),
.B(n_1204),
.Y(n_1319)
);

AO22x2_ASAP7_75t_L g1320 ( 
.A1(n_1206),
.A2(n_795),
.B1(n_654),
.B2(n_898),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1084),
.B(n_991),
.Y(n_1321)
);

BUFx10_ASAP7_75t_L g1322 ( 
.A(n_1125),
.Y(n_1322)
);

AOI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1218),
.A2(n_1136),
.B(n_1224),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1101),
.B(n_971),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1093),
.A2(n_1224),
.B(n_1216),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1093),
.A2(n_1224),
.B(n_1216),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1129),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1330)
);

BUFx24_ASAP7_75t_L g1331 ( 
.A(n_1120),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1159),
.A2(n_746),
.B(n_884),
.C(n_752),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1141),
.A2(n_1214),
.B(n_1204),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1083),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1093),
.A2(n_1224),
.B(n_1216),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1085),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1103),
.Y(n_1337)
);

AO32x2_ASAP7_75t_L g1338 ( 
.A1(n_1187),
.A2(n_1134),
.A3(n_1135),
.B1(n_1219),
.B2(n_1163),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1083),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1093),
.A2(n_1224),
.B(n_1216),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1083),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1084),
.B(n_991),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1103),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1084),
.B(n_991),
.Y(n_1347)
);

OAI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1158),
.A2(n_746),
.B1(n_619),
.B2(n_681),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1141),
.A2(n_1214),
.B(n_1204),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1084),
.B(n_991),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1091),
.B(n_908),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1083),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1103),
.B(n_884),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1083),
.Y(n_1355)
);

OR2x6_ASAP7_75t_L g1356 ( 
.A(n_1120),
.B(n_968),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1141),
.A2(n_1214),
.B(n_1204),
.Y(n_1357)
);

O2A1O1Ixp5_ASAP7_75t_SL g1358 ( 
.A1(n_1162),
.A2(n_1222),
.B(n_1168),
.C(n_1141),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1084),
.B(n_991),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1160),
.A2(n_746),
.B1(n_818),
.B2(n_783),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1159),
.A2(n_746),
.B(n_884),
.C(n_752),
.Y(n_1363)
);

INVxp67_ASAP7_75t_L g1364 ( 
.A(n_1091),
.Y(n_1364)
);

CKINVDCx6p67_ASAP7_75t_R g1365 ( 
.A(n_1094),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1162),
.A2(n_1205),
.B(n_1221),
.Y(n_1366)
);

BUFx10_ASAP7_75t_L g1367 ( 
.A(n_1125),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1160),
.B(n_762),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1158),
.B(n_1012),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1083),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1109),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1083),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1084),
.B(n_991),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1083),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_SL g1378 ( 
.A1(n_1097),
.A2(n_746),
.B(n_884),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1120),
.B(n_787),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1083),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1141),
.A2(n_1214),
.B(n_1204),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1083),
.Y(n_1382)
);

INVx4_ASAP7_75t_SL g1383 ( 
.A(n_1166),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1384)
);

INVx4_ASAP7_75t_L g1385 ( 
.A(n_1085),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1103),
.B(n_884),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1093),
.A2(n_1224),
.B(n_1216),
.Y(n_1387)
);

AO32x2_ASAP7_75t_L g1388 ( 
.A1(n_1187),
.A2(n_1134),
.A3(n_1135),
.B1(n_1219),
.B2(n_1163),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1129),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1187),
.A2(n_746),
.B(n_1136),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1093),
.A2(n_1224),
.B(n_1216),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1129),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1083),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1162),
.A2(n_1205),
.B(n_1221),
.Y(n_1394)
);

OAI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1262),
.A2(n_1271),
.B1(n_1348),
.B2(n_1266),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1233),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1383),
.B(n_1324),
.Y(n_1397)
);

BUFx12f_ASAP7_75t_L g1398 ( 
.A(n_1322),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1365),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1253),
.A2(n_1320),
.B1(n_1266),
.B2(n_1243),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1378),
.A2(n_1357),
.B1(n_1309),
.B2(n_1319),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1337),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_1351),
.Y(n_1403)
);

OAI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1356),
.A2(n_1284),
.B1(n_1362),
.B2(n_1333),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1315),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1320),
.A2(n_1243),
.B1(n_1369),
.B2(n_1375),
.Y(n_1406)
);

CKINVDCx6p67_ASAP7_75t_R g1407 ( 
.A(n_1331),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1345),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1322),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1309),
.A2(n_1357),
.B1(n_1349),
.B2(n_1333),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1319),
.A2(n_1381),
.B1(n_1349),
.B2(n_1362),
.Y(n_1411)
);

INVx4_ASAP7_75t_L g1412 ( 
.A(n_1385),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1367),
.Y(n_1413)
);

INVx6_ASAP7_75t_L g1414 ( 
.A(n_1383),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1381),
.A2(n_1347),
.B1(n_1350),
.B2(n_1360),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1249),
.A2(n_1263),
.B1(n_1321),
.B2(n_1375),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1321),
.A2(n_1360),
.B1(n_1344),
.B2(n_1347),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1344),
.A2(n_1350),
.B1(n_1270),
.B2(n_1249),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1373),
.A2(n_1252),
.B1(n_1264),
.B2(n_1379),
.Y(n_1419)
);

BUFx12f_ASAP7_75t_L g1420 ( 
.A(n_1367),
.Y(n_1420)
);

BUFx12f_ASAP7_75t_L g1421 ( 
.A(n_1305),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1252),
.A2(n_1313),
.B1(n_1356),
.B2(n_1383),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1267),
.Y(n_1423)
);

OAI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1356),
.A2(n_1238),
.B1(n_1285),
.B2(n_1260),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1279),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1296),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1256),
.A2(n_1274),
.B1(n_1273),
.B2(n_1280),
.Y(n_1427)
);

CKINVDCx11_ASAP7_75t_R g1428 ( 
.A(n_1336),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1334),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1256),
.A2(n_1273),
.B1(n_1280),
.B2(n_1254),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1254),
.A2(n_1304),
.B1(n_1290),
.B2(n_1295),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1269),
.A2(n_1354),
.B1(n_1386),
.B2(n_1272),
.Y(n_1432)
);

OAI22xp33_ASAP7_75t_R g1433 ( 
.A1(n_1245),
.A2(n_1293),
.B1(n_1363),
.B2(n_1332),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1289),
.A2(n_1282),
.B1(n_1240),
.B2(n_1393),
.Y(n_1434)
);

CKINVDCx11_ASAP7_75t_R g1435 ( 
.A(n_1250),
.Y(n_1435)
);

BUFx2_ASAP7_75t_SL g1436 ( 
.A(n_1255),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1281),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_1364),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1286),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1340),
.A2(n_1374),
.B1(n_1342),
.B2(n_1382),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_SL g1441 ( 
.A1(n_1289),
.A2(n_1377),
.B1(n_1352),
.B2(n_1370),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1355),
.Y(n_1442)
);

BUFx2_ASAP7_75t_SL g1443 ( 
.A(n_1328),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1380),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1278),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1261),
.A2(n_1251),
.B1(n_1248),
.B2(n_1235),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1258),
.A2(n_1311),
.B1(n_1390),
.B2(n_1384),
.Y(n_1447)
);

BUFx8_ASAP7_75t_L g1448 ( 
.A(n_1328),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1294),
.Y(n_1449)
);

CKINVDCx6p67_ASAP7_75t_R g1450 ( 
.A(n_1389),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1276),
.A2(n_1291),
.B1(n_1343),
.B2(n_1376),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1234),
.A2(n_1299),
.B1(n_1291),
.B2(n_1268),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1288),
.B(n_1301),
.Y(n_1453)
);

INVx6_ASAP7_75t_L g1454 ( 
.A(n_1389),
.Y(n_1454)
);

INVx6_ASAP7_75t_L g1455 ( 
.A(n_1307),
.Y(n_1455)
);

CKINVDCx11_ASAP7_75t_R g1456 ( 
.A(n_1303),
.Y(n_1456)
);

BUFx4f_ASAP7_75t_SL g1457 ( 
.A(n_1277),
.Y(n_1457)
);

OAI22x1_ASAP7_75t_L g1458 ( 
.A1(n_1277),
.A2(n_1392),
.B1(n_1306),
.B2(n_1388),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1392),
.B(n_1316),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1308),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1283),
.A2(n_1257),
.B1(n_1366),
.B2(n_1394),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1366),
.A2(n_1394),
.B1(n_1372),
.B2(n_1371),
.Y(n_1462)
);

CKINVDCx20_ASAP7_75t_R g1463 ( 
.A(n_1300),
.Y(n_1463)
);

INVx6_ASAP7_75t_L g1464 ( 
.A(n_1298),
.Y(n_1464)
);

INVx5_ASAP7_75t_L g1465 ( 
.A(n_1298),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1310),
.A2(n_1359),
.B(n_1330),
.Y(n_1466)
);

OAI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1325),
.A2(n_1339),
.B1(n_1361),
.B2(n_1353),
.Y(n_1467)
);

INVx6_ASAP7_75t_L g1468 ( 
.A(n_1302),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1329),
.A2(n_1346),
.B1(n_1388),
.B2(n_1338),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1306),
.A2(n_1338),
.B1(n_1388),
.B2(n_1297),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1265),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1287),
.A2(n_1275),
.B1(n_1306),
.B2(n_1247),
.Y(n_1472)
);

BUFx8_ASAP7_75t_L g1473 ( 
.A(n_1338),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1292),
.A2(n_1312),
.B1(n_1323),
.B2(n_1358),
.Y(n_1474)
);

INVx6_ASAP7_75t_L g1475 ( 
.A(n_1236),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_SL g1476 ( 
.A1(n_1246),
.A2(n_1312),
.B1(n_1242),
.B2(n_1236),
.Y(n_1476)
);

INVxp67_ASAP7_75t_SL g1477 ( 
.A(n_1237),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1236),
.A2(n_1314),
.B1(n_1318),
.B2(n_1326),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1327),
.A2(n_1335),
.B1(n_1341),
.B2(n_1387),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1391),
.Y(n_1480)
);

BUFx8_ASAP7_75t_L g1481 ( 
.A(n_1337),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1239),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1262),
.A2(n_746),
.B1(n_619),
.B2(n_1271),
.Y(n_1483)
);

CKINVDCx11_ASAP7_75t_R g1484 ( 
.A(n_1317),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1241),
.A2(n_1348),
.B1(n_762),
.B2(n_769),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1239),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1351),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1241),
.A2(n_1348),
.B1(n_762),
.B2(n_769),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1244),
.A2(n_746),
.B1(n_1241),
.B2(n_884),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1313),
.B(n_1379),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1324),
.Y(n_1491)
);

INVx6_ASAP7_75t_L g1492 ( 
.A(n_1385),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1348),
.A2(n_762),
.B1(n_769),
.B2(n_681),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1348),
.A2(n_762),
.B1(n_769),
.B2(n_681),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1239),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1243),
.B(n_1368),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1241),
.A2(n_1348),
.B1(n_762),
.B2(n_769),
.Y(n_1497)
);

INVx6_ASAP7_75t_L g1498 ( 
.A(n_1385),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_1317),
.Y(n_1499)
);

BUFx4f_ASAP7_75t_L g1500 ( 
.A(n_1365),
.Y(n_1500)
);

OAI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1244),
.A2(n_746),
.B(n_884),
.Y(n_1501)
);

OAI21xp33_ASAP7_75t_L g1502 ( 
.A1(n_1244),
.A2(n_746),
.B(n_1378),
.Y(n_1502)
);

BUFx8_ASAP7_75t_L g1503 ( 
.A(n_1337),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1259),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1241),
.A2(n_1348),
.B1(n_762),
.B2(n_769),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1241),
.A2(n_1348),
.B1(n_762),
.B2(n_769),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1324),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1337),
.Y(n_1508)
);

CKINVDCx11_ASAP7_75t_R g1509 ( 
.A(n_1317),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1317),
.Y(n_1510)
);

INVxp67_ASAP7_75t_SL g1511 ( 
.A(n_1242),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1239),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1241),
.A2(n_1348),
.B1(n_762),
.B2(n_769),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1239),
.Y(n_1514)
);

CKINVDCx8_ASAP7_75t_R g1515 ( 
.A(n_1315),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1244),
.A2(n_746),
.B1(n_1241),
.B2(n_884),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1244),
.A2(n_746),
.B1(n_1241),
.B2(n_884),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1244),
.A2(n_746),
.B1(n_1241),
.B2(n_884),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1241),
.A2(n_746),
.B(n_931),
.Y(n_1519)
);

BUFx2_ASAP7_75t_SL g1520 ( 
.A(n_1317),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1239),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1348),
.A2(n_772),
.B1(n_762),
.B2(n_769),
.Y(n_1522)
);

OAI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1262),
.A2(n_746),
.B1(n_619),
.B2(n_1271),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1337),
.Y(n_1524)
);

CKINVDCx6p67_ASAP7_75t_R g1525 ( 
.A(n_1233),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1348),
.A2(n_762),
.B1(n_769),
.B2(n_681),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1262),
.A2(n_746),
.B1(n_619),
.B2(n_1271),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1348),
.A2(n_762),
.B1(n_769),
.B2(n_681),
.Y(n_1528)
);

INVx4_ASAP7_75t_L g1529 ( 
.A(n_1385),
.Y(n_1529)
);

INVx4_ASAP7_75t_L g1530 ( 
.A(n_1385),
.Y(n_1530)
);

INVx4_ASAP7_75t_L g1531 ( 
.A(n_1385),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1317),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_SL g1533 ( 
.A1(n_1320),
.A2(n_681),
.B1(n_769),
.B2(n_762),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1317),
.Y(n_1534)
);

INVx4_ASAP7_75t_L g1535 ( 
.A(n_1385),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1233),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1281),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1317),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1241),
.A2(n_1348),
.B1(n_762),
.B2(n_769),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1239),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1351),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1317),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1281),
.Y(n_1543)
);

AOI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1474),
.A2(n_1447),
.B(n_1480),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1470),
.B(n_1504),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1466),
.A2(n_1472),
.B(n_1479),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1453),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1465),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1470),
.B(n_1504),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1465),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1471),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_SL g1552 ( 
.A(n_1515),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1475),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1423),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1429),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1401),
.B(n_1411),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1442),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1445),
.Y(n_1558)
);

INVx4_ASAP7_75t_L g1559 ( 
.A(n_1464),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1444),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1482),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1486),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1495),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1512),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1514),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1496),
.B(n_1418),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1410),
.B(n_1411),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1521),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1458),
.Y(n_1569)
);

AO21x2_ASAP7_75t_L g1570 ( 
.A1(n_1469),
.A2(n_1467),
.B(n_1424),
.Y(n_1570)
);

INVx4_ASAP7_75t_SL g1571 ( 
.A(n_1464),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1540),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1459),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1508),
.Y(n_1574)
);

OAI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1462),
.A2(n_1461),
.B(n_1452),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1464),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1400),
.B(n_1410),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1475),
.B(n_1415),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1460),
.Y(n_1579)
);

CKINVDCx11_ASAP7_75t_R g1580 ( 
.A(n_1396),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1460),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1511),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1511),
.Y(n_1583)
);

AOI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1489),
.A2(n_1516),
.B(n_1518),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1524),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1469),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1473),
.Y(n_1587)
);

OR2x6_ASAP7_75t_L g1588 ( 
.A(n_1414),
.B(n_1468),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1468),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1418),
.B(n_1417),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1473),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1446),
.Y(n_1592)
);

AOI211x1_ASAP7_75t_L g1593 ( 
.A1(n_1483),
.A2(n_1527),
.B(n_1523),
.C(n_1517),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1446),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1477),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1463),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1397),
.B(n_1537),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1468),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1533),
.A2(n_1494),
.B1(n_1493),
.B2(n_1528),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1402),
.Y(n_1600)
);

OAI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1522),
.A2(n_1502),
.B(n_1501),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1403),
.B(n_1487),
.Y(n_1602)
);

AO21x2_ASAP7_75t_L g1603 ( 
.A1(n_1467),
.A2(n_1424),
.B(n_1395),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1533),
.A2(n_1526),
.B1(n_1485),
.B2(n_1488),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1448),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1448),
.Y(n_1606)
);

OA21x2_ASAP7_75t_L g1607 ( 
.A1(n_1477),
.A2(n_1406),
.B(n_1415),
.Y(n_1607)
);

CKINVDCx11_ASAP7_75t_R g1608 ( 
.A(n_1484),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1440),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1441),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1456),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1441),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1436),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1543),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1434),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1434),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1476),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1476),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1509),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1408),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1478),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1478),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1417),
.A2(n_1430),
.B(n_1427),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1537),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1416),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1416),
.B(n_1541),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1451),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1490),
.B(n_1419),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1451),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1404),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1454),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1481),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1404),
.A2(n_1527),
.B(n_1523),
.Y(n_1633)
);

INVx4_ASAP7_75t_L g1634 ( 
.A(n_1414),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1422),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1422),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1443),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1419),
.B(n_1426),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1483),
.B(n_1432),
.Y(n_1639)
);

AO21x2_ASAP7_75t_L g1640 ( 
.A1(n_1519),
.A2(n_1431),
.B(n_1539),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1450),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1499),
.B(n_1538),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1481),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1503),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1433),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1485),
.A2(n_1488),
.B(n_1539),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_SL g1647 ( 
.A(n_1536),
.B(n_1500),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1510),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1457),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1407),
.B(n_1437),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1435),
.B(n_1491),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1457),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1503),
.B(n_1505),
.Y(n_1653)
);

OA21x2_ASAP7_75t_L g1654 ( 
.A1(n_1497),
.A2(n_1505),
.B(n_1513),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1491),
.B(n_1507),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1578),
.B(n_1449),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1633),
.A2(n_1497),
.B(n_1506),
.Y(n_1657)
);

OA21x2_ASAP7_75t_L g1658 ( 
.A1(n_1546),
.A2(n_1513),
.B(n_1506),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1573),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1596),
.B(n_1520),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1558),
.B(n_1439),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1639),
.A2(n_1500),
.B(n_1438),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1596),
.B(n_1542),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_R g1664 ( 
.A(n_1580),
.B(n_1525),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1566),
.B(n_1425),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1596),
.B(n_1534),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1601),
.A2(n_1646),
.B(n_1604),
.C(n_1577),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1651),
.B(n_1428),
.Y(n_1668)
);

AOI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1645),
.A2(n_1413),
.B1(n_1409),
.B2(n_1399),
.C(n_1405),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1651),
.B(n_1455),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1600),
.B(n_1455),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_SL g1672 ( 
.A1(n_1603),
.A2(n_1535),
.B(n_1412),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1573),
.Y(n_1673)
);

A2O1A1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1646),
.A2(n_1532),
.B(n_1498),
.C(n_1492),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1554),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1603),
.A2(n_1529),
.B(n_1530),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1574),
.B(n_1421),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1567),
.B(n_1585),
.Y(n_1678)
);

AOI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1645),
.A2(n_1529),
.B1(n_1531),
.B2(n_1398),
.C(n_1420),
.Y(n_1679)
);

AOI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1610),
.A2(n_1612),
.B1(n_1590),
.B2(n_1593),
.C(n_1586),
.Y(n_1680)
);

OAI21x1_ASAP7_75t_SL g1681 ( 
.A1(n_1584),
.A2(n_1576),
.B(n_1556),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1611),
.B(n_1620),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1613),
.Y(n_1683)
);

AOI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1612),
.A2(n_1593),
.B1(n_1586),
.B2(n_1625),
.C(n_1621),
.Y(n_1684)
);

OA21x2_ASAP7_75t_L g1685 ( 
.A1(n_1546),
.A2(n_1575),
.B(n_1627),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1582),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1576),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1599),
.A2(n_1654),
.B1(n_1584),
.B2(n_1577),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1615),
.A2(n_1616),
.B(n_1654),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1611),
.B(n_1628),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1587),
.B(n_1591),
.Y(n_1691)
);

AO21x1_ASAP7_75t_L g1692 ( 
.A1(n_1627),
.A2(n_1629),
.B(n_1622),
.Y(n_1692)
);

AO22x2_ASAP7_75t_L g1693 ( 
.A1(n_1622),
.A2(n_1618),
.B1(n_1617),
.B2(n_1545),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1654),
.A2(n_1640),
.B1(n_1598),
.B2(n_1589),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1640),
.B(n_1653),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1571),
.B(n_1548),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1650),
.B(n_1655),
.Y(n_1697)
);

OA21x2_ASAP7_75t_L g1698 ( 
.A1(n_1575),
.A2(n_1629),
.B(n_1544),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1630),
.A2(n_1625),
.B(n_1618),
.C(n_1617),
.Y(n_1699)
);

A2O1A1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1630),
.A2(n_1594),
.B(n_1592),
.C(n_1545),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1555),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1582),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1650),
.B(n_1655),
.Y(n_1703)
);

AOI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1569),
.A2(n_1549),
.B1(n_1570),
.B2(n_1626),
.C(n_1609),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1597),
.B(n_1561),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1549),
.A2(n_1598),
.B(n_1589),
.C(n_1638),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1597),
.B(n_1563),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1597),
.B(n_1565),
.Y(n_1708)
);

AO32x2_ASAP7_75t_L g1709 ( 
.A1(n_1559),
.A2(n_1634),
.A3(n_1606),
.B1(n_1605),
.B2(n_1638),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1583),
.Y(n_1710)
);

O2A1O1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1643),
.A2(n_1644),
.B(n_1649),
.C(n_1652),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1572),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_SL g1713 ( 
.A1(n_1623),
.A2(n_1589),
.B1(n_1598),
.B2(n_1607),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1631),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1649),
.A2(n_1652),
.B1(n_1632),
.B2(n_1641),
.Y(n_1715)
);

OA21x2_ASAP7_75t_L g1716 ( 
.A1(n_1544),
.A2(n_1583),
.B(n_1595),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1637),
.B(n_1641),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1623),
.A2(n_1609),
.B1(n_1635),
.B2(n_1636),
.Y(n_1718)
);

INVx5_ASAP7_75t_L g1719 ( 
.A(n_1550),
.Y(n_1719)
);

AOI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1547),
.A2(n_1635),
.B1(n_1568),
.B2(n_1560),
.C(n_1557),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1579),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1705),
.B(n_1595),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1659),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1678),
.B(n_1607),
.Y(n_1724)
);

NOR2x1_ASAP7_75t_L g1725 ( 
.A(n_1672),
.B(n_1614),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1707),
.B(n_1607),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1657),
.A2(n_1623),
.B1(n_1607),
.B2(n_1588),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1659),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1673),
.Y(n_1729)
);

INVx4_ASAP7_75t_L g1730 ( 
.A(n_1719),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1686),
.B(n_1564),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1686),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1695),
.B(n_1547),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1702),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1708),
.B(n_1581),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1702),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1710),
.Y(n_1737)
);

INVx3_ASAP7_75t_L g1738 ( 
.A(n_1721),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1690),
.B(n_1581),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1710),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1675),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1695),
.B(n_1562),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1719),
.B(n_1579),
.Y(n_1743)
);

INVx2_ASAP7_75t_SL g1744 ( 
.A(n_1719),
.Y(n_1744)
);

INVxp67_ASAP7_75t_SL g1745 ( 
.A(n_1716),
.Y(n_1745)
);

INVx2_ASAP7_75t_R g1746 ( 
.A(n_1701),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1665),
.B(n_1608),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1704),
.A2(n_1623),
.B1(n_1588),
.B2(n_1553),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1668),
.B(n_1552),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1691),
.B(n_1579),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1716),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_SL g1752 ( 
.A1(n_1667),
.A2(n_1637),
.B1(n_1642),
.B2(n_1551),
.C(n_1624),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1693),
.A2(n_1692),
.B1(n_1688),
.B2(n_1680),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1712),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1697),
.B(n_1579),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1703),
.B(n_1551),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1681),
.Y(n_1757)
);

INVxp67_ASAP7_75t_SL g1758 ( 
.A(n_1716),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1660),
.B(n_1619),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1687),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1685),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1714),
.Y(n_1762)
);

INVxp67_ASAP7_75t_SL g1763 ( 
.A(n_1698),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1685),
.Y(n_1764)
);

OAI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1727),
.A2(n_1658),
.B1(n_1694),
.B2(n_1689),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1732),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1726),
.B(n_1713),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1723),
.B(n_1667),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1764),
.Y(n_1769)
);

INVx4_ASAP7_75t_SL g1770 ( 
.A(n_1743),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1730),
.B(n_1696),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1732),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1734),
.Y(n_1773)
);

OAI31xp33_ASAP7_75t_L g1774 ( 
.A1(n_1753),
.A2(n_1700),
.A3(n_1699),
.B(n_1693),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1734),
.Y(n_1775)
);

AO21x2_ASAP7_75t_L g1776 ( 
.A1(n_1745),
.A2(n_1699),
.B(n_1700),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1736),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1761),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1736),
.Y(n_1779)
);

BUFx3_ASAP7_75t_L g1780 ( 
.A(n_1744),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1757),
.B(n_1711),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1757),
.B(n_1715),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1737),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1761),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1737),
.Y(n_1785)
);

OAI321xp33_ASAP7_75t_L g1786 ( 
.A1(n_1727),
.A2(n_1684),
.A3(n_1718),
.B1(n_1674),
.B2(n_1662),
.C(n_1706),
.Y(n_1786)
);

AOI33xp33_ASAP7_75t_L g1787 ( 
.A1(n_1748),
.A2(n_1718),
.A3(n_1682),
.B1(n_1666),
.B2(n_1663),
.B3(n_1679),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1740),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1724),
.A2(n_1658),
.B1(n_1693),
.B2(n_1698),
.Y(n_1789)
);

NAND2xp33_ASAP7_75t_R g1790 ( 
.A(n_1743),
.B(n_1664),
.Y(n_1790)
);

AO21x2_ASAP7_75t_L g1791 ( 
.A1(n_1745),
.A2(n_1758),
.B(n_1763),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1728),
.B(n_1698),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1747),
.B(n_1717),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1751),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1746),
.B(n_1709),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1746),
.B(n_1709),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1746),
.B(n_1709),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1728),
.B(n_1720),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1740),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1724),
.B(n_1683),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1756),
.B(n_1709),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1729),
.B(n_1717),
.Y(n_1802)
);

INVxp67_ASAP7_75t_SL g1803 ( 
.A(n_1751),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1733),
.B(n_1706),
.Y(n_1804)
);

NAND3xp33_ASAP7_75t_L g1805 ( 
.A(n_1752),
.B(n_1658),
.C(n_1674),
.Y(n_1805)
);

INVx4_ASAP7_75t_L g1806 ( 
.A(n_1743),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1768),
.B(n_1754),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1788),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1798),
.B(n_1733),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1791),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1798),
.B(n_1731),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1801),
.B(n_1795),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1801),
.B(n_1760),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1770),
.B(n_1758),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1768),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1801),
.B(n_1760),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1795),
.B(n_1760),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1792),
.B(n_1766),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1792),
.B(n_1731),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1795),
.B(n_1762),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1776),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1796),
.B(n_1797),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1783),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1796),
.B(n_1722),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1796),
.B(n_1722),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1797),
.B(n_1755),
.Y(n_1826)
);

INVxp67_ASAP7_75t_L g1827 ( 
.A(n_1781),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1799),
.B(n_1741),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1766),
.B(n_1742),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1770),
.B(n_1744),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1797),
.B(n_1755),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1767),
.B(n_1750),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1767),
.B(n_1750),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1767),
.B(n_1739),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1776),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1799),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1770),
.B(n_1752),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1776),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1783),
.Y(n_1839)
);

NAND2x1_ASAP7_75t_L g1840 ( 
.A(n_1806),
.B(n_1725),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1772),
.B(n_1742),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1773),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1770),
.B(n_1735),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1770),
.B(n_1735),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1770),
.B(n_1738),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1775),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1775),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1777),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1808),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1827),
.B(n_1815),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1827),
.B(n_1781),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1815),
.B(n_1779),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1807),
.B(n_1800),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1834),
.B(n_1770),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1808),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1809),
.B(n_1782),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1846),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1836),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1807),
.B(n_1779),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1809),
.B(n_1785),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1834),
.B(n_1806),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_1811),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1809),
.B(n_1785),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1834),
.B(n_1832),
.Y(n_1864)
);

NAND2x1_ASAP7_75t_L g1865 ( 
.A(n_1830),
.B(n_1806),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1832),
.B(n_1806),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1832),
.B(n_1806),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1836),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1811),
.B(n_1803),
.Y(n_1869)
);

NOR2x1p5_ASAP7_75t_L g1870 ( 
.A(n_1840),
.B(n_1805),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1833),
.B(n_1782),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1828),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1830),
.B(n_1771),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1837),
.A2(n_1805),
.B1(n_1793),
.B2(n_1789),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1833),
.B(n_1780),
.Y(n_1875)
);

AND2x2_ASAP7_75t_SL g1876 ( 
.A(n_1830),
.B(n_1787),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1811),
.B(n_1800),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1829),
.B(n_1800),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1828),
.Y(n_1879)
);

INVx2_ASAP7_75t_SL g1880 ( 
.A(n_1830),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1810),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1833),
.B(n_1787),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1843),
.B(n_1780),
.Y(n_1883)
);

BUFx2_ASAP7_75t_SL g1884 ( 
.A(n_1837),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1846),
.B(n_1803),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1810),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1810),
.Y(n_1887)
);

INVxp67_ASAP7_75t_L g1888 ( 
.A(n_1823),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1823),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1842),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1829),
.B(n_1802),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1843),
.B(n_1844),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1810),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1842),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1810),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1842),
.Y(n_1896)
);

INVx5_ASAP7_75t_L g1897 ( 
.A(n_1814),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1857),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1849),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1862),
.B(n_1829),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1849),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1864),
.Y(n_1902)
);

NAND2x1p5_ASAP7_75t_L g1903 ( 
.A(n_1870),
.B(n_1840),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1856),
.B(n_1841),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1864),
.B(n_1830),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1862),
.B(n_1813),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1855),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1871),
.B(n_1812),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1854),
.B(n_1814),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1850),
.B(n_1877),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1855),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1871),
.B(n_1812),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1858),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1854),
.B(n_1812),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1870),
.B(n_1814),
.Y(n_1915)
);

INVxp67_ASAP7_75t_SL g1916 ( 
.A(n_1851),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1882),
.B(n_1813),
.Y(n_1917)
);

OAI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1876),
.A2(n_1822),
.B1(n_1789),
.B2(n_1793),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1889),
.B(n_1813),
.Y(n_1919)
);

AOI211xp5_ASAP7_75t_L g1920 ( 
.A1(n_1874),
.A2(n_1822),
.B(n_1765),
.C(n_1821),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1884),
.B(n_1843),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1889),
.B(n_1816),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1876),
.B(n_1816),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1874),
.A2(n_1774),
.B1(n_1838),
.B2(n_1821),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1858),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1877),
.B(n_1891),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1884),
.B(n_1844),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1860),
.B(n_1841),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1868),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1868),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1876),
.B(n_1814),
.Y(n_1931)
);

OAI33xp33_ASAP7_75t_L g1932 ( 
.A1(n_1888),
.A2(n_1835),
.A3(n_1838),
.B1(n_1821),
.B2(n_1818),
.B3(n_1848),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1880),
.B(n_1749),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1890),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1890),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1852),
.B(n_1816),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1860),
.B(n_1841),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1852),
.B(n_1820),
.Y(n_1938)
);

OAI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1918),
.A2(n_1786),
.B1(n_1835),
.B2(n_1821),
.Y(n_1939)
);

AOI221xp5_ASAP7_75t_L g1940 ( 
.A1(n_1924),
.A2(n_1835),
.B1(n_1838),
.B2(n_1822),
.C(n_1765),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1914),
.Y(n_1941)
);

OAI22xp33_ASAP7_75t_L g1942 ( 
.A1(n_1923),
.A2(n_1786),
.B1(n_1838),
.B2(n_1835),
.Y(n_1942)
);

INVxp67_ASAP7_75t_L g1943 ( 
.A(n_1933),
.Y(n_1943)
);

OAI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1931),
.A2(n_1774),
.B(n_1869),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1931),
.A2(n_1869),
.B(n_1863),
.Y(n_1945)
);

AOI221xp5_ASAP7_75t_L g1946 ( 
.A1(n_1924),
.A2(n_1881),
.B1(n_1886),
.B2(n_1895),
.C(n_1887),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1920),
.A2(n_1776),
.B1(n_1763),
.B2(n_1656),
.Y(n_1947)
);

AOI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1932),
.A2(n_1863),
.B(n_1885),
.Y(n_1948)
);

OAI21xp5_ASAP7_75t_SL g1949 ( 
.A1(n_1903),
.A2(n_1814),
.B(n_1875),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1916),
.B(n_1872),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1934),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1935),
.Y(n_1952)
);

O2A1O1Ixp33_ASAP7_75t_L g1953 ( 
.A1(n_1903),
.A2(n_1885),
.B(n_1794),
.C(n_1895),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1917),
.A2(n_1776),
.B1(n_1656),
.B2(n_1791),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1908),
.B(n_1872),
.Y(n_1955)
);

NAND2x1_ASAP7_75t_L g1956 ( 
.A(n_1915),
.B(n_1921),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1899),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1908),
.B(n_1875),
.Y(n_1958)
);

INVxp67_ASAP7_75t_SL g1959 ( 
.A(n_1933),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1912),
.B(n_1879),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1901),
.Y(n_1961)
);

AOI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1919),
.A2(n_1865),
.B(n_1873),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1907),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1912),
.B(n_1879),
.Y(n_1964)
);

AOI211xp5_ASAP7_75t_L g1965 ( 
.A1(n_1915),
.A2(n_1853),
.B(n_1880),
.C(n_1794),
.Y(n_1965)
);

A2O1A1Ixp33_ASAP7_75t_L g1966 ( 
.A1(n_1915),
.A2(n_1804),
.B(n_1853),
.C(n_1817),
.Y(n_1966)
);

OR2x6_ASAP7_75t_L g1967 ( 
.A(n_1910),
.B(n_1664),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1951),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1943),
.B(n_1910),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1952),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1957),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1942),
.A2(n_1906),
.B1(n_1791),
.B2(n_1900),
.Y(n_1972)
);

AOI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1939),
.A2(n_1914),
.B1(n_1927),
.B2(n_1921),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1961),
.Y(n_1974)
);

NAND3xp33_ASAP7_75t_SL g1975 ( 
.A(n_1947),
.B(n_1927),
.C(n_1922),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1963),
.Y(n_1976)
);

INVx2_ASAP7_75t_SL g1977 ( 
.A(n_1967),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1955),
.Y(n_1978)
);

AOI221xp5_ASAP7_75t_L g1979 ( 
.A1(n_1940),
.A2(n_1944),
.B1(n_1948),
.B2(n_1954),
.C(n_1946),
.Y(n_1979)
);

OAI21xp33_ASAP7_75t_L g1980 ( 
.A1(n_1959),
.A2(n_1904),
.B(n_1926),
.Y(n_1980)
);

AOI211xp5_ASAP7_75t_L g1981 ( 
.A1(n_1953),
.A2(n_1900),
.B(n_1938),
.C(n_1936),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1960),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1941),
.B(n_1898),
.Y(n_1983)
);

CKINVDCx14_ASAP7_75t_R g1984 ( 
.A(n_1967),
.Y(n_1984)
);

OAI31xp33_ASAP7_75t_L g1985 ( 
.A1(n_1966),
.A2(n_1937),
.A3(n_1928),
.B(n_1804),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1958),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1964),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1945),
.B(n_1902),
.Y(n_1988)
);

OAI21xp33_ASAP7_75t_L g1989 ( 
.A1(n_1967),
.A2(n_1902),
.B(n_1937),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1956),
.Y(n_1990)
);

AOI21xp33_ASAP7_75t_L g1991 ( 
.A1(n_1950),
.A2(n_1913),
.B(n_1911),
.Y(n_1991)
);

AOI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1979),
.A2(n_1975),
.B1(n_1972),
.B2(n_1973),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1969),
.B(n_1965),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_L g1994 ( 
.A(n_1984),
.B(n_1949),
.Y(n_1994)
);

INVxp33_ASAP7_75t_L g1995 ( 
.A(n_1969),
.Y(n_1995)
);

OAI322xp33_ASAP7_75t_L g1996 ( 
.A1(n_1988),
.A2(n_1925),
.A3(n_1930),
.B1(n_1929),
.B2(n_1962),
.C1(n_1881),
.C2(n_1895),
.Y(n_1996)
);

OAI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1984),
.A2(n_1949),
.B1(n_1909),
.B2(n_1897),
.Y(n_1997)
);

INVxp67_ASAP7_75t_L g1998 ( 
.A(n_1977),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1986),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1986),
.B(n_1905),
.Y(n_2000)
);

AOI22xp33_ASAP7_75t_SL g2001 ( 
.A1(n_1990),
.A2(n_1982),
.B1(n_1978),
.B2(n_1987),
.Y(n_2001)
);

AOI22xp33_ASAP7_75t_SL g2002 ( 
.A1(n_1968),
.A2(n_1881),
.B1(n_1886),
.B2(n_1887),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1980),
.B(n_1905),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1989),
.B(n_1981),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1983),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1970),
.Y(n_2006)
);

AOI21xp5_ASAP7_75t_L g2007 ( 
.A1(n_1985),
.A2(n_1865),
.B(n_1839),
.Y(n_2007)
);

NOR3x1_ASAP7_75t_L g2008 ( 
.A(n_1993),
.B(n_1974),
.C(n_1971),
.Y(n_2008)
);

XNOR2xp5_ASAP7_75t_L g2009 ( 
.A(n_1995),
.B(n_1972),
.Y(n_2009)
);

NOR3xp33_ASAP7_75t_L g2010 ( 
.A(n_1998),
.B(n_1991),
.C(n_1976),
.Y(n_2010)
);

NAND4xp25_ASAP7_75t_L g2011 ( 
.A(n_1994),
.B(n_1647),
.C(n_1909),
.D(n_1669),
.Y(n_2011)
);

NAND4xp25_ASAP7_75t_L g2012 ( 
.A(n_1992),
.B(n_2001),
.C(n_2004),
.D(n_2003),
.Y(n_2012)
);

NAND3xp33_ASAP7_75t_SL g2013 ( 
.A(n_2001),
.B(n_1648),
.C(n_1840),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1999),
.Y(n_2014)
);

AOI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1996),
.A2(n_1887),
.B(n_1886),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_2000),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_2006),
.Y(n_2017)
);

NAND4xp25_ASAP7_75t_SL g2018 ( 
.A(n_2007),
.B(n_1892),
.C(n_1883),
.D(n_1867),
.Y(n_2018)
);

O2A1O1Ixp33_ASAP7_75t_L g2019 ( 
.A1(n_2005),
.A2(n_1893),
.B(n_1859),
.C(n_1896),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_2002),
.B(n_1866),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_2002),
.B(n_1866),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2016),
.Y(n_2022)
);

OAI211xp5_ASAP7_75t_L g2023 ( 
.A1(n_2012),
.A2(n_1997),
.B(n_1897),
.C(n_1892),
.Y(n_2023)
);

NOR4xp25_ASAP7_75t_L g2024 ( 
.A(n_2014),
.B(n_1893),
.C(n_1896),
.D(n_1894),
.Y(n_2024)
);

AOI31xp33_ASAP7_75t_L g2025 ( 
.A1(n_2017),
.A2(n_1909),
.A3(n_1790),
.B(n_1883),
.Y(n_2025)
);

AOI31xp33_ASAP7_75t_L g2026 ( 
.A1(n_2009),
.A2(n_1790),
.A3(n_1867),
.B(n_1759),
.Y(n_2026)
);

NOR2x1_ASAP7_75t_L g2027 ( 
.A(n_2013),
.B(n_1894),
.Y(n_2027)
);

NOR4xp25_ASAP7_75t_L g2028 ( 
.A(n_2019),
.B(n_1893),
.C(n_1859),
.D(n_1861),
.Y(n_2028)
);

OAI221xp5_ASAP7_75t_L g2029 ( 
.A1(n_2010),
.A2(n_1897),
.B1(n_1878),
.B2(n_1778),
.C(n_1784),
.Y(n_2029)
);

OAI31xp33_ASAP7_75t_L g2030 ( 
.A1(n_2023),
.A2(n_2015),
.A3(n_2020),
.B(n_2021),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2022),
.Y(n_2031)
);

AOI211xp5_ASAP7_75t_L g2032 ( 
.A1(n_2029),
.A2(n_2011),
.B(n_2018),
.C(n_2008),
.Y(n_2032)
);

NAND3xp33_ASAP7_75t_L g2033 ( 
.A(n_2027),
.B(n_1897),
.C(n_1839),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_2028),
.B(n_1897),
.Y(n_2034)
);

OAI211xp5_ASAP7_75t_SL g2035 ( 
.A1(n_2024),
.A2(n_1878),
.B(n_1661),
.C(n_1818),
.Y(n_2035)
);

AOI221xp5_ASAP7_75t_L g2036 ( 
.A1(n_2026),
.A2(n_1791),
.B1(n_1784),
.B2(n_1778),
.C(n_1897),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2025),
.Y(n_2037)
);

AOI21xp33_ASAP7_75t_L g2038 ( 
.A1(n_2023),
.A2(n_1791),
.B(n_1784),
.Y(n_2038)
);

XNOR2xp5_ASAP7_75t_L g2039 ( 
.A(n_2032),
.B(n_1677),
.Y(n_2039)
);

AND2x2_ASAP7_75t_SL g2040 ( 
.A(n_2037),
.B(n_1861),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_2031),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_2034),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2030),
.B(n_2033),
.Y(n_2043)
);

NAND2x1p5_ASAP7_75t_L g2044 ( 
.A(n_2038),
.B(n_1671),
.Y(n_2044)
);

OAI22xp5_ASAP7_75t_SL g2045 ( 
.A1(n_2035),
.A2(n_1778),
.B1(n_1784),
.B2(n_1818),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_2040),
.B(n_2036),
.Y(n_2046)
);

NOR3xp33_ASAP7_75t_L g2047 ( 
.A(n_2041),
.B(n_1670),
.C(n_1778),
.Y(n_2047)
);

OAI221xp5_ASAP7_75t_L g2048 ( 
.A1(n_2044),
.A2(n_1819),
.B1(n_1817),
.B2(n_1820),
.C(n_1769),
.Y(n_2048)
);

AOI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_2046),
.A2(n_2042),
.B(n_2039),
.Y(n_2049)
);

AOI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_2049),
.A2(n_2043),
.B1(n_2039),
.B2(n_2048),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2050),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_2050),
.A2(n_2045),
.B1(n_2047),
.B2(n_1819),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_2051),
.A2(n_2052),
.B1(n_1819),
.B2(n_1820),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2051),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_SL g2055 ( 
.A1(n_2054),
.A2(n_1847),
.B1(n_1848),
.B2(n_1802),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_2053),
.A2(n_1817),
.B(n_1826),
.Y(n_2056)
);

OAI21x1_ASAP7_75t_L g2057 ( 
.A1(n_2056),
.A2(n_1825),
.B(n_1824),
.Y(n_2057)
);

OAI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_2057),
.A2(n_2055),
.B(n_1831),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_2058),
.Y(n_2059)
);

OAI221xp5_ASAP7_75t_R g2060 ( 
.A1(n_2059),
.A2(n_1847),
.B1(n_1825),
.B2(n_1824),
.C(n_1831),
.Y(n_2060)
);

AOI211xp5_ASAP7_75t_L g2061 ( 
.A1(n_2060),
.A2(n_1676),
.B(n_1845),
.C(n_1602),
.Y(n_2061)
);


endmodule