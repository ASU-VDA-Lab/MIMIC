module fake_jpeg_22798_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_60),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_28),
.B1(n_31),
.B2(n_27),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_45),
.B1(n_44),
.B2(n_19),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_27),
.B1(n_31),
.B2(n_26),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_48),
.B1(n_27),
.B2(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_47),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_82),
.B1(n_86),
.B2(n_94),
.Y(n_109)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_70),
.Y(n_111)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_28),
.B1(n_24),
.B2(n_36),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_89),
.B1(n_93),
.B2(n_33),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_77),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_47),
.B(n_41),
.C(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_76),
.B(n_79),
.Y(n_122)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_39),
.B1(n_44),
.B2(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_87),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_43),
.B1(n_39),
.B2(n_36),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_38),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_17),
.B1(n_24),
.B2(n_36),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_91),
.Y(n_101)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_96),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_52),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_64),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_102),
.A2(n_32),
.B1(n_34),
.B2(n_33),
.Y(n_153)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_104),
.B(n_114),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_43),
.B1(n_32),
.B2(n_17),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_110),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_46),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_42),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_72),
.B(n_45),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_40),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_75),
.Y(n_133)
);

CKINVDCx12_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

OR2x4_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_19),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_35),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_46),
.B(n_42),
.C(n_37),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_19),
.B1(n_73),
.B2(n_37),
.Y(n_137)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_124),
.Y(n_147)
);

CKINVDCx12_ASAP7_75t_R g123 ( 
.A(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_125),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_92),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_24),
.C(n_32),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_128),
.B1(n_34),
.B2(n_46),
.Y(n_155)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_132),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_154),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_70),
.B1(n_85),
.B2(n_84),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_148),
.B1(n_127),
.B2(n_113),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_139),
.B1(n_153),
.B2(n_128),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_40),
.B1(n_38),
.B2(n_37),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_109),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_142),
.B(n_150),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_29),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_143),
.B(n_152),
.Y(n_175)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_145),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_38),
.B1(n_40),
.B2(n_33),
.Y(n_148)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_122),
.B(n_17),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_42),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_111),
.B(n_35),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_139),
.A2(n_104),
.B1(n_112),
.B2(n_101),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_160),
.A2(n_162),
.B1(n_167),
.B2(n_181),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_18),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_112),
.B1(n_101),
.B2(n_115),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_20),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_SL g216 ( 
.A1(n_165),
.A2(n_170),
.B(n_171),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_146),
.A2(n_110),
.B1(n_106),
.B2(n_100),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_100),
.B(n_129),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_168),
.A2(n_169),
.B(n_174),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_130),
.B(n_126),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_121),
.Y(n_173)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_25),
.B(n_20),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_131),
.B(n_108),
.C(n_121),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_187),
.B(n_188),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_124),
.B1(n_131),
.B2(n_108),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_135),
.A2(n_25),
.B1(n_108),
.B2(n_23),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_137),
.B1(n_149),
.B2(n_157),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_18),
.Y(n_183)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_143),
.B(n_9),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_186),
.B(n_157),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_138),
.A2(n_20),
.B(n_18),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_148),
.A2(n_152),
.B(n_142),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_172),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_190),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_150),
.C(n_141),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_207),
.C(n_161),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_134),
.Y(n_192)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_193),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_156),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_197),
.B(n_198),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_175),
.B(n_136),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_202),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_136),
.B(n_132),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_206),
.B(n_214),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_183),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_210),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_188),
.A2(n_132),
.B(n_20),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_175),
.B(n_8),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_23),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_180),
.B(n_187),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_217),
.B(n_219),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_163),
.A2(n_0),
.B(n_1),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_220),
.A2(n_176),
.B1(n_174),
.B2(n_171),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_223),
.C(n_226),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_166),
.C(n_178),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_166),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_243),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_178),
.C(n_167),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_204),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_176),
.C(n_185),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_233),
.C(n_213),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_220),
.B1(n_203),
.B2(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_176),
.C(n_185),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_176),
.B1(n_103),
.B2(n_23),
.Y(n_236)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_218),
.A2(n_103),
.B1(n_23),
.B2(n_2),
.Y(n_239)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_218),
.B(n_9),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_192),
.B(n_212),
.CI(n_195),
.CON(n_244),
.SN(n_244)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_244),
.B(n_212),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_191),
.B(n_9),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_243),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_230),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_250),
.A2(n_251),
.B(n_262),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_240),
.A2(n_199),
.B(n_214),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_199),
.B(n_206),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_260),
.B(n_263),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_258),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_235),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_259),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_193),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_205),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_264),
.A2(n_266),
.B(n_267),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_219),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_223),
.C(n_226),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_229),
.B(n_190),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_201),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_1),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_233),
.C(n_232),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_274),
.C(n_275),
.Y(n_296)
);

NOR3xp33_ASAP7_75t_SL g272 ( 
.A(n_253),
.B(n_225),
.C(n_237),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_279),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_247),
.A2(n_239),
.B1(n_242),
.B2(n_231),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_280),
.B1(n_10),
.B2(n_13),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_189),
.C(n_224),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_263),
.C(n_189),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_248),
.A2(n_236),
.B1(n_227),
.B2(n_241),
.Y(n_276)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_276),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_260),
.B(n_244),
.CI(n_238),
.CON(n_278),
.SN(n_278)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_255),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_209),
.C(n_244),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_209),
.B1(n_246),
.B2(n_4),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_251),
.A2(n_7),
.B(n_13),
.Y(n_282)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_261),
.Y(n_288)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_283),
.A2(n_252),
.B1(n_254),
.B2(n_265),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_289),
.A2(n_270),
.B1(n_285),
.B2(n_278),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_278),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_292),
.C(n_300),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_254),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_7),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_6),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_298),
.Y(n_309)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_1),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_275),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_299),
.A2(n_283),
.B1(n_271),
.B2(n_268),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_272),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_301),
.A2(n_296),
.B(n_11),
.Y(n_319)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_287),
.A2(n_277),
.B1(n_285),
.B2(n_273),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_304),
.B(n_308),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_312),
.C(n_292),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_286),
.A2(n_289),
.B1(n_294),
.B2(n_280),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_310),
.B(n_311),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_311),
.B(n_293),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_3),
.C(n_4),
.Y(n_312)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_317),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_300),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_306),
.C(n_312),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_320),
.B(n_321),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_301),
.A2(n_11),
.B(n_12),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_12),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_306),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_325),
.C(n_3),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_SL g324 ( 
.A(n_316),
.B(n_305),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_303),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_313),
.B(n_302),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_14),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_14),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_326),
.B(n_332),
.Y(n_335)
);

OAI21xp33_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_322),
.B(n_334),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_330),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_327),
.C(n_4),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_4),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_5),
.C(n_332),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_5),
.C(n_332),
.Y(n_341)
);


endmodule