module fake_jpeg_4858_n_209 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_1),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_29),
.B1(n_32),
.B2(n_19),
.Y(n_33)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_35),
.B(n_36),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_13),
.C(n_20),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_13),
.B1(n_14),
.B2(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_32),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_25),
.A2(n_14),
.B1(n_15),
.B2(n_20),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_19),
.B1(n_15),
.B2(n_26),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_24),
.A2(n_22),
.B1(n_14),
.B2(n_15),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_22),
.B1(n_16),
.B2(n_23),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_26),
.B(n_25),
.C(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_36),
.B(n_40),
.C(n_35),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_23),
.B1(n_39),
.B2(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_50),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_57),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_29),
.B1(n_24),
.B2(n_32),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_24),
.B1(n_27),
.B2(n_32),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_39),
.B1(n_38),
.B2(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_21),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_70),
.B1(n_75),
.B2(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_73),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_33),
.B1(n_39),
.B2(n_38),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_42),
.C(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_76),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_31),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_33),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_74),
.B1(n_39),
.B2(n_48),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_91),
.B1(n_70),
.B2(n_72),
.Y(n_93)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_59),
.B(n_63),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_73),
.B(n_61),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_56),
.C(n_30),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_75),
.Y(n_96)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_74),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_56),
.Y(n_87)
);

OR2x6_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_72),
.Y(n_97)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_66),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_91),
.B1(n_86),
.B2(n_88),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_52),
.B1(n_45),
.B2(n_44),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_62),
.B(n_64),
.Y(n_114)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_103),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_72),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_97),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_28),
.C(n_31),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_102),
.B(n_88),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_71),
.B1(n_75),
.B2(n_54),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_76),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_65),
.Y(n_120)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_90),
.B1(n_78),
.B2(n_87),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_82),
.B1(n_83),
.B2(n_71),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_113),
.B(n_114),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_124),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_27),
.B1(n_38),
.B2(n_37),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_83),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_58),
.B1(n_55),
.B2(n_85),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_98),
.B1(n_38),
.B2(n_80),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_96),
.C(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_55),
.B1(n_58),
.B2(n_38),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_50),
.B(n_107),
.C(n_38),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_84),
.B(n_21),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_103),
.B1(n_95),
.B2(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_134),
.C(n_135),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_138),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_93),
.B1(n_102),
.B2(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_140),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_115),
.B1(n_117),
.B2(n_27),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_98),
.C(n_37),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_37),
.C(n_101),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_77),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_37),
.C(n_43),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_113),
.C(n_43),
.Y(n_150)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_142),
.A2(n_121),
.B1(n_115),
.B2(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_124),
.B(n_114),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_149),
.A2(n_133),
.B(n_43),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_151),
.C(n_154),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_113),
.C(n_99),
.Y(n_151)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_156),
.B1(n_133),
.B2(n_142),
.Y(n_159)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_125),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_43),
.B1(n_77),
.B2(n_17),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_141),
.A2(n_43),
.B1(n_21),
.B2(n_3),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_139),
.B(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_135),
.B(n_137),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_166),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_148),
.B1(n_155),
.B2(n_153),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_157),
.B1(n_152),
.B2(n_143),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_136),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_1),
.Y(n_175)
);

AOI21x1_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_1),
.B(n_2),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_17),
.C(n_12),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_170),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_145),
.B(n_17),
.CI(n_2),
.CON(n_170),
.SN(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_162),
.B(n_6),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_168),
.C(n_169),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_179),
.Y(n_184)
);

OAI321xp33_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_170),
.A3(n_160),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_6),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_183),
.B(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_164),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_166),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_171),
.B(n_170),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_186),
.A2(n_8),
.B(n_9),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_163),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_1),
.C(n_2),
.Y(n_192)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_176),
.A3(n_172),
.B1(n_177),
.B2(n_167),
.C1(n_161),
.C2(n_174),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_8),
.B(n_10),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_163),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_191),
.B(n_192),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_184),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_188),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_196),
.B(n_11),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_195),
.A2(n_189),
.B(n_9),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_11),
.Y(n_202)
);

AOI21x1_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_8),
.B(n_10),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_202),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_203),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_3),
.C(n_4),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_197),
.A3(n_204),
.B1(n_11),
.B2(n_5),
.C1(n_3),
.C2(n_4),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_206),
.B(n_204),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_5),
.Y(n_209)
);


endmodule