module fake_jpeg_23943_n_282 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_282);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_0),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_22),
.C(n_31),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_42),
.B(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_16),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_21),
.B1(n_23),
.B2(n_20),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_47),
.A2(n_49),
.B1(n_58),
.B2(n_59),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_21),
.B1(n_20),
.B2(n_23),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_60),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_21),
.B1(n_23),
.B2(n_19),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_54),
.B1(n_38),
.B2(n_33),
.Y(n_78)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_52),
.B(n_56),
.Y(n_92)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_18),
.B1(n_19),
.B2(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_17),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_29),
.B(n_28),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_18),
.B1(n_19),
.B2(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_18),
.B1(n_32),
.B2(n_19),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_63),
.B(n_73),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_32),
.B1(n_18),
.B2(n_27),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_27),
.B1(n_31),
.B2(n_22),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_42),
.B1(n_40),
.B2(n_39),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_66),
.A2(n_75),
.B1(n_35),
.B2(n_30),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_22),
.B1(n_31),
.B2(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_29),
.B1(n_43),
.B2(n_38),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_74),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_42),
.B1(n_40),
.B2(n_43),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_71),
.A2(n_78),
.B1(n_81),
.B2(n_41),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_91),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_59),
.B1(n_54),
.B2(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_76),
.B(n_77),
.Y(n_122)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_83),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

CKINVDCx10_ASAP7_75t_R g121 ( 
.A(n_80),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_26),
.B1(n_17),
.B2(n_25),
.Y(n_81)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_35),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_38),
.B1(n_26),
.B2(n_34),
.Y(n_85)
);

OAI22x1_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_88),
.B1(n_89),
.B2(n_71),
.Y(n_101)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_90),
.Y(n_114)
);

OR2x2_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_24),
.Y(n_87)
);

NAND2x1_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_41),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_34),
.B1(n_33),
.B2(n_30),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_55),
.A2(n_30),
.B1(n_35),
.B2(n_11),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_11),
.B(n_15),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_48),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_96),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_9),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_98),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_116),
.B1(n_99),
.B2(n_66),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_41),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_104),
.B(n_117),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_111),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_106),
.A2(n_115),
.B1(n_79),
.B2(n_83),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_76),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_8),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_110),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_8),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_113),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_41),
.B1(n_36),
.B2(n_2),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_117),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_41),
.C(n_36),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_36),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_69),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_129),
.A2(n_115),
.B(n_104),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_132),
.Y(n_165)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_133),
.A2(n_137),
.B1(n_152),
.B2(n_109),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_140),
.Y(n_175)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_148),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_78),
.B1(n_99),
.B2(n_96),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_147),
.B1(n_128),
.B2(n_125),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_73),
.B1(n_72),
.B2(n_84),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_92),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_82),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_143),
.B(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_82),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_153),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_112),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_86),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_101),
.A2(n_87),
.B1(n_90),
.B2(n_74),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_100),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_117),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_41),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_164),
.B1(n_171),
.B2(n_146),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_107),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_160),
.B(n_163),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_119),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_169),
.C(n_144),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_142),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_153),
.A2(n_128),
.B1(n_127),
.B2(n_110),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_178),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_179),
.B1(n_136),
.B2(n_131),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_98),
.B1(n_77),
.B2(n_111),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_105),
.B(n_103),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_176),
.B(n_169),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_105),
.B(n_123),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_139),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_133),
.A2(n_123),
.B1(n_113),
.B2(n_36),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_140),
.B(n_36),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_36),
.Y(n_189)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_135),
.B(n_152),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_146),
.B(n_145),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_173),
.B(n_132),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_203),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_188),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_179),
.B1(n_164),
.B2(n_166),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_191),
.A2(n_194),
.B(n_174),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_202),
.B1(n_204),
.B2(n_182),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_0),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_0),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_195),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_199),
.C(n_200),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_1),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_41),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_41),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_138),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_194),
.C(n_196),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_159),
.A2(n_138),
.B1(n_36),
.B2(n_1),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_138),
.B1(n_2),
.B2(n_1),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_156),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_215),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_174),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_209),
.A2(n_211),
.B(n_217),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_218),
.B1(n_205),
.B2(n_203),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_156),
.B1(n_168),
.B2(n_162),
.Y(n_214)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_178),
.B1(n_167),
.B2(n_177),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_190),
.A2(n_168),
.B1(n_172),
.B2(n_162),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_167),
.Y(n_219)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_36),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_180),
.C(n_163),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_201),
.C(n_186),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_225),
.A2(n_233),
.B1(n_220),
.B2(n_224),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_208),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_227),
.B(n_235),
.Y(n_251)
);

OAI322xp33_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_188),
.A3(n_191),
.B1(n_195),
.B2(n_193),
.C1(n_197),
.C2(n_206),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_232),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_186),
.Y(n_230)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_165),
.B1(n_189),
.B2(n_1),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_165),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_9),
.B(n_3),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_236),
.A2(n_218),
.B(n_214),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_213),
.B(n_9),
.Y(n_237)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_2),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_226),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_247),
.B(n_235),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_230),
.A2(n_209),
.B(n_216),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_226),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_242),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_232),
.C(n_221),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_258),
.B(n_259),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_231),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_257),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_245),
.B(n_229),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_233),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_261),
.A2(n_243),
.B1(n_244),
.B2(n_234),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_251),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_264),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_241),
.Y(n_263)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_263),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_243),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_221),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_240),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_265),
.Y(n_271)
);

OAI211xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_267),
.B(n_268),
.C(n_260),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_272),
.A2(n_273),
.A3(n_209),
.B1(n_252),
.B2(n_234),
.C1(n_266),
.C2(n_239),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_275),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_269),
.A2(n_247),
.B(n_241),
.Y(n_275)
);

AOI321xp33_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_271),
.A3(n_270),
.B1(n_239),
.B2(n_216),
.C(n_6),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_278),
.C(n_3),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_SL g281 ( 
.A1(n_279),
.A2(n_280),
.B(n_13),
.C(n_4),
.Y(n_281)
);

OAI311xp33_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_12),
.A3(n_4),
.B1(n_5),
.C1(n_6),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_281),
.Y(n_282)
);


endmodule