module fake_jpeg_26501_n_105 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_9),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_25),
.Y(n_36)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_1),
.B(n_2),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_16),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_31),
.B(n_16),
.C(n_18),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_19),
.B1(n_13),
.B2(n_20),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_19),
.B1(n_15),
.B2(n_18),
.Y(n_32)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx12_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_24),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_19),
.B1(n_20),
.B2(n_13),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_16),
.C(n_18),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_36),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_29),
.B(n_38),
.Y(n_56)
);

OA21x2_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_29),
.B(n_35),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_34),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_29),
.B1(n_17),
.B2(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_23),
.B1(n_41),
.B2(n_30),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_56),
.B(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_54),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_57),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_55),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_24),
.C(n_46),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_67),
.C(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_72),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_14),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_18),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_63),
.C(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_75),
.B(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_12),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_58),
.B(n_3),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_83),
.B1(n_84),
.B2(n_21),
.Y(n_89)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_30),
.B(n_34),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_30),
.B1(n_33),
.B2(n_21),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_74),
.B1(n_73),
.B2(n_16),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_82),
.B1(n_12),
.B2(n_4),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_22),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_88),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_10),
.C(n_8),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_89),
.B(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_2),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_3),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_95),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_8),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_92),
.B(n_85),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_96),
.Y(n_100)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_93),
.B(n_5),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_102),
.B(n_6),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_90),
.B1(n_12),
.B2(n_6),
.Y(n_102)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_97),
.B(n_5),
.C(n_6),
.D(n_4),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);


endmodule