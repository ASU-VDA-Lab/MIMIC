module fake_aes_7735_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g11 ( .A(n_7), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_10), .B(n_8), .Y(n_12) );
INVxp67_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
BUFx10_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_7), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_1), .Y(n_16) );
NAND2xp33_ASAP7_75t_R g17 ( .A(n_6), .B(n_8), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_12), .A2(n_13), .B(n_16), .Y(n_18) );
O2A1O1Ixp33_ASAP7_75t_SL g19 ( .A1(n_13), .A2(n_0), .B(n_1), .C(n_2), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_14), .B(n_0), .Y(n_20) );
INVx1_ASAP7_75t_SL g21 ( .A(n_14), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g22 ( .A(n_14), .B(n_0), .Y(n_22) );
NOR3xp33_ASAP7_75t_SL g23 ( .A(n_20), .B(n_17), .C(n_15), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
NOR2xp33_ASAP7_75t_R g25 ( .A(n_21), .B(n_17), .Y(n_25) );
NOR2x1_ASAP7_75t_L g26 ( .A(n_24), .B(n_21), .Y(n_26) );
NOR2xp33_ASAP7_75t_R g27 ( .A(n_24), .B(n_22), .Y(n_27) );
HB1xp67_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
AOI31xp33_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_12), .A3(n_18), .B(n_23), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_26), .Y(n_30) );
AOI22xp33_ASAP7_75t_SL g31 ( .A1(n_30), .A2(n_27), .B1(n_14), .B2(n_12), .Y(n_31) );
OAI321xp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_11), .A3(n_2), .B1(n_1), .B2(n_4), .C(n_3), .Y(n_32) );
OAI221xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_29), .B1(n_11), .B2(n_2), .C(n_6), .Y(n_33) );
HB1xp67_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
OAI22xp5_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_11), .B1(n_9), .B2(n_10), .Y(n_35) );
AOI22xp5_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_34), .B1(n_11), .B2(n_5), .Y(n_36) );
endmodule