module real_jpeg_11104_n_18 (n_17, n_8, n_0, n_2, n_338, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_339, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_338;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_339;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_2),
.A2(n_25),
.B1(n_35),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_2),
.A2(n_60),
.B1(n_68),
.B2(n_69),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_2),
.A2(n_52),
.B1(n_53),
.B2(n_60),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_60),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_52),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_3),
.B(n_52),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_3),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_3),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_3),
.A2(n_30),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_3),
.B(n_30),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_32),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_3),
.A2(n_27),
.B(n_31),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_3),
.A2(n_25),
.B1(n_35),
.B2(n_117),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_4),
.A2(n_25),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_4),
.A2(n_34),
.B1(n_52),
.B2(n_53),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_4),
.A2(n_34),
.B1(n_68),
.B2(n_69),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_5),
.Y(n_94)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

BUFx6f_ASAP7_75t_SL g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_10),
.A2(n_68),
.B1(n_69),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_10),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_97),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_97),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_10),
.A2(n_25),
.B1(n_35),
.B2(n_97),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_11),
.A2(n_68),
.B1(n_69),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_11),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_133),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_133),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_11),
.A2(n_25),
.B1(n_35),
.B2(n_133),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_12),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_12),
.A2(n_68),
.B1(n_69),
.B2(n_104),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_104),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_12),
.A2(n_25),
.B1(n_35),
.B2(n_104),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_13),
.A2(n_25),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_13),
.A2(n_38),
.B1(n_68),
.B2(n_69),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_13),
.A2(n_38),
.B1(n_52),
.B2(n_53),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_14),
.A2(n_25),
.B1(n_35),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_14),
.A2(n_62),
.B1(n_68),
.B2(n_69),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_62),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_16),
.A2(n_68),
.B1(n_69),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_16),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_16),
.A2(n_52),
.B1(n_53),
.B2(n_92),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_92),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_16),
.A2(n_25),
.B1(n_35),
.B2(n_92),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_17),
.A2(n_68),
.B1(n_69),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_17),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_17),
.A2(n_52),
.B1(n_53),
.B2(n_152),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_17),
.A2(n_30),
.B1(n_31),
.B2(n_152),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_17),
.A2(n_25),
.B1(n_35),
.B2(n_152),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_32),
.B(n_33),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_23),
.A2(n_32),
.B1(n_37),
.B2(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_23),
.A2(n_32),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_24),
.A2(n_29),
.B1(n_59),
.B2(n_61),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_24),
.A2(n_29),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_24),
.A2(n_29),
.B1(n_215),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_24),
.A2(n_29),
.B1(n_240),
.B2(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_24),
.A2(n_29),
.B1(n_258),
.B2(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_24),
.A2(n_29),
.B1(n_59),
.B2(n_284),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_25),
.A2(n_26),
.B(n_117),
.C(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_49),
.Y(n_50)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_36),
.B(n_43),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_79),
.B(n_336),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_72),
.C(n_74),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_44),
.A2(n_45),
.B1(n_331),
.B2(n_333),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_57),
.C(n_63),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_46),
.A2(n_47),
.B1(n_63),
.B2(n_311),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_47)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_48),
.A2(n_51),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_48),
.A2(n_51),
.B1(n_143),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_48),
.A2(n_51),
.B1(n_160),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_48),
.A2(n_51),
.B1(n_200),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_48),
.A2(n_51),
.B1(n_211),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_48),
.A2(n_51),
.B1(n_237),
.B2(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_48),
.A2(n_51),
.B1(n_55),
.B2(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_50),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_51),
.B(n_117),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_52),
.B(n_54),
.Y(n_147)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_53),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_57),
.A2(n_58),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_63),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_63),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_67),
.B(n_71),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_67),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_64),
.A2(n_67),
.B1(n_103),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_64),
.A2(n_67),
.B1(n_130),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_64),
.A2(n_67),
.B1(n_139),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_64),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_64),
.A2(n_67),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_64),
.A2(n_67),
.B1(n_223),
.B2(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_64),
.A2(n_67),
.B1(n_232),
.B2(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_67),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_67),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_70),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_68),
.B(n_121),
.Y(n_120)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_71),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_72),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_76),
.A2(n_77),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_329),
.B(n_335),
.Y(n_79)
);

OAI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_302),
.A3(n_322),
.B1(n_327),
.B2(n_328),
.C(n_338),
.Y(n_80)
);

AOI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_248),
.A3(n_290),
.B1(n_296),
.B2(n_301),
.C(n_339),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_205),
.C(n_244),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_175),
.B(n_204),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_154),
.B(n_174),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_135),
.B(n_153),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_124),
.B(n_134),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_110),
.B(n_123),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_98),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_89),
.B(n_98),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_93),
.A2(n_94),
.B1(n_151),
.B2(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_114),
.B1(n_115),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_105),
.B2(n_109),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_109),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_102),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_105),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_118),
.B(n_122),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_116),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_115),
.B1(n_132),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_114),
.A2(n_115),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_114),
.A2(n_115),
.B1(n_186),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_114),
.A2(n_115),
.B1(n_220),
.B2(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_114),
.A2(n_115),
.B(n_230),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_117),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_126),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_129),
.C(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_137),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_140),
.CI(n_144),
.CON(n_137),
.SN(n_137)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_142),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_149),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_155),
.B(n_156),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_167),
.B2(n_168),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_170),
.C(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_161),
.B1(n_162),
.B2(n_166),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_159),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_164),
.C(n_166),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_169),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_170),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_176),
.B(n_177),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_190),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_179),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_179),
.B(n_189),
.C(n_190),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_184),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_201),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_198),
.B2(n_199),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_198),
.C(n_201),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_195),
.A2(n_197),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_196),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_203),
.Y(n_214)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_206),
.A2(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_225),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_207),
.B(n_225),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_218),
.C(n_224),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_217),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_212),
.B1(n_213),
.B2(n_216),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_210),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_SL g242 ( 
.A(n_212),
.B(n_216),
.C(n_217),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_224),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_221),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_242),
.B2(n_243),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_228),
.B(n_233),
.C(n_243),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_231),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_238),
.C(n_241),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_238),
.B1(n_239),
.B2(n_241),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_236),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_242),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_245),
.B(n_246),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_267),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_249),
.B(n_267),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_260),
.C(n_266),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_250),
.A2(n_251),
.B1(n_260),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_256),
.C(n_259),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_254),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_255),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_260),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_265),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_262),
.B1(n_283),
.B2(n_285),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_261),
.A2(n_283),
.B(n_286),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_263),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_263),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_264),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_288),
.B2(n_289),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_279),
.B2(n_280),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_270),
.B(n_280),
.C(n_289),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_275),
.B(n_278),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_275),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_277),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_278),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_278),
.A2(n_304),
.B1(n_313),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_286),
.B2(n_287),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_283),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_288),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_297),
.B(n_300),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_292),
.B(n_293),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_315),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_315),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_313),
.C(n_314),
.Y(n_303)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_304),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_306),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_311),
.C(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_317),
.C(n_321),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_309),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_323),
.B(n_324),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_334),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_334),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_331),
.Y(n_333)
);


endmodule