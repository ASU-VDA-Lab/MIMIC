module fake_jpeg_1483_n_208 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_208);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_1),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx11_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_78),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_0),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_69),
.B1(n_61),
.B2(n_70),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_84),
.B1(n_91),
.B2(n_74),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_90),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_70),
.B1(n_66),
.B2(n_67),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_66),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_65),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_66),
.B1(n_79),
.B2(n_80),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_102),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_97),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_62),
.C(n_54),
.Y(n_99)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_53),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_79),
.B1(n_80),
.B2(n_88),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_55),
.B1(n_68),
.B2(n_51),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_63),
.B1(n_58),
.B2(n_86),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_51),
.B1(n_68),
.B2(n_58),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_72),
.B1(n_56),
.B2(n_59),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_108),
.Y(n_116)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_87),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_53),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_85),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_64),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_126),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_71),
.B1(n_89),
.B2(n_72),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_115),
.B1(n_121),
.B2(n_129),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_76),
.B(n_89),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_132),
.B(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_108),
.A2(n_53),
.B1(n_57),
.B2(n_76),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_0),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_8),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_15),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_28),
.B(n_45),
.C(n_44),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_134),
.B(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_9),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_144),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_153),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_116),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_151),
.C(n_123),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_11),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_142),
.Y(n_154)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_145),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_95),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_95),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_12),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_13),
.B(n_14),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_17),
.B(n_18),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_13),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_150),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_32),
.C(n_43),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_36),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_163),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_138),
.A2(n_125),
.B1(n_132),
.B2(n_19),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_152),
.B(n_148),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_SL g181 ( 
.A1(n_158),
.A2(n_165),
.B(n_166),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_35),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_150),
.B1(n_153),
.B2(n_151),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_19),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_170),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_153),
.B(n_22),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_168),
.B(n_37),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_40),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_176),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_31),
.C(n_34),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_180),
.C(n_184),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_179),
.B(n_182),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_38),
.C(n_39),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_160),
.B(n_49),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_42),
.C(n_165),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_162),
.Y(n_185)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_167),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_181),
.B1(n_159),
.B2(n_171),
.Y(n_195)
);

OA21x2_ASAP7_75t_SL g191 ( 
.A1(n_177),
.A2(n_164),
.B(n_157),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_164),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_195),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_187),
.Y(n_194)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_194),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_186),
.B(n_190),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_197),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_201),
.A2(n_202),
.B(n_200),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_199),
.B(n_196),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_173),
.C(n_189),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_168),
.B(n_192),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_206),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_192),
.Y(n_208)
);


endmodule