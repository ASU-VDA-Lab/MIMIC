module fake_jpeg_26730_n_144 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_56),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_55),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_43),
.B1(n_47),
.B2(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_65),
.B1(n_62),
.B2(n_47),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_79),
.B1(n_83),
.B2(n_84),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_46),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_54),
.B1(n_58),
.B2(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_0),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_48),
.B1(n_50),
.B2(n_49),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_59),
.B1(n_56),
.B2(n_20),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_19),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_99),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_89),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_39),
.B1(n_18),
.B2(n_21),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_94),
.B1(n_96),
.B2(n_102),
.Y(n_112)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_1),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_97),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_94)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_22),
.B1(n_34),
.B2(n_33),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_4),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

AO22x1_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_5),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_5),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_15),
.B1(n_29),
.B2(n_26),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_100),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_7),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_99),
.B1(n_100),
.B2(n_95),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_86),
.B1(n_94),
.B2(n_99),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_117),
.B(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_116),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_88),
.Y(n_116)
);

INVxp33_ASAP7_75t_SL g117 ( 
.A(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_124),
.Y(n_130)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_127),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_121),
.B1(n_112),
.B2(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_124),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_130),
.C(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_128),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_135),
.B1(n_134),
.B2(n_127),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_13),
.C(n_25),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_10),
.B(n_23),
.Y(n_144)
);


endmodule