module real_jpeg_4938_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AND2x2_ASAP7_75t_L g143 ( 
.A(n_0),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_0),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_0),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_0),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_0),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_0),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_0),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_0),
.B(n_33),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_1),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_1),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_1),
.B(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_1),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_1),
.B(n_125),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_1),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_1),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_2),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_2),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_2),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_2),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g365 ( 
.A(n_2),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_2),
.B(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_3),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_3),
.B(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_3),
.B(n_204),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_3),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_3),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_3),
.B(n_57),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_3),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_3),
.B(n_52),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_4),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_4),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_4),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_4),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_4),
.B(n_353),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_4),
.B(n_410),
.Y(n_409)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_5),
.Y(n_100)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_5),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_5),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_5),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_5),
.Y(n_366)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_6),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_6),
.Y(n_433)
);

BUFx5_ASAP7_75t_L g473 ( 
.A(n_6),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_7),
.B(n_37),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_7),
.B(n_135),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_7),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_7),
.B(n_98),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_7),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_7),
.B(n_198),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_7),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_7),
.B(n_63),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_8),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_9),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_9),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g292 ( 
.A(n_9),
.B(n_202),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_9),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_9),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_9),
.B(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_9),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_9),
.B(n_503),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_10),
.Y(n_181)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_10),
.Y(n_490)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_11),
.Y(n_546)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_12),
.Y(n_127)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_12),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_12),
.Y(n_198)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_14),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_14),
.B(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_14),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_14),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_14),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_14),
.B(n_392),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_14),
.B(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_14),
.B(n_489),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_15),
.Y(n_95)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_15),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_15),
.Y(n_364)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_17),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_17),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_17),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_17),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_17),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_17),
.B(n_339),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_17),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_17),
.B(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_18),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_18),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_18),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_18),
.B(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_18),
.B(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_18),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_18),
.B(n_33),
.Y(n_289)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_545),
.B(n_547),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_79),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_78),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_45),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_45),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_35),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_26),
.A2(n_27),
.B1(n_36),
.B2(n_61),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_36),
.C(n_41),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_28),
.B(n_386),
.Y(n_385)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_29),
.Y(n_312)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_55),
.B1(n_56),
.B2(n_61),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_36),
.B(n_49),
.C(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_39),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_39),
.Y(n_319)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_40),
.Y(n_340)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_40),
.Y(n_412)
);

BUFx5_ASAP7_75t_L g442 ( 
.A(n_40),
.Y(n_442)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_40),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_74),
.C(n_76),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_46),
.B(n_535),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_62),
.C(n_64),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_47),
.A2(n_48),
.B1(n_531),
.B2(n_532),
.Y(n_530)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_65),
.C(n_70),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_55),
.A2(n_56),
.B1(n_70),
.B2(n_491),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_59),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_59),
.Y(n_355)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_60),
.Y(n_159)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_60),
.Y(n_176)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_60),
.Y(n_255)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_60),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_62),
.B(n_64),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_65),
.A2(n_66),
.B1(n_493),
.B2(n_494),
.Y(n_492)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_70),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_70),
.A2(n_444),
.B1(n_445),
.B2(n_491),
.Y(n_509)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_72),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

INVx11_ASAP7_75t_L g227 ( 
.A(n_73),
.Y(n_227)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_73),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_536),
.Y(n_535)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_76),
.Y(n_536)
);

AO21x1_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_463),
.B(n_538),
.Y(n_79)
);

OAI21x1_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_419),
.B(n_462),
.Y(n_80)
);

AOI21x1_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_374),
.B(n_418),
.Y(n_81)
);

OAI21x1_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_323),
.B(n_373),
.Y(n_82)
);

AOI21x1_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_282),
.B(n_322),
.Y(n_83)
);

AO21x1_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_207),
.B(n_281),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_191),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_86),
.B(n_191),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_130),
.B2(n_190),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_87),
.B(n_131),
.C(n_170),
.Y(n_321)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_108),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_89),
.B(n_109),
.C(n_129),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_101),
.C(n_105),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_90),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_196)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_93),
.Y(n_215)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_95),
.Y(n_204)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_100),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_101),
.B(n_105),
.Y(n_206)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_107),
.B(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_113),
.B1(n_128),
.B2(n_129),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B(n_112),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_111),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_112),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_112),
.B(n_287),
.C(n_296),
.Y(n_330)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_114),
.B(n_120),
.C(n_124),
.Y(n_320)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_126),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_127),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_127),
.Y(n_447)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_170),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_148),
.C(n_160),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_132),
.B(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_143),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_138),
.C(n_143),
.Y(n_189)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_149),
.B1(n_160),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_156),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_150),
.A2(n_151),
.B1(n_156),
.B2(n_157),
.Y(n_274)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_153),
.B(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_167),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_162),
.B(n_452),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_162),
.B(n_472),
.Y(n_471)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2x1_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_187),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_171),
.B(n_188),
.C(n_189),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_177),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_172),
.B(n_182),
.C(n_185),
.Y(n_296)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_175),
.Y(n_476)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_181),
.Y(n_351)
);

INVx3_ASAP7_75t_SL g452 ( 
.A(n_181),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_182),
.Y(n_186)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_184),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.C(n_205),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_192),
.B(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_195),
.B(n_205),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.C(n_199),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_196),
.B(n_197),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_199),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_203),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21x1_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_276),
.B(n_280),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_261),
.B(n_275),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_245),
.B(n_260),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_236),
.B(n_244),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_217),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_216),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_228),
.B2(n_229),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_223),
.C(n_228),
.Y(n_259)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_227),
.Y(n_306)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_234),
.Y(n_249)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_240),
.B(n_243),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_259),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_259),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_249),
.C(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_256),
.C(n_258),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_254),
.Y(n_258)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_264),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_271),
.C(n_272),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_278),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_321),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_321),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_298),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_286),
.C(n_298),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_295),
.B2(n_297),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_289),
.B(n_292),
.C(n_293),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_301),
.C(n_313),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_313),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_307),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_302),
.B(n_308),
.C(n_311),
.Y(n_357)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx6_ASAP7_75t_L g459 ( 
.A(n_306),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_311),
.Y(n_307)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_320),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_317),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_317),
.C(n_320),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_324),
.B(n_325),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_326),
.B(n_343),
.C(n_371),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_343),
.B1(n_371),
.B2(n_372),
.Y(n_327)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_328),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_331),
.B2(n_342),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_329),
.B(n_332),
.C(n_333),
.Y(n_376)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_331),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_341),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_335),
.B(n_338),
.C(n_341),
.Y(n_405)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_343),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_356),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_344),
.B(n_357),
.C(n_358),
.Y(n_403)
);

BUFx24_ASAP7_75t_SL g552 ( 
.A(n_344),
.Y(n_552)
);

FAx1_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_349),
.CI(n_352),
.CON(n_344),
.SN(n_344)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_345),
.B(n_349),
.C(n_352),
.Y(n_415)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx5_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_369),
.B2(n_370),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_365),
.B1(n_367),
.B2(n_368),
.Y(n_360)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_361),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_361),
.B(n_368),
.C(n_369),
.Y(n_388)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_365),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_365),
.A2(n_368),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_368),
.B(n_381),
.C(n_385),
.Y(n_430)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_417),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_375),
.B(n_417),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_376),
.B(n_378),
.C(n_401),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_401),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_380),
.B1(n_387),
.B2(n_400),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_379),
.B(n_388),
.C(n_389),
.Y(n_424)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_383),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_384),
.A2(n_385),
.B1(n_444),
.B2(n_445),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_384),
.B(n_437),
.C(n_444),
.Y(n_510)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_387),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_397),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_395),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_391),
.B(n_395),
.C(n_397),
.Y(n_449)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_403),
.B1(n_404),
.B2(n_416),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_405),
.C(n_406),
.Y(n_421)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_404),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_415),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_409),
.B1(n_413),
.B2(n_414),
.Y(n_407)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_408),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_409),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_413),
.C(n_428),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_409),
.A2(n_414),
.B1(n_432),
.B2(n_434),
.Y(n_431)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx6_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_414),
.B(n_430),
.C(n_434),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_415),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_461),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_420),
.B(n_461),
.Y(n_462)
);

BUFx24_ASAP7_75t_SL g553 ( 
.A(n_420),
.Y(n_553)
);

FAx1_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_422),
.CI(n_435),
.CON(n_420),
.SN(n_420)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_421),
.B(n_422),
.C(n_435),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_425),
.B2(n_426),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_423),
.B(n_427),
.C(n_429),
.Y(n_518)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_429),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_432),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_448),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_449),
.C(n_450),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_443),
.Y(n_436)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx6_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_442),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_444),
.B(n_488),
.C(n_491),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_453),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_451),
.B(n_455),
.C(n_460),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_454),
.A2(n_455),
.B1(n_456),
.B2(n_460),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g460 ( 
.A(n_454),
.Y(n_460)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

NOR3xp33_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_523),
.C(n_533),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_519),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_466),
.A2(n_542),
.B(n_543),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_467),
.B(n_512),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_467),
.B(n_512),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_484),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_468),
.B(n_485),
.C(n_507),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.C(n_482),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_469),
.B(n_514),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_470),
.A2(n_482),
.B1(n_483),
.B2(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_470),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_474),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_475),
.C(n_477),
.Y(n_498)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_477),
.Y(n_474)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_507),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_497),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_487),
.A2(n_492),
.B1(n_495),
.B2(n_496),
.Y(n_486)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_487),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_487),
.B(n_496),
.C(n_497),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_488),
.B(n_509),
.Y(n_508)
);

INVx6_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_492),
.Y(n_496)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_498),
.B(n_499),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_498),
.B(n_501),
.C(n_506),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_501),
.B1(n_502),
.B2(n_506),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_500),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_502),
.Y(n_501)
);

INVx8_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_510),
.C(n_511),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_508),
.B(n_517),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_511),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_516),
.C(n_518),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_516),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_518),
.B(n_521),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_522),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_520),
.B(n_522),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_524),
.B(n_541),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_526),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_525),
.B(n_526),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_528),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_527),
.B(n_529),
.C(n_530),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_530),
.Y(n_528)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

A2O1A1Ixp33_ASAP7_75t_L g538 ( 
.A1(n_533),
.A2(n_539),
.B(n_540),
.C(n_544),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_537),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_534),
.B(n_537),
.Y(n_544)
);

INVx13_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_546),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_550),
.Y(n_547)
);

BUFx12f_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);


endmodule