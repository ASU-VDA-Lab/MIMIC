module real_aes_144_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_726;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_782;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_713;
wire n_404;
wire n_598;
wire n_288;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_692;
wire n_789;
wire n_544;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_762;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_475;
wire n_554;
wire n_798;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g288 ( .A(n_0), .B(n_289), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_1), .A2(n_253), .B1(n_347), .B2(n_429), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_2), .A2(n_208), .B1(n_393), .B2(n_479), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_3), .A2(n_245), .B1(n_425), .B2(n_483), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_4), .A2(n_149), .B1(n_611), .B2(n_665), .Y(n_664) );
XNOR2x1_ASAP7_75t_L g661 ( .A(n_5), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_6), .B(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_7), .A2(n_23), .B1(n_325), .B2(n_333), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_8), .A2(n_114), .B1(n_366), .B2(n_368), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_9), .A2(n_175), .B1(n_597), .B2(n_598), .Y(n_596) );
AO22x2_ASAP7_75t_L g306 ( .A1(n_10), .A2(n_191), .B1(n_296), .B2(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g743 ( .A(n_10), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_11), .A2(n_192), .B1(n_392), .B2(n_393), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_12), .A2(n_111), .B1(n_348), .B2(n_389), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_13), .A2(n_48), .B1(n_456), .B2(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g631 ( .A(n_14), .Y(n_631) );
INVx1_ASAP7_75t_L g648 ( .A(n_15), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_16), .A2(n_237), .B1(n_771), .B2(n_772), .Y(n_770) );
INVx1_ASAP7_75t_L g627 ( .A(n_17), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_18), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_19), .A2(n_80), .B1(n_362), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_20), .A2(n_177), .B1(n_389), .B2(n_442), .Y(n_676) );
AO22x2_ASAP7_75t_L g303 ( .A1(n_21), .A2(n_58), .B1(n_296), .B2(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_21), .B(n_742), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_22), .A2(n_227), .B1(n_381), .B2(n_382), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_24), .A2(n_142), .B1(n_321), .B2(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_25), .A2(n_226), .B1(n_432), .B2(n_503), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_26), .A2(n_190), .B1(n_456), .B2(n_457), .Y(n_455) );
AO222x2_ASAP7_75t_SL g534 ( .A1(n_27), .A2(n_43), .B1(n_157), .B2(n_400), .C1(n_403), .C2(n_419), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_28), .A2(n_158), .B1(n_345), .B2(n_606), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_29), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_30), .A2(n_120), .B1(n_453), .B2(n_597), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_31), .A2(n_82), .B1(n_389), .B2(n_427), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_32), .A2(n_162), .B1(n_523), .B2(n_526), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_33), .A2(n_151), .B1(n_392), .B2(n_517), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_34), .A2(n_42), .B1(n_343), .B2(n_346), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_35), .A2(n_256), .B1(n_583), .B2(n_585), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_36), .A2(n_59), .B1(n_343), .B2(n_634), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_37), .A2(n_164), .B1(n_462), .B2(n_611), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_38), .A2(n_152), .B1(n_427), .B2(n_429), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_39), .A2(n_132), .B1(n_453), .B2(n_604), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_40), .A2(n_76), .B1(n_332), .B2(n_337), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_41), .A2(n_128), .B1(n_425), .B2(n_483), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_44), .A2(n_180), .B1(n_432), .B2(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_45), .A2(n_70), .B1(n_424), .B2(n_425), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_46), .A2(n_61), .B1(n_444), .B2(n_446), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_47), .A2(n_106), .B1(n_581), .B2(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_49), .A2(n_107), .B1(n_392), .B2(n_393), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_50), .A2(n_129), .B1(n_351), .B2(n_355), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_51), .A2(n_89), .B1(n_416), .B2(n_417), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_52), .A2(n_252), .B1(n_367), .B2(n_389), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_53), .A2(n_165), .B1(n_431), .B2(n_432), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_54), .A2(n_123), .B1(n_416), .B2(n_417), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_55), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_56), .A2(n_66), .B1(n_604), .B2(n_605), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_57), .A2(n_147), .B1(n_403), .B2(n_419), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_60), .A2(n_103), .B1(n_479), .B2(n_517), .Y(n_516) );
AO222x2_ASAP7_75t_SL g514 ( .A1(n_62), .A2(n_183), .B1(n_204), .B2(n_400), .C1(n_403), .C2(n_419), .Y(n_514) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_63), .A2(n_271), .B(n_280), .C(n_745), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_64), .A2(n_141), .B1(n_448), .B2(n_449), .Y(n_447) );
OA22x2_ASAP7_75t_L g677 ( .A1(n_65), .A2(n_678), .B1(n_679), .B2(n_700), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_65), .Y(n_678) );
INVx3_ASAP7_75t_L g296 ( .A(n_67), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_68), .A2(n_97), .B1(n_351), .B2(n_446), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_69), .A2(n_257), .B1(n_497), .B2(n_576), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_71), .A2(n_138), .B1(n_431), .B2(n_432), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_72), .A2(n_234), .B1(n_403), .B2(n_419), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_73), .A2(n_197), .B1(n_427), .B2(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g641 ( .A(n_74), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_75), .A2(n_186), .B1(n_565), .B2(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_77), .A2(n_214), .B1(n_321), .B2(n_713), .Y(n_777) );
AOI222xp33_ASAP7_75t_L g398 ( .A1(n_78), .A2(n_95), .B1(n_193), .B2(n_399), .C1(n_401), .C2(n_404), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_79), .A2(n_126), .B1(n_580), .B2(n_581), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_81), .A2(n_188), .B1(n_397), .B2(n_584), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g709 ( .A1(n_83), .A2(n_710), .B1(n_726), .B2(n_727), .Y(n_709) );
INVx1_ASAP7_75t_L g726 ( .A(n_83), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_84), .A2(n_241), .B1(n_425), .B2(n_483), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_85), .A2(n_160), .B1(n_309), .B2(n_316), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_86), .A2(n_94), .B1(n_389), .B2(n_427), .Y(n_498) );
INVx1_ASAP7_75t_SL g297 ( .A(n_87), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_87), .B(n_125), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_88), .A2(n_115), .B1(n_392), .B2(n_393), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_90), .A2(n_127), .B1(n_397), .B2(n_584), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_91), .A2(n_266), .B1(n_378), .B2(n_445), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_92), .A2(n_172), .B1(n_667), .B2(n_668), .Y(n_666) );
INVx2_ASAP7_75t_L g276 ( .A(n_93), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_96), .A2(n_136), .B1(n_441), .B2(n_442), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_98), .A2(n_218), .B1(n_416), .B2(n_477), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_99), .A2(n_130), .B1(n_403), .B2(n_404), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_100), .A2(n_146), .B1(n_431), .B2(n_432), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_101), .A2(n_179), .B1(n_600), .B2(n_602), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_102), .A2(n_194), .B1(n_441), .B2(n_442), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_104), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_105), .A2(n_135), .B1(n_584), .B2(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_108), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_109), .A2(n_118), .B1(n_370), .B2(n_572), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_110), .A2(n_239), .B1(n_311), .B2(n_316), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_112), .B(n_289), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_113), .A2(n_242), .B1(n_395), .B2(n_397), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_116), .A2(n_133), .B1(n_449), .B2(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_117), .A2(n_230), .B1(n_333), .B2(n_466), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_119), .A2(n_182), .B1(n_459), .B2(n_461), .Y(n_458) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_121), .A2(n_558), .B(n_586), .Y(n_557) );
INVx1_ASAP7_75t_L g588 ( .A(n_121), .Y(n_588) );
AOI22xp33_ASAP7_75t_SL g482 ( .A1(n_122), .A2(n_173), .B1(n_425), .B2(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_124), .A2(n_248), .B1(n_337), .B2(n_580), .Y(n_753) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_125), .A2(n_207), .B1(n_296), .B2(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g561 ( .A(n_131), .B(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_134), .A2(n_224), .B1(n_427), .B2(n_429), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_137), .A2(n_260), .B1(n_451), .B2(n_452), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_139), .A2(n_184), .B1(n_316), .B2(n_717), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_140), .A2(n_265), .B1(n_381), .B2(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_143), .Y(n_792) );
XOR2xp5_ASAP7_75t_L g766 ( .A(n_144), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g803 ( .A(n_144), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_145), .A2(n_268), .B1(n_352), .B2(n_378), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_148), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_150), .A2(n_217), .B1(n_321), .B2(n_325), .Y(n_320) );
INVx1_ASAP7_75t_L g298 ( .A(n_153), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_154), .A2(n_250), .B1(n_581), .B2(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g650 ( .A(n_155), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_156), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_159), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_161), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_163), .A2(n_225), .B1(n_385), .B2(n_386), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_166), .A2(n_251), .B1(n_381), .B2(n_449), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_167), .Y(n_793) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_168), .A2(n_747), .B1(n_748), .B2(n_762), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_168), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_169), .A2(n_255), .B1(n_456), .B2(n_466), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_170), .B(n_290), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_171), .B(n_290), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_174), .A2(n_235), .B1(n_359), .B2(n_362), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_176), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_178), .A2(n_187), .B1(n_355), .B2(n_575), .Y(n_574) );
AO22x1_ASAP7_75t_L g564 ( .A1(n_181), .A2(n_240), .B1(n_459), .B2(n_565), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_185), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_189), .A2(n_254), .B1(n_445), .B2(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_195), .B(n_289), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_196), .A2(n_202), .B1(n_429), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_198), .A2(n_222), .B1(n_348), .B2(n_500), .Y(n_499) );
XNOR2x1_ASAP7_75t_L g621 ( .A(n_199), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g615 ( .A(n_200), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_201), .A2(n_209), .B1(n_416), .B2(n_477), .Y(n_476) );
AOI221x1_ASAP7_75t_L g635 ( .A1(n_203), .A2(n_228), .B1(n_448), .B2(n_636), .C(n_637), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_205), .A2(n_206), .B1(n_656), .B2(n_657), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_210), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g626 ( .A(n_211), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_212), .A2(n_269), .B1(n_636), .B2(n_725), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_213), .A2(n_216), .B1(n_449), .B2(n_595), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_215), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_219), .A2(n_262), .B1(n_389), .B2(n_427), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_220), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_221), .B(n_290), .Y(n_718) );
AND2x4_ASAP7_75t_L g278 ( .A(n_223), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g739 ( .A(n_223), .Y(n_739) );
AO21x1_ASAP7_75t_L g801 ( .A1(n_223), .A2(n_274), .B(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g279 ( .A(n_229), .Y(n_279) );
AND2x2_ASAP7_75t_R g764 ( .A(n_229), .B(n_739), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_231), .B(n_399), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_232), .B(n_752), .Y(n_751) );
XNOR2x1_ASAP7_75t_L g285 ( .A(n_233), .B(n_286), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_236), .A2(n_264), .B1(n_429), .B2(n_488), .Y(n_487) );
INVxp67_ASAP7_75t_L g275 ( .A(n_238), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_243), .Y(n_691) );
XNOR2xp5_ASAP7_75t_L g437 ( .A(n_244), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g640 ( .A(n_246), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_247), .A2(n_263), .B1(n_431), .B2(n_432), .Y(n_527) );
INVx1_ASAP7_75t_L g630 ( .A(n_249), .Y(n_630) );
INVx1_ASAP7_75t_L g644 ( .A(n_258), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_259), .B(n_290), .Y(n_473) );
OA22x2_ASAP7_75t_L g373 ( .A1(n_261), .A2(n_374), .B1(n_375), .B2(n_405), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_261), .Y(n_374) );
AO21x2_ASAP7_75t_L g408 ( .A1(n_261), .A2(n_375), .B(n_409), .Y(n_408) );
AOI22x1_ASAP7_75t_L g511 ( .A1(n_267), .A2(n_512), .B1(n_528), .B2(n_529), .Y(n_511) );
INVx1_ASAP7_75t_L g529 ( .A(n_267), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_279), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g802 ( .A(n_279), .Y(n_802) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_552), .B1(n_734), .B2(n_735), .C(n_736), .Y(n_280) );
INVx1_ASAP7_75t_L g734 ( .A(n_281), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_435), .B1(n_550), .B2(n_551), .Y(n_281) );
INVx4_ASAP7_75t_L g550 ( .A(n_282), .Y(n_550) );
OA22x2_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_411), .B2(n_434), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_373), .B1(n_406), .B2(n_407), .Y(n_284) );
INVx1_ASAP7_75t_SL g406 ( .A(n_285), .Y(n_406) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_341), .Y(n_286) );
NAND4xp25_ASAP7_75t_L g287 ( .A(n_288), .B(n_308), .C(n_320), .D(n_331), .Y(n_287) );
BUFx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx4_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
INVx3_ASAP7_75t_L g563 ( .A(n_291), .Y(n_563) );
INVx3_ASAP7_75t_SL g647 ( .A(n_291), .Y(n_647) );
INVx4_ASAP7_75t_SL g671 ( .A(n_291), .Y(n_671) );
INVx3_ASAP7_75t_L g752 ( .A(n_291), .Y(n_752) );
BUFx2_ASAP7_75t_L g775 ( .A(n_291), .Y(n_775) );
INVx6_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_301), .Y(n_292) );
AND2x4_ASAP7_75t_L g328 ( .A(n_293), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g339 ( .A(n_293), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g393 ( .A(n_293), .B(n_340), .Y(n_393) );
AND2x4_ASAP7_75t_L g400 ( .A(n_293), .B(n_301), .Y(n_400) );
AND2x2_ASAP7_75t_L g417 ( .A(n_293), .B(n_329), .Y(n_417) );
AND2x2_ASAP7_75t_L g477 ( .A(n_293), .B(n_329), .Y(n_477) );
AND2x2_ASAP7_75t_L g517 ( .A(n_293), .B(n_340), .Y(n_517) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_299), .Y(n_293) );
AND2x2_ASAP7_75t_L g314 ( .A(n_294), .B(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_294), .Y(n_319) );
INVx2_ASAP7_75t_L g336 ( .A(n_294), .Y(n_336) );
OAI22x1_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B1(n_297), .B2(n_298), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g300 ( .A(n_296), .Y(n_300) );
INVx2_ASAP7_75t_L g304 ( .A(n_296), .Y(n_304) );
INVx1_ASAP7_75t_L g307 ( .A(n_296), .Y(n_307) );
INVx2_ASAP7_75t_L g315 ( .A(n_299), .Y(n_315) );
AND2x2_ASAP7_75t_L g335 ( .A(n_299), .B(n_336), .Y(n_335) );
BUFx2_ASAP7_75t_L g357 ( .A(n_299), .Y(n_357) );
AND2x4_ASAP7_75t_L g345 ( .A(n_301), .B(n_314), .Y(n_345) );
AND2x2_ASAP7_75t_L g361 ( .A(n_301), .B(n_335), .Y(n_361) );
AND2x4_ASAP7_75t_L g372 ( .A(n_301), .B(n_349), .Y(n_372) );
AND2x6_ASAP7_75t_L g429 ( .A(n_301), .B(n_335), .Y(n_429) );
AND2x2_ASAP7_75t_L g431 ( .A(n_301), .B(n_314), .Y(n_431) );
AND2x2_ASAP7_75t_L g503 ( .A(n_301), .B(n_314), .Y(n_503) );
AND2x2_ASAP7_75t_L g523 ( .A(n_301), .B(n_349), .Y(n_523) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_305), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x4_ASAP7_75t_L g313 ( .A(n_303), .B(n_305), .Y(n_313) );
AND2x2_ASAP7_75t_L g318 ( .A(n_303), .B(n_306), .Y(n_318) );
INVx1_ASAP7_75t_L g324 ( .A(n_303), .Y(n_324) );
INVxp67_ASAP7_75t_L g340 ( .A(n_305), .Y(n_340) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g323 ( .A(n_306), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g463 ( .A(n_312), .Y(n_463) );
BUFx3_ASAP7_75t_L g566 ( .A(n_312), .Y(n_566) );
BUFx5_ASAP7_75t_L g717 ( .A(n_312), .Y(n_717) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AND2x4_ASAP7_75t_L g334 ( .A(n_313), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g348 ( .A(n_313), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g392 ( .A(n_313), .B(n_335), .Y(n_392) );
AND2x4_ASAP7_75t_L g403 ( .A(n_313), .B(n_314), .Y(n_403) );
AND2x2_ASAP7_75t_L g479 ( .A(n_313), .B(n_335), .Y(n_479) );
AND2x2_ASAP7_75t_L g526 ( .A(n_313), .B(n_349), .Y(n_526) );
AND2x2_ASAP7_75t_L g322 ( .A(n_314), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g416 ( .A(n_314), .B(n_323), .Y(n_416) );
AND2x4_ASAP7_75t_L g349 ( .A(n_315), .B(n_336), .Y(n_349) );
INVx2_ASAP7_75t_L g460 ( .A(n_316), .Y(n_460) );
BUFx3_ASAP7_75t_L g772 ( .A(n_316), .Y(n_772) );
BUFx12f_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx3_ASAP7_75t_L g612 ( .A(n_317), .Y(n_612) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x4_ASAP7_75t_L g356 ( .A(n_318), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g367 ( .A(n_318), .B(n_349), .Y(n_367) );
AND2x2_ASAP7_75t_SL g404 ( .A(n_318), .B(n_319), .Y(n_404) );
AND2x2_ASAP7_75t_SL g419 ( .A(n_318), .B(n_319), .Y(n_419) );
AND2x4_ASAP7_75t_L g425 ( .A(n_318), .B(n_357), .Y(n_425) );
AND2x4_ASAP7_75t_L g432 ( .A(n_318), .B(n_349), .Y(n_432) );
BUFx6f_ASAP7_75t_SL g456 ( .A(n_321), .Y(n_456) );
INVx1_ASAP7_75t_L g686 ( .A(n_321), .Y(n_686) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx3_ASAP7_75t_L g396 ( .A(n_322), .Y(n_396) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_322), .Y(n_584) );
AND2x2_ASAP7_75t_L g354 ( .A(n_323), .B(n_335), .Y(n_354) );
AND2x4_ASAP7_75t_L g364 ( .A(n_323), .B(n_349), .Y(n_364) );
AND2x2_ASAP7_75t_L g424 ( .A(n_323), .B(n_335), .Y(n_424) );
AND2x6_ASAP7_75t_L g427 ( .A(n_323), .B(n_349), .Y(n_427) );
AND2x2_ASAP7_75t_SL g483 ( .A(n_323), .B(n_335), .Y(n_483) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_324), .Y(n_330) );
INVx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g457 ( .A(n_327), .Y(n_457) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx3_ASAP7_75t_L g397 ( .A(n_328), .Y(n_397) );
BUFx6f_ASAP7_75t_SL g509 ( .A(n_328), .Y(n_509) );
INVx1_ASAP7_75t_L g654 ( .A(n_328), .Y(n_654) );
BUFx4f_ASAP7_75t_L g713 ( .A(n_328), .Y(n_713) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx2_ASAP7_75t_L g656 ( .A(n_333), .Y(n_656) );
BUFx4f_ASAP7_75t_SL g779 ( .A(n_333), .Y(n_779) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx2_ASAP7_75t_L g580 ( .A(n_334), .Y(n_580) );
BUFx3_ASAP7_75t_L g667 ( .A(n_334), .Y(n_667) );
BUFx2_ASAP7_75t_L g715 ( .A(n_334), .Y(n_715) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_SL g466 ( .A(n_338), .Y(n_466) );
INVx2_ASAP7_75t_SL g581 ( .A(n_338), .Y(n_581) );
INVx2_ASAP7_75t_L g657 ( .A(n_338), .Y(n_657) );
INVx2_ASAP7_75t_L g668 ( .A(n_338), .Y(n_668) );
INVx6_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND4xp25_ASAP7_75t_L g341 ( .A(n_342), .B(n_350), .C(n_358), .D(n_365), .Y(n_341) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g441 ( .A(n_344), .Y(n_441) );
INVx3_ASAP7_75t_L g604 ( .A(n_344), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_344), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_344), .A2(n_782), .B1(n_783), .B2(n_784), .Y(n_781) );
INVx6_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx3_ASAP7_75t_L g385 ( .A(n_345), .Y(n_385) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g573 ( .A(n_347), .Y(n_573) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g387 ( .A(n_348), .Y(n_387) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_348), .Y(n_453) );
BUFx3_ASAP7_75t_L g634 ( .A(n_348), .Y(n_634) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g639 ( .A(n_352), .Y(n_639) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g601 ( .A(n_353), .Y(n_601) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_354), .Y(n_445) );
BUFx3_ASAP7_75t_L g576 ( .A(n_354), .Y(n_576) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx5_ASAP7_75t_SL g379 ( .A(n_356), .Y(n_379) );
BUFx2_ASAP7_75t_L g446 ( .A(n_356), .Y(n_446) );
BUFx3_ASAP7_75t_L g497 ( .A(n_356), .Y(n_497) );
INVx2_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx3_ASAP7_75t_L g381 ( .A(n_360), .Y(n_381) );
INVx2_ASAP7_75t_L g570 ( .A(n_360), .Y(n_570) );
INVx2_ASAP7_75t_SL g723 ( .A(n_360), .Y(n_723) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g451 ( .A(n_361), .Y(n_451) );
BUFx2_ASAP7_75t_L g595 ( .A(n_361), .Y(n_595) );
INVx1_ASAP7_75t_L g628 ( .A(n_362), .Y(n_628) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g382 ( .A(n_363), .Y(n_382) );
INVx2_ASAP7_75t_L g449 ( .A(n_363), .Y(n_449) );
INVx2_ASAP7_75t_SL g759 ( .A(n_363), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_363), .A2(n_786), .B1(n_787), .B2(n_789), .Y(n_785) );
INVx8_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
BUFx3_ASAP7_75t_L g442 ( .A(n_367), .Y(n_442) );
BUFx3_ASAP7_75t_L g606 ( .A(n_367), .Y(n_606) );
BUFx2_ASAP7_75t_SL g636 ( .A(n_367), .Y(n_636) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g725 ( .A(n_370), .Y(n_725) );
INVx4_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx3_ASAP7_75t_L g389 ( .A(n_371), .Y(n_389) );
INVx3_ASAP7_75t_SL g448 ( .A(n_371), .Y(n_448) );
INVx2_ASAP7_75t_L g597 ( .A(n_371), .Y(n_597) );
INVx8_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_374), .Y(n_410) );
INVx1_ASAP7_75t_L g405 ( .A(n_375), .Y(n_405) );
NOR2x1_ASAP7_75t_SL g409 ( .A(n_375), .B(n_410), .Y(n_409) );
NAND4xp75_ASAP7_75t_L g375 ( .A(n_376), .B(n_383), .C(n_390), .D(n_398), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_380), .Y(n_376) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g602 ( .A(n_379), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_379), .A2(n_638), .B1(n_640), .B2(n_641), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_379), .A2(n_638), .B1(n_792), .B2(n_793), .Y(n_791) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_388), .Y(n_383) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_386), .Y(n_598) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g488 ( .A(n_387), .Y(n_488) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_394), .Y(n_390) );
INVxp67_ASAP7_75t_L g690 ( .A(n_392), .Y(n_690) );
INVx4_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g434 ( .A(n_411), .Y(n_434) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
XNOR2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_433), .Y(n_412) );
NOR2x1_ASAP7_75t_L g413 ( .A(n_414), .B(n_422), .Y(n_413) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .C(n_420), .D(n_421), .Y(n_414) );
NAND4xp25_ASAP7_75t_L g422 ( .A(n_423), .B(n_426), .C(n_428), .D(n_430), .Y(n_422) );
INVx1_ASAP7_75t_L g501 ( .A(n_429), .Y(n_501) );
INVx1_ASAP7_75t_L g551 ( .A(n_435), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_467), .B1(n_548), .B2(n_549), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_437), .Y(n_548) );
NOR2xp67_ASAP7_75t_L g438 ( .A(n_439), .B(n_454), .Y(n_438) );
NAND4xp25_ASAP7_75t_L g439 ( .A(n_440), .B(n_443), .C(n_447), .D(n_450), .Y(n_439) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx3_ASAP7_75t_L g788 ( .A(n_451), .Y(n_788) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND4xp25_ASAP7_75t_L g454 ( .A(n_455), .B(n_458), .C(n_464), .D(n_465), .Y(n_454) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI222xp33_ASAP7_75t_L g643 ( .A1(n_460), .A2(n_644), .B1(n_645), .B2(n_648), .C1(n_649), .C2(n_650), .Y(n_643) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g649 ( .A(n_462), .Y(n_649) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g665 ( .A(n_463), .Y(n_665) );
INVx1_ASAP7_75t_L g771 ( .A(n_463), .Y(n_771) );
INVx1_ASAP7_75t_L g549 ( .A(n_467), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_490), .B2(n_547), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
XOR2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_489), .Y(n_469) );
NAND2x1_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .Y(n_470) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
NOR2x1_ASAP7_75t_L g480 ( .A(n_481), .B(n_485), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
INVx1_ASAP7_75t_L g547 ( .A(n_490), .Y(n_547) );
XNOR2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_510), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
XNOR2x1_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
OR2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_504), .Y(n_494) );
NAND4xp25_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .C(n_499), .D(n_502), .Y(n_495) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND4xp25_ASAP7_75t_SL g504 ( .A(n_505), .B(n_506), .C(n_507), .D(n_508), .Y(n_504) );
BUFx2_ASAP7_75t_SL g585 ( .A(n_509), .Y(n_585) );
AO22x2_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_530), .B1(n_531), .B2(n_546), .Y(n_510) );
INVx1_ASAP7_75t_L g546 ( .A(n_511), .Y(n_546) );
INVx1_ASAP7_75t_L g528 ( .A(n_512), .Y(n_528) );
NAND2x1_ASAP7_75t_SL g512 ( .A(n_513), .B(n_519), .Y(n_512) );
NOR2xp67_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_518), .Y(n_515) );
INVxp67_ASAP7_75t_L g692 ( .A(n_517), .Y(n_692) );
NOR2x1_ASAP7_75t_L g519 ( .A(n_520), .B(n_524), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
XOR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_545), .Y(n_531) );
NAND2x1_ASAP7_75t_L g532 ( .A(n_533), .B(n_538), .Y(n_532) );
NOR2x1_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
NOR2x1_ASAP7_75t_L g538 ( .A(n_539), .B(n_542), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g735 ( .A(n_552), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_618), .B1(n_732), .B2(n_733), .Y(n_552) );
INVx1_ASAP7_75t_L g732 ( .A(n_553), .Y(n_732) );
OAI22xp5_ASAP7_75t_SL g553 ( .A1(n_554), .A2(n_589), .B1(n_590), .B2(n_616), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g617 ( .A(n_557), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_558), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_578), .Y(n_559) );
NOR3xp33_ASAP7_75t_SL g560 ( .A(n_561), .B(n_564), .C(n_567), .Y(n_560) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND4xp25_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .C(n_574), .D(n_577), .Y(n_567) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_573), .A2(n_795), .B1(n_796), .B2(n_797), .Y(n_794) );
BUFx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
XNOR2x1_ASAP7_75t_L g591 ( .A(n_592), .B(n_615), .Y(n_591) );
NOR2xp67_ASAP7_75t_L g592 ( .A(n_593), .B(n_607), .Y(n_592) );
NAND4xp25_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .C(n_599), .D(n_603), .Y(n_593) );
INVx2_ASAP7_75t_L g625 ( .A(n_595), .Y(n_625) );
INVx1_ASAP7_75t_L g796 ( .A(n_597), .Y(n_796) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVxp67_ASAP7_75t_L g784 ( .A(n_605), .Y(n_784) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND4xp25_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .C(n_613), .D(n_614), .Y(n_607) );
BUFx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g733 ( .A(n_618), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_704), .B1(n_730), .B2(n_731), .Y(n_618) );
INVx1_ASAP7_75t_L g731 ( .A(n_619), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_658), .B1(n_659), .B2(n_702), .Y(n_619) );
INVxp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g703 ( .A(n_621), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_635), .C(n_642), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_629), .Y(n_623) );
OAI22xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B1(n_627), .B2(n_628), .Y(n_624) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_651), .Y(n_642) );
INVx3_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_655), .Y(n_651) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_654), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_684) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AO22x2_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_677), .B2(n_701), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_672), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .C(n_669), .D(n_670), .Y(n_663) );
NAND4xp25_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .C(n_675), .D(n_676), .Y(n_672) );
INVx2_ASAP7_75t_L g701 ( .A(n_677), .Y(n_701) );
INVx1_ASAP7_75t_L g729 ( .A(n_677), .Y(n_729) );
INVx1_ASAP7_75t_L g700 ( .A(n_679), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_693), .Y(n_679) );
NOR3xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_684), .C(n_688), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_682), .B(n_683), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B1(n_691), .B2(n_692), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx2_ASAP7_75t_L g706 ( .A(n_701), .Y(n_706) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g730 ( .A(n_704), .Y(n_730) );
OA21x2_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B(n_728), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_709), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g727 ( .A(n_710), .Y(n_727) );
NOR2xp67_ASAP7_75t_L g710 ( .A(n_711), .B(n_719), .Y(n_710) );
NAND4xp25_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .C(n_716), .D(n_718), .Y(n_711) );
NAND4xp25_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .C(n_722), .D(n_724), .Y(n_719) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_740), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_738), .B(n_741), .Y(n_800) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
OAI222xp33_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_763), .B1(n_765), .B2(n_798), .C1(n_801), .C2(n_803), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_756), .Y(n_749) );
NAND4xp25_ASAP7_75t_L g750 ( .A(n_751), .B(n_753), .C(n_754), .D(n_755), .Y(n_750) );
NAND4xp25_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .C(n_760), .D(n_761), .Y(n_756) );
INVx1_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_780), .C(n_790), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_776), .Y(n_768) );
NAND2xp5_ASAP7_75t_SL g769 ( .A(n_770), .B(n_773), .Y(n_769) );
INVx2_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_785), .Y(n_780) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_794), .Y(n_790) );
INVx1_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
CKINVDCx6p67_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
endmodule