module fake_jpeg_18897_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_39),
.B(n_45),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_16),
.B1(n_15),
.B2(n_20),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_43),
.B1(n_27),
.B2(n_33),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_16),
.B1(n_26),
.B2(n_20),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_23),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_63),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_28),
.C(n_36),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_15),
.B1(n_13),
.B2(n_26),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_36),
.B(n_30),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_72),
.B(n_73),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_22),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_15),
.B1(n_27),
.B2(n_21),
.Y(n_65)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_30),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_2),
.B(n_3),
.Y(n_88)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_47),
.B(n_2),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_17),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

AOI22x1_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_59),
.B1(n_58),
.B2(n_54),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_58),
.B(n_66),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_96),
.B(n_86),
.C(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_93),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_70),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_97),
.C(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_98),
.B1(n_75),
.B2(n_85),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_53),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_84),
.C(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_102),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_90),
.B1(n_97),
.B2(n_89),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_74),
.B(n_82),
.C(n_86),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_96),
.B(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_107),
.Y(n_114)
);

A2O1A1O1Ixp25_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_81),
.B(n_88),
.C(n_62),
.D(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_113),
.Y(n_117)
);

AO221x1_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_83),
.B1(n_69),
.B2(n_64),
.C(n_52),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_14),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_104),
.B(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_116),
.B(n_118),
.Y(n_121)
);

OAI221xp5_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_14),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_5),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_114),
.C(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_122),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_108),
.C(n_68),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_10),
.Y(n_124)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

BUFx6f_ASAP7_75t_SL g127 ( 
.A(n_124),
.Y(n_127)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_11),
.B(n_121),
.C(n_125),
.D(n_126),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_11),
.Y(n_129)
);


endmodule