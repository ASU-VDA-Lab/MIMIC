module fake_jpeg_5186_n_61 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_61);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_61;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_38;
wire n_36;
wire n_31;
wire n_56;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_7),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_46),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_38),
.C(n_39),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_32),
.C(n_31),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_52),
.C(n_53),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_8),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_56),
.B(n_16),
.Y(n_57)
);

AOI322xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_55),
.A3(n_18),
.B1(n_20),
.B2(n_21),
.C1(n_22),
.C2(n_17),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_60),
.B(n_28),
.Y(n_61)
);


endmodule