module fake_jpeg_14277_n_31 (n_3, n_2, n_1, n_0, n_4, n_5, n_31);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_31;

wire n_13;
wire n_21;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_SL g6 ( 
.A(n_1),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx24_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx14_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_15),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_17),
.B1(n_18),
.B2(n_6),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_9),
.A2(n_1),
.B(n_3),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_7),
.B(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_9),
.A2(n_5),
.B1(n_8),
.B2(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_21),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_23),
.B(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_25),
.C(n_20),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_26),
.A2(n_21),
.B1(n_23),
.B2(n_18),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_28),
.B(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_17),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_10),
.B(n_8),
.C(n_15),
.Y(n_31)
);


endmodule