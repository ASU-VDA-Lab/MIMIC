module fake_jpeg_31633_n_509 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_509);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_509;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_21),
.B(n_7),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_54),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_7),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_25),
.B(n_7),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_58),
.B(n_76),
.Y(n_117)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_82),
.Y(n_107)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_25),
.B(n_6),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_23),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_30),
.B(n_6),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_88),
.B(n_99),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_19),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_93),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_6),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_30),
.B(n_10),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_43),
.B(n_10),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_50),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_64),
.A2(n_26),
.B1(n_49),
.B2(n_33),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g200 ( 
.A1(n_109),
.A2(n_63),
.B1(n_17),
.B2(n_41),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_35),
.B1(n_34),
.B2(n_36),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_111),
.A2(n_131),
.B1(n_145),
.B2(n_100),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_122),
.B(n_41),
.Y(n_205)
);

INVx6_ASAP7_75t_SL g123 ( 
.A(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_123),
.B(n_136),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_92),
.A2(n_35),
.B1(n_34),
.B2(n_89),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_103),
.B(n_43),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_135),
.B(n_150),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_56),
.A2(n_35),
.B1(n_41),
.B2(n_38),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_60),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_149),
.A2(n_152),
.B1(n_24),
.B2(n_20),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_103),
.B(n_51),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_61),
.A2(n_45),
.B1(n_52),
.B2(n_26),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_93),
.B(n_49),
.C(n_33),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_17),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_72),
.B(n_50),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_156),
.B(n_161),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_101),
.B(n_51),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_SL g162 ( 
.A(n_63),
.Y(n_162)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g249 ( 
.A(n_166),
.Y(n_249)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_113),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_185),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_175),
.Y(n_218)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_172),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_70),
.B(n_71),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_174),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_105),
.B(n_47),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_176),
.B(n_178),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_159),
.A2(n_94),
.B1(n_87),
.B2(n_81),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_177),
.A2(n_206),
.B1(n_216),
.B2(n_147),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_127),
.B(n_140),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_192),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_184),
.A2(n_190),
.B1(n_193),
.B2(n_114),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_109),
.B(n_152),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_109),
.A2(n_98),
.B1(n_97),
.B2(n_77),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_L g253 ( 
.A1(n_187),
.A2(n_195),
.B1(n_129),
.B2(n_158),
.Y(n_253)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_111),
.A2(n_91),
.B1(n_86),
.B2(n_84),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_110),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_130),
.A2(n_95),
.B1(n_75),
.B2(n_74),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_142),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_194),
.B(n_199),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_130),
.A2(n_23),
.B1(n_47),
.B2(n_45),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_196),
.Y(n_230)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_198),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_138),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_212),
.Y(n_226)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_112),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_201),
.B(n_202),
.Y(n_252)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_215),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_115),
.B(n_24),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_217),
.C(n_174),
.Y(n_247)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_144),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_208),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_138),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_213),
.Y(n_227)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_121),
.B(n_24),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_118),
.B(n_41),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_126),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_214),
.B(n_125),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_131),
.A2(n_38),
.B1(n_36),
.B2(n_20),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_106),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_114),
.B(n_24),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_223),
.A2(n_132),
.B1(n_146),
.B2(n_210),
.Y(n_285)
);

CKINVDCx12_ASAP7_75t_R g224 ( 
.A(n_178),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_224),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_168),
.B(n_165),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_238),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_236),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_141),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_185),
.A2(n_159),
.B1(n_164),
.B2(n_129),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_251),
.B1(n_253),
.B2(n_198),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_141),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_254),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_247),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_215),
.A2(n_145),
.B1(n_158),
.B2(n_148),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_170),
.B(n_143),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_200),
.B(n_148),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_226),
.Y(n_273)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_260),
.A2(n_268),
.B1(n_278),
.B2(n_282),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_224),
.A2(n_180),
.B1(n_196),
.B2(n_203),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_262),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_202),
.C(n_207),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_272),
.C(n_286),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_248),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_288),
.Y(n_297)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_237),
.A2(n_200),
.B1(n_181),
.B2(n_207),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_221),
.A2(n_217),
.B(n_189),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_269),
.A2(n_276),
.B(n_243),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_223),
.A2(n_172),
.B1(n_166),
.B2(n_204),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_270),
.A2(n_280),
.B(n_281),
.Y(n_321)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_202),
.C(n_171),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_273),
.A2(n_222),
.B1(n_235),
.B2(n_241),
.Y(n_309)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_251),
.A2(n_217),
.B1(n_208),
.B2(n_157),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_237),
.A2(n_192),
.B1(n_201),
.B2(n_167),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_249),
.A2(n_216),
.B1(n_197),
.B2(n_116),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_249),
.A2(n_220),
.B1(n_231),
.B2(n_245),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_237),
.A2(n_182),
.B1(n_186),
.B2(n_191),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_249),
.A2(n_106),
.B1(n_116),
.B2(n_163),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_283),
.A2(n_290),
.B1(n_169),
.B2(n_173),
.Y(n_323)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_229),
.Y(n_284)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_284),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_236),
.B1(n_233),
.B2(n_231),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_222),
.B(n_188),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_146),
.C(n_132),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_252),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_244),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_248),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_228),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_220),
.A2(n_179),
.B1(n_206),
.B2(n_36),
.Y(n_290)
);

AND2x2_ASAP7_75t_SL g293 ( 
.A(n_267),
.B(n_226),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_293),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_258),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_298),
.B(n_315),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_269),
.A2(n_221),
.B(n_257),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_299),
.A2(n_303),
.B(n_313),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_300),
.B(n_306),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_302),
.B(n_309),
.Y(n_350)
);

AOI32xp33_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_221),
.A3(n_252),
.B1(n_242),
.B2(n_228),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_304),
.A2(n_319),
.B1(n_276),
.B2(n_275),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_267),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_305),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_254),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_278),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_311),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_218),
.Y(n_311)
);

AOI32xp33_ASAP7_75t_L g313 ( 
.A1(n_291),
.A2(n_242),
.A3(n_218),
.B1(n_238),
.B2(n_227),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_282),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_314),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_275),
.B(n_227),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_316),
.A2(n_317),
.B1(n_285),
.B2(n_277),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_260),
.A2(n_149),
.B1(n_240),
.B2(n_230),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_262),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_318),
.B(n_259),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_273),
.A2(n_229),
.B1(n_240),
.B2(n_230),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_323),
.A2(n_277),
.B1(n_274),
.B2(n_271),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_325),
.A2(n_343),
.B1(n_323),
.B2(n_322),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_279),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_327),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_328),
.A2(n_346),
.B1(n_347),
.B2(n_349),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_292),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_329),
.B(n_333),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_330),
.A2(n_312),
.B1(n_316),
.B2(n_304),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_264),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_332),
.C(n_337),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_286),
.C(n_272),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_244),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_292),
.Y(n_334)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_334),
.Y(n_359)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_335),
.Y(n_362)
);

OAI21xp33_ASAP7_75t_L g336 ( 
.A1(n_311),
.A2(n_263),
.B(n_268),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_336),
.A2(n_299),
.B(n_293),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_263),
.C(n_287),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_294),
.Y(n_338)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_338),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_341),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_305),
.A2(n_266),
.B1(n_284),
.B2(n_229),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_345),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_307),
.A2(n_244),
.B1(n_256),
.B2(n_246),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_307),
.A2(n_256),
.B1(n_250),
.B2(n_246),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_302),
.B(n_250),
.C(n_219),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_353),
.C(n_319),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_317),
.A2(n_256),
.B1(n_219),
.B2(n_220),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_300),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_351),
.B(n_318),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_303),
.B(n_313),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_297),
.B(n_220),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_320),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_357),
.A2(n_343),
.B1(n_349),
.B2(n_347),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_326),
.A2(n_310),
.B1(n_314),
.B2(n_293),
.Y(n_358)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_358),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_340),
.B(n_297),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_360),
.B(n_329),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_351),
.B(n_344),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_361),
.B(n_371),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_331),
.B(n_302),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_372),
.Y(n_386)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_339),
.A2(n_326),
.B1(n_352),
.B2(n_344),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_365),
.A2(n_383),
.B1(n_322),
.B2(n_173),
.Y(n_398)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_367),
.Y(n_400)
);

AO21x1_ASAP7_75t_L g368 ( 
.A1(n_342),
.A2(n_299),
.B(n_321),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_368),
.B(n_382),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_339),
.B(n_293),
.Y(n_373)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_373),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_332),
.B(n_309),
.C(n_319),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_375),
.B(n_376),
.C(n_378),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_309),
.C(n_298),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_295),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_381),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_296),
.C(n_308),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_320),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_24),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_353),
.C(n_342),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_38),
.C(n_48),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_296),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_354),
.B(n_308),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_368),
.A2(n_324),
.B(n_330),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_385),
.B(n_395),
.Y(n_425)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_388),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_369),
.A2(n_321),
.B1(n_338),
.B2(n_335),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_373),
.A2(n_328),
.B1(n_324),
.B2(n_346),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_390),
.A2(n_398),
.B1(n_404),
.B2(n_355),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_392),
.A2(n_355),
.B1(n_367),
.B2(n_382),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_360),
.B(n_345),
.Y(n_393)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_393),
.Y(n_423)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_374),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_334),
.Y(n_397)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_397),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_363),
.B(n_125),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_406),
.Y(n_419)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_383),
.A2(n_38),
.B1(n_36),
.B2(n_0),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_368),
.A2(n_11),
.B(n_15),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_410),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_356),
.B(n_48),
.C(n_1),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_408),
.B(n_409),
.C(n_378),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_48),
.C(n_1),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_365),
.B(n_0),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_381),
.B(n_48),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_362),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_387),
.B(n_380),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_412),
.B(n_428),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_396),
.Y(n_414)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_414),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_415),
.B(n_429),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_376),
.C(n_372),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_422),
.C(n_426),
.Y(n_438)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_420),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_421),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_401),
.B(n_375),
.C(n_377),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_390),
.A2(n_364),
.B1(n_370),
.B2(n_384),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_394),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_386),
.B(n_371),
.C(n_384),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_386),
.B(n_370),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_393),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_362),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_391),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_388),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_359),
.C(n_1),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_433),
.B(n_359),
.C(n_397),
.Y(n_442)
);

XNOR2x1_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_444),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_433),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_447),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_450),
.Y(n_452)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_423),
.Y(n_443)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_443),
.Y(n_462)
);

XOR2x1_ASAP7_75t_L g444 ( 
.A(n_430),
.B(n_391),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_425),
.B(n_403),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_445),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_406),
.C(n_394),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_451),
.C(n_419),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_418),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_414),
.B(n_396),
.Y(n_448)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_448),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_424),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_400),
.C(n_409),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_449),
.B(n_431),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_453),
.B(n_458),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_440),
.A2(n_421),
.B1(n_413),
.B2(n_427),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_454),
.A2(n_5),
.B1(n_2),
.B2(n_3),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_464),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_457),
.B(n_404),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_440),
.A2(n_413),
.B1(n_420),
.B2(n_405),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_437),
.A2(n_405),
.B1(n_410),
.B2(n_392),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_459),
.B(n_454),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_428),
.C(n_426),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_465),
.C(n_451),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_439),
.B(n_412),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_419),
.C(n_415),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_434),
.A2(n_385),
.B(n_407),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_467),
.A2(n_416),
.B(n_400),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_471),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_456),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_470),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_442),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_474),
.C(n_476),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_473),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_446),
.C(n_439),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_460),
.A2(n_435),
.B(n_444),
.C(n_398),
.Y(n_475)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_475),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_436),
.C(n_408),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_477),
.B(n_478),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_5),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_5),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_480),
.B(n_460),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_481),
.A2(n_462),
.B1(n_466),
.B2(n_467),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_470),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_452),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_486),
.A2(n_472),
.B(n_474),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_489),
.B(n_476),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_SL g490 ( 
.A(n_475),
.B(n_461),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_490),
.B(n_480),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_492),
.A2(n_493),
.B(n_494),
.Y(n_501)
);

AOI21x1_ASAP7_75t_SL g499 ( 
.A1(n_495),
.A2(n_496),
.B(n_497),
.Y(n_499)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_486),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_483),
.A2(n_468),
.B(n_464),
.Y(n_497)
);

A2O1A1Ixp33_ASAP7_75t_SL g498 ( 
.A1(n_495),
.A2(n_490),
.B(n_491),
.C(n_484),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_498),
.A2(n_500),
.B(n_468),
.Y(n_503)
);

A2O1A1Ixp33_ASAP7_75t_SL g500 ( 
.A1(n_495),
.A2(n_485),
.B(n_488),
.C(n_487),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_499),
.B(n_488),
.Y(n_502)
);

OAI311xp33_ASAP7_75t_L g504 ( 
.A1(n_502),
.A2(n_503),
.A3(n_501),
.B1(n_2),
.C1(n_3),
.Y(n_504)
);

AOI321xp33_ASAP7_75t_L g505 ( 
.A1(n_504),
.A2(n_4),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_505),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_506),
.A2(n_4),
.B(n_12),
.Y(n_507)
);

XOR2x2_ASAP7_75t_L g508 ( 
.A(n_507),
.B(n_4),
.Y(n_508)
);

AO21x1_ASAP7_75t_L g509 ( 
.A1(n_508),
.A2(n_13),
.B(n_15),
.Y(n_509)
);


endmodule