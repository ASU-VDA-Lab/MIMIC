module fake_netlist_1_1004_n_1540 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_137, n_277, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_210, n_184, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1540, n_995);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_210;
input n_184;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1540;
output n_995;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_311;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_315;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1533;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1203;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_606;
wire n_332;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1275;
wire n_955;
wire n_1093;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_325;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1335;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_1531;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g311 ( .A(n_273), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_98), .Y(n_312) );
CKINVDCx14_ASAP7_75t_R g313 ( .A(n_113), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_210), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_239), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_204), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_185), .B(n_81), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_191), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_184), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_201), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_103), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_254), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_42), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_297), .Y(n_324) );
CKINVDCx14_ASAP7_75t_R g325 ( .A(n_302), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_296), .Y(n_326) );
INVxp33_ASAP7_75t_SL g327 ( .A(n_252), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_55), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_251), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_77), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_130), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_12), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_186), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_277), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_290), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_260), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_236), .Y(n_337) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_161), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_280), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_143), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_309), .Y(n_341) );
CKINVDCx16_ASAP7_75t_R g342 ( .A(n_74), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_220), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_117), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_247), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_303), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_310), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_109), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_305), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_165), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_291), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_101), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_150), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_171), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_174), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_237), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_284), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_192), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_49), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_222), .Y(n_360) );
CKINVDCx16_ASAP7_75t_R g361 ( .A(n_98), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_166), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_228), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_187), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_101), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_42), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_103), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_221), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_196), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_235), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_78), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_94), .Y(n_372) );
INVx2_ASAP7_75t_SL g373 ( .A(n_209), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_111), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_6), .Y(n_375) );
BUFx10_ASAP7_75t_L g376 ( .A(n_5), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_26), .Y(n_377) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_226), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_275), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_225), .Y(n_380) );
INVx1_ASAP7_75t_SL g381 ( .A(n_224), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_4), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_227), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_300), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_207), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_68), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_122), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_266), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_84), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_160), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_71), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_141), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_172), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_261), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_159), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_142), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_217), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_262), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_234), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_7), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_246), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_272), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_243), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_241), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_293), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_59), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_203), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_265), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_181), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_211), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_294), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_286), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_230), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_244), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_80), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_182), .Y(n_416) );
INVx2_ASAP7_75t_SL g417 ( .A(n_269), .Y(n_417) );
INVxp33_ASAP7_75t_L g418 ( .A(n_30), .Y(n_418) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_183), .Y(n_419) );
CKINVDCx16_ASAP7_75t_R g420 ( .A(n_89), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_249), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_264), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_140), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_177), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_90), .Y(n_425) );
CKINVDCx16_ASAP7_75t_R g426 ( .A(n_308), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_248), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_46), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_70), .Y(n_429) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_45), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_36), .Y(n_431) );
CKINVDCx16_ASAP7_75t_R g432 ( .A(n_77), .Y(n_432) );
BUFx2_ASAP7_75t_SL g433 ( .A(n_154), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_281), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_255), .Y(n_435) );
BUFx2_ASAP7_75t_L g436 ( .A(n_292), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_146), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_128), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_188), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_218), .Y(n_440) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_274), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_21), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_44), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_48), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_288), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_37), .Y(n_446) );
BUFx2_ASAP7_75t_L g447 ( .A(n_44), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_176), .Y(n_448) );
BUFx3_ASAP7_75t_L g449 ( .A(n_223), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_283), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_158), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_81), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_208), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_91), .Y(n_454) );
BUFx3_ASAP7_75t_L g455 ( .A(n_25), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_282), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_232), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_100), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_73), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_87), .Y(n_460) );
BUFx10_ASAP7_75t_L g461 ( .A(n_268), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_134), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_132), .Y(n_463) );
INVxp67_ASAP7_75t_SL g464 ( .A(n_129), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_93), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_152), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_259), .Y(n_467) );
INVxp67_ASAP7_75t_L g468 ( .A(n_162), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_133), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_180), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_6), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_168), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_123), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_82), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_306), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_11), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_3), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_307), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_276), .Y(n_479) );
INVxp67_ASAP7_75t_SL g480 ( .A(n_169), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_212), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_12), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_117), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_270), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_256), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_111), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_75), .Y(n_487) );
INVx1_ASAP7_75t_SL g488 ( .A(n_271), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_94), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_233), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_133), .Y(n_491) );
INVx3_ASAP7_75t_L g492 ( .A(n_461), .Y(n_492) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_318), .A2(n_144), .B(n_139), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_426), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_323), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_373), .B(n_0), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_313), .Y(n_497) );
AO22x1_ASAP7_75t_L g498 ( .A1(n_418), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_341), .B(n_1), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_461), .Y(n_500) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_318), .A2(n_147), .B(n_145), .Y(n_501) );
INVx3_ASAP7_75t_L g502 ( .A(n_461), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_313), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_360), .Y(n_504) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_360), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_323), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_353), .B(n_3), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_370), .B(n_4), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_374), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_418), .B(n_5), .Y(n_510) );
NOR2x1_ASAP7_75t_L g511 ( .A(n_455), .B(n_7), .Y(n_511) );
INVx4_ASAP7_75t_L g512 ( .A(n_436), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_342), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_441), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_360), .Y(n_515) );
INVx3_ASAP7_75t_L g516 ( .A(n_455), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_329), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_374), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_346), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_409), .B(n_8), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_473), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_361), .A2(n_11), .B1(n_9), .B2(n_10), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_420), .A2(n_15), .B1(n_13), .B2(n_14), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_360), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_417), .B(n_13), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_462), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_393), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_473), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_477), .Y(n_529) );
NOR2x1_ASAP7_75t_L g530 ( .A(n_462), .B(n_14), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_393), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_477), .B(n_15), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_432), .A2(n_18), .B1(n_16), .B2(n_17), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_366), .B(n_16), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_311), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_447), .B(n_491), .Y(n_536) );
BUFx2_ASAP7_75t_L g537 ( .A(n_497), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_535), .B(n_337), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_505), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_535), .B(n_337), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_516), .B(n_354), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_516), .B(n_354), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_505), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_497), .B(n_325), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_516), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_512), .B(n_334), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_517), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_532), .A2(n_330), .B1(n_332), .B2(n_312), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_532), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_516), .B(n_357), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_505), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_503), .B(n_325), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_526), .B(n_357), .Y(n_553) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_505), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_532), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_512), .B(n_448), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_526), .B(n_363), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_512), .B(n_468), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_492), .B(n_343), .Y(n_559) );
BUFx10_ASAP7_75t_L g560 ( .A(n_503), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_532), .A2(n_344), .B1(n_352), .B2(n_348), .Y(n_561) );
INVx5_ASAP7_75t_L g562 ( .A(n_505), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_505), .Y(n_563) );
BUFx10_ASAP7_75t_L g564 ( .A(n_519), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_526), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_492), .B(n_343), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_504), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_505), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_504), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_504), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_515), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_510), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_512), .B(n_475), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_515), .Y(n_574) );
AND3x1_ASAP7_75t_L g575 ( .A(n_522), .B(n_533), .C(n_523), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_515), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_494), .Y(n_577) );
BUFx3_ASAP7_75t_L g578 ( .A(n_493), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_524), .Y(n_579) );
BUFx4f_ASAP7_75t_L g580 ( .A(n_493), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_524), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_572), .B(n_544), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_572), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_573), .B(n_492), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_549), .A2(n_510), .B1(n_534), .B2(n_506), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_544), .B(n_492), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_564), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_544), .B(n_500), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_552), .B(n_500), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_552), .A2(n_510), .B1(n_519), .B2(n_534), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_573), .B(n_500), .Y(n_591) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_578), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_546), .B(n_502), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_548), .A2(n_388), .B1(n_395), .B2(n_329), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_564), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_560), .B(n_502), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_SL g597 ( .A1(n_556), .A2(n_496), .B(n_502), .C(n_520), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_552), .A2(n_519), .B1(n_534), .B2(n_514), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_558), .B(n_536), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_559), .B(n_536), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_549), .A2(n_506), .B1(n_509), .B2(n_495), .Y(n_601) );
INVx3_ASAP7_75t_L g602 ( .A(n_549), .Y(n_602) );
BUFx2_ASAP7_75t_L g603 ( .A(n_537), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_555), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_537), .B(n_499), .Y(n_605) );
AND2x6_ASAP7_75t_SL g606 ( .A(n_575), .B(n_499), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_560), .B(n_507), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_547), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_545), .Y(n_609) );
INVx2_ASAP7_75t_SL g610 ( .A(n_560), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_560), .B(n_508), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_566), .B(n_525), .Y(n_612) );
AND2x6_ASAP7_75t_L g613 ( .A(n_578), .B(n_511), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_561), .B(n_347), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_545), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_538), .B(n_327), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_565), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_561), .B(n_347), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_575), .A2(n_523), .B1(n_533), .B2(n_522), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_538), .B(n_351), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_540), .B(n_327), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_565), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_578), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_541), .Y(n_624) );
OAI22xp5_ASAP7_75t_SL g625 ( .A1(n_577), .A2(n_458), .B1(n_331), .B2(n_513), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_540), .A2(n_513), .B1(n_443), .B2(n_452), .C(n_438), .Y(n_626) );
INVx3_ASAP7_75t_L g627 ( .A(n_541), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_542), .B(n_355), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_580), .A2(n_501), .B(n_493), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_580), .A2(n_501), .B(n_493), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_580), .A2(n_509), .B1(n_518), .B2(n_495), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_550), .B(n_355), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_550), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_580), .A2(n_501), .B(n_493), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_553), .B(n_358), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_553), .B(n_358), .Y(n_636) );
AND2x6_ASAP7_75t_SL g637 ( .A(n_557), .B(n_359), .Y(n_637) );
HB1xp67_ASAP7_75t_SL g638 ( .A(n_567), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_567), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_570), .B(n_362), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_570), .B(n_376), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_581), .B(n_428), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_581), .A2(n_518), .B1(n_528), .B2(n_521), .Y(n_643) );
AO22x1_ASAP7_75t_L g644 ( .A1(n_571), .A2(n_438), .B1(n_443), .B2(n_428), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_576), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_576), .B(n_396), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_579), .B(n_405), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_579), .B(n_405), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_569), .B(n_407), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_574), .A2(n_395), .B1(n_478), .B2(n_388), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_574), .B(n_407), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_539), .A2(n_521), .B1(n_529), .B2(n_528), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_562), .B(n_484), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_568), .A2(n_478), .B1(n_454), .B2(n_452), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_539), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_539), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_543), .A2(n_529), .B1(n_530), .B2(n_511), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_543), .A2(n_530), .B1(n_371), .B2(n_377), .Y(n_658) );
BUFx8_ASAP7_75t_L g659 ( .A(n_543), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_562), .B(n_484), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_624), .A2(n_458), .B1(n_331), .B2(n_454), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_627), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_610), .B(n_464), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_611), .B(n_498), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_595), .B(n_490), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_608), .Y(n_666) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_592), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_607), .B(n_490), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_650), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_629), .A2(n_501), .B(n_378), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_603), .B(n_489), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_594), .B(n_489), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_599), .A2(n_321), .B1(n_365), .B2(n_328), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_599), .B(n_375), .Y(n_674) );
O2A1O1Ixp5_ASAP7_75t_L g675 ( .A1(n_634), .A2(n_338), .B(n_480), .C(n_419), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_633), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_630), .A2(n_501), .B(n_551), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_616), .B(n_382), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_638), .A2(n_372), .B1(n_391), .B2(n_386), .Y(n_679) );
INVxp67_ASAP7_75t_L g680 ( .A(n_654), .Y(n_680) );
AND2x2_ASAP7_75t_SL g681 ( .A(n_619), .B(n_317), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_597), .A2(n_563), .B(n_551), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_602), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_613), .A2(n_406), .B1(n_415), .B2(n_400), .Y(n_684) );
O2A1O1Ixp33_ASAP7_75t_L g685 ( .A1(n_582), .A2(n_429), .B(n_431), .C(n_425), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_616), .B(n_389), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_583), .Y(n_687) );
O2A1O1Ixp33_ASAP7_75t_L g688 ( .A1(n_600), .A2(n_442), .B(n_446), .C(n_444), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_659), .B(n_587), .Y(n_689) );
BUFx3_ASAP7_75t_L g690 ( .A(n_659), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_598), .B(n_459), .Y(n_691) );
OAI321xp33_ASAP7_75t_L g692 ( .A1(n_657), .A2(n_460), .A3(n_469), .B1(n_474), .B2(n_471), .C(n_465), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_621), .B(n_463), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_585), .A2(n_486), .B1(n_487), .B2(n_483), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_584), .A2(n_315), .B(n_314), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_584), .A2(n_317), .B(n_319), .C(n_316), .Y(n_696) );
BUFx8_ASAP7_75t_L g697 ( .A(n_641), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_591), .A2(n_322), .B(n_320), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_585), .B(n_476), .Y(n_699) );
OAI21xp5_ASAP7_75t_L g700 ( .A1(n_604), .A2(n_326), .B(n_324), .Y(n_700) );
INVx1_ASAP7_75t_SL g701 ( .A(n_642), .Y(n_701) );
NOR2xp33_ASAP7_75t_SL g702 ( .A(n_592), .B(n_376), .Y(n_702) );
BUFx6f_ASAP7_75t_L g703 ( .A(n_592), .Y(n_703) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_592), .Y(n_704) );
AND2x6_ASAP7_75t_L g705 ( .A(n_623), .B(n_349), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_590), .B(n_376), .Y(n_706) );
OAI21xp33_ASAP7_75t_L g707 ( .A1(n_620), .A2(n_379), .B(n_340), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_628), .B(n_383), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_586), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_588), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_614), .B(n_336), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_632), .B(n_390), .Y(n_712) );
AND2x4_ASAP7_75t_L g713 ( .A(n_596), .B(n_333), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_635), .B(n_392), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_589), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_591), .A2(n_339), .B(n_335), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_609), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_636), .B(n_421), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_593), .A2(n_350), .B(n_345), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_644), .B(n_17), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_593), .A2(n_369), .B(n_368), .Y(n_721) );
BUFx3_ASAP7_75t_L g722 ( .A(n_613), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_631), .A2(n_387), .B1(n_430), .B2(n_367), .Y(n_723) );
INVx1_ASAP7_75t_SL g724 ( .A(n_623), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_618), .B(n_356), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_637), .B(n_364), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_615), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_631), .A2(n_387), .B1(n_430), .B2(n_367), .Y(n_728) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_623), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_612), .B(n_479), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_606), .B(n_640), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_601), .B(n_481), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_601), .A2(n_387), .B1(n_430), .B2(n_367), .Y(n_733) );
AOI21x1_ASAP7_75t_L g734 ( .A1(n_617), .A2(n_394), .B(n_380), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_626), .A2(n_397), .B1(n_399), .B2(n_398), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_622), .A2(n_403), .B(n_402), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_639), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_645), .Y(n_738) );
NAND3xp33_ASAP7_75t_L g739 ( .A(n_658), .B(n_482), .C(n_412), .Y(n_739) );
O2A1O1Ixp33_ASAP7_75t_L g740 ( .A1(n_646), .A2(n_414), .B(n_416), .C(n_411), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_647), .B(n_381), .Y(n_741) );
O2A1O1Ixp33_ASAP7_75t_L g742 ( .A1(n_648), .A2(n_423), .B(n_424), .C(n_422), .Y(n_742) );
AOI21x1_ASAP7_75t_L g743 ( .A1(n_655), .A2(n_435), .B(n_427), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_613), .B(n_404), .Y(n_744) );
AOI21x1_ASAP7_75t_L g745 ( .A1(n_656), .A2(n_440), .B(n_439), .Y(n_745) );
CKINVDCx8_ASAP7_75t_R g746 ( .A(n_625), .Y(n_746) );
AND2x4_ASAP7_75t_L g747 ( .A(n_649), .B(n_450), .Y(n_747) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_651), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_657), .A2(n_453), .B1(n_457), .B2(n_456), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_643), .B(n_488), .Y(n_750) );
BUFx3_ASAP7_75t_L g751 ( .A(n_653), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_643), .B(n_482), .Y(n_752) );
CKINVDCx10_ASAP7_75t_R g753 ( .A(n_652), .Y(n_753) );
OAI21xp33_ASAP7_75t_L g754 ( .A1(n_660), .A2(n_472), .B(n_470), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_629), .A2(n_384), .B(n_363), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_627), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_611), .B(n_433), .Y(n_757) );
A2O1A1Ixp33_ASAP7_75t_SL g758 ( .A1(n_593), .A2(n_527), .B(n_531), .C(n_524), .Y(n_758) );
NOR2xp67_ASAP7_75t_L g759 ( .A(n_650), .B(n_18), .Y(n_759) );
OAI21x1_ASAP7_75t_L g760 ( .A1(n_629), .A2(n_401), .B(n_384), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_605), .B(n_19), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_624), .A2(n_410), .B1(n_413), .B2(n_408), .Y(n_762) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_629), .A2(n_413), .B(n_410), .Y(n_763) );
INVx3_ASAP7_75t_L g764 ( .A(n_659), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_603), .Y(n_765) );
NOR2xp33_ASAP7_75t_R g766 ( .A(n_608), .B(n_19), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_611), .B(n_349), .Y(n_767) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_608), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_611), .B(n_385), .Y(n_769) );
NAND2xp33_ASAP7_75t_L g770 ( .A(n_595), .B(n_393), .Y(n_770) );
BUFx2_ASAP7_75t_L g771 ( .A(n_603), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_624), .A2(n_437), .B1(n_466), .B2(n_445), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_627), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_624), .A2(n_445), .B1(n_467), .B2(n_466), .Y(n_774) );
BUFx2_ASAP7_75t_L g775 ( .A(n_603), .Y(n_775) );
AOI21xp5_ASAP7_75t_L g776 ( .A1(n_629), .A2(n_485), .B(n_449), .Y(n_776) );
BUFx4f_ASAP7_75t_L g777 ( .A(n_603), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_611), .B(n_385), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_611), .B(n_20), .Y(n_779) );
AND2x4_ASAP7_75t_L g780 ( .A(n_610), .B(n_20), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_602), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_611), .A2(n_434), .B1(n_451), .B2(n_393), .Y(n_782) );
BUFx2_ASAP7_75t_L g783 ( .A(n_603), .Y(n_783) );
CKINVDCx8_ASAP7_75t_R g784 ( .A(n_608), .Y(n_784) );
AOI221xp5_ASAP7_75t_L g785 ( .A1(n_688), .A2(n_451), .B1(n_434), .B2(n_531), .C(n_527), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_677), .A2(n_554), .B(n_562), .Y(n_786) );
AND2x4_ASAP7_75t_L g787 ( .A(n_690), .B(n_22), .Y(n_787) );
A2O1A1Ixp33_ASAP7_75t_L g788 ( .A1(n_761), .A2(n_527), .B(n_451), .C(n_434), .Y(n_788) );
O2A1O1Ixp33_ASAP7_75t_SL g789 ( .A1(n_758), .A2(n_149), .B(n_151), .C(n_148), .Y(n_789) );
A2O1A1Ixp33_ASAP7_75t_L g790 ( .A1(n_740), .A2(n_562), .B(n_554), .C(n_24), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_676), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_701), .B(n_22), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_701), .B(n_23), .Y(n_793) );
AO22x2_ASAP7_75t_L g794 ( .A1(n_661), .A2(n_25), .B1(n_23), .B2(n_24), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_727), .Y(n_795) );
OAI21x1_ASAP7_75t_L g796 ( .A1(n_760), .A2(n_554), .B(n_155), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_680), .A2(n_28), .B1(n_26), .B2(n_27), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_687), .Y(n_798) );
AO31x2_ASAP7_75t_L g799 ( .A1(n_755), .A2(n_29), .A3(n_27), .B(n_28), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_717), .Y(n_800) );
OAI21xp5_ASAP7_75t_L g801 ( .A1(n_675), .A2(n_156), .B(n_153), .Y(n_801) );
OAI21x1_ASAP7_75t_L g802 ( .A1(n_682), .A2(n_554), .B(n_157), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_681), .B(n_29), .Y(n_803) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_765), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_669), .A2(n_32), .B1(n_30), .B2(n_31), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_709), .B(n_31), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_737), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_738), .Y(n_808) );
OAI21xp5_ASAP7_75t_L g809 ( .A1(n_763), .A2(n_32), .B(n_33), .Y(n_809) );
AOI221x1_ASAP7_75t_L g810 ( .A1(n_776), .A2(n_33), .B1(n_34), .B2(n_35), .C(n_36), .Y(n_810) );
NAND3xp33_ASAP7_75t_L g811 ( .A(n_696), .B(n_34), .C(n_35), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_771), .B(n_775), .Y(n_812) );
A2O1A1Ixp33_ASAP7_75t_L g813 ( .A1(n_742), .A2(n_39), .B(n_37), .C(n_38), .Y(n_813) );
BUFx10_ASAP7_75t_L g814 ( .A(n_780), .Y(n_814) );
CKINVDCx8_ASAP7_75t_R g815 ( .A(n_753), .Y(n_815) );
BUFx6f_ASAP7_75t_SL g816 ( .A(n_780), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_783), .B(n_40), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_662), .Y(n_818) );
O2A1O1Ixp33_ASAP7_75t_L g819 ( .A1(n_685), .A2(n_45), .B(n_41), .C(n_43), .Y(n_819) );
AND2x4_ASAP7_75t_L g820 ( .A(n_764), .B(n_41), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_756), .Y(n_821) );
INVx4_ASAP7_75t_L g822 ( .A(n_764), .Y(n_822) );
OAI21x1_ASAP7_75t_L g823 ( .A1(n_743), .A2(n_164), .B(n_163), .Y(n_823) );
OAI21x1_ASAP7_75t_L g824 ( .A1(n_745), .A2(n_170), .B(n_167), .Y(n_824) );
BUFx2_ASAP7_75t_L g825 ( .A(n_777), .Y(n_825) );
OA21x2_ASAP7_75t_L g826 ( .A1(n_734), .A2(n_175), .B(n_173), .Y(n_826) );
AO31x2_ASAP7_75t_L g827 ( .A1(n_723), .A2(n_47), .A3(n_43), .B(n_46), .Y(n_827) );
OAI21xp5_ASAP7_75t_L g828 ( .A1(n_664), .A2(n_47), .B(n_48), .Y(n_828) );
AOI22xp33_ASAP7_75t_SL g829 ( .A1(n_777), .A2(n_51), .B1(n_49), .B2(n_50), .Y(n_829) );
INVx1_ASAP7_75t_SL g830 ( .A(n_705), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_710), .B(n_50), .Y(n_831) );
AND2x4_ASAP7_75t_SL g832 ( .A(n_671), .B(n_52), .Y(n_832) );
OAI21x1_ASAP7_75t_L g833 ( .A1(n_752), .A2(n_179), .B(n_178), .Y(n_833) );
OAI21xp5_ASAP7_75t_L g834 ( .A1(n_715), .A2(n_52), .B(n_53), .Y(n_834) );
OAI22x1_ASAP7_75t_L g835 ( .A1(n_720), .A2(n_56), .B1(n_54), .B2(n_55), .Y(n_835) );
AOI221x1_ASAP7_75t_L g836 ( .A1(n_728), .A2(n_54), .B1(n_56), .B2(n_57), .C(n_58), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_674), .B(n_57), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_773), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g839 ( .A(n_672), .B(n_58), .Y(n_839) );
NOR2x1_ASAP7_75t_SL g840 ( .A(n_689), .B(n_60), .Y(n_840) );
NAND3x1_ASAP7_75t_L g841 ( .A(n_731), .B(n_60), .C(n_61), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_735), .B(n_61), .Y(n_842) );
OA21x2_ASAP7_75t_L g843 ( .A1(n_700), .A2(n_190), .B(n_189), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_779), .Y(n_844) );
CKINVDCx5p33_ASAP7_75t_R g845 ( .A(n_784), .Y(n_845) );
BUFx8_ASAP7_75t_L g846 ( .A(n_663), .Y(n_846) );
OAI22xp33_ASAP7_75t_L g847 ( .A1(n_746), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_847) );
AO31x2_ASAP7_75t_L g848 ( .A1(n_733), .A2(n_63), .A3(n_64), .B(n_65), .Y(n_848) );
AOI21xp5_ASAP7_75t_L g849 ( .A1(n_770), .A2(n_194), .B(n_193), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_694), .B(n_65), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_757), .Y(n_851) );
AOI21xp5_ASAP7_75t_L g852 ( .A1(n_712), .A2(n_197), .B(n_195), .Y(n_852) );
OAI21xp5_ASAP7_75t_L g853 ( .A1(n_695), .A2(n_199), .B(n_198), .Y(n_853) );
CKINVDCx8_ASAP7_75t_R g854 ( .A(n_666), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_767), .Y(n_855) );
INVx5_ASAP7_75t_L g856 ( .A(n_705), .Y(n_856) );
AO21x1_ASAP7_75t_L g857 ( .A1(n_698), .A2(n_716), .B(n_719), .Y(n_857) );
A2O1A1Ixp33_ASAP7_75t_L g858 ( .A1(n_759), .A2(n_66), .B(n_67), .C(n_68), .Y(n_858) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_697), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_768), .Y(n_860) );
INVx5_ASAP7_75t_L g861 ( .A(n_705), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_769), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g863 ( .A1(n_714), .A2(n_202), .B(n_200), .Y(n_863) );
AOI21xp5_ASAP7_75t_L g864 ( .A1(n_718), .A2(n_206), .B(n_205), .Y(n_864) );
AOI221xp5_ASAP7_75t_SL g865 ( .A1(n_721), .A2(n_66), .B1(n_67), .B2(n_69), .C(n_70), .Y(n_865) );
OR2x2_ASAP7_75t_L g866 ( .A(n_673), .B(n_69), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_748), .B(n_71), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_778), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_699), .B(n_72), .Y(n_869) );
CKINVDCx11_ASAP7_75t_R g870 ( .A(n_663), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_747), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g872 ( .A(n_691), .B(n_697), .Y(n_872) );
BUFx3_ASAP7_75t_L g873 ( .A(n_705), .Y(n_873) );
AOI221x1_ASAP7_75t_L g874 ( .A1(n_754), .A2(n_739), .B1(n_774), .B2(n_772), .C(n_762), .Y(n_874) );
AND2x4_ASAP7_75t_L g875 ( .A(n_722), .B(n_72), .Y(n_875) );
OAI22x1_ASAP7_75t_L g876 ( .A1(n_726), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_683), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_706), .B(n_76), .Y(n_878) );
CKINVDCx11_ASAP7_75t_R g879 ( .A(n_713), .Y(n_879) );
BUFx2_ASAP7_75t_L g880 ( .A(n_766), .Y(n_880) );
BUFx2_ASAP7_75t_L g881 ( .A(n_713), .Y(n_881) );
BUFx6f_ASAP7_75t_L g882 ( .A(n_667), .Y(n_882) );
BUFx2_ASAP7_75t_R g883 ( .A(n_744), .Y(n_883) );
NOR2x1_ASAP7_75t_SL g884 ( .A(n_667), .B(n_76), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_678), .B(n_78), .Y(n_885) );
BUFx2_ASAP7_75t_L g886 ( .A(n_751), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_686), .B(n_79), .Y(n_887) );
NAND2xp5_ASAP7_75t_SL g888 ( .A(n_702), .B(n_79), .Y(n_888) );
INVxp67_ASAP7_75t_SL g889 ( .A(n_703), .Y(n_889) );
AO21x1_ASAP7_75t_L g890 ( .A1(n_782), .A2(n_214), .B(n_213), .Y(n_890) );
OR2x2_ASAP7_75t_L g891 ( .A(n_679), .B(n_693), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_750), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_711), .B(n_725), .Y(n_893) );
INVx3_ASAP7_75t_SL g894 ( .A(n_665), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_781), .Y(n_895) );
A2O1A1Ixp33_ASAP7_75t_L g896 ( .A1(n_736), .A2(n_83), .B(n_84), .C(n_85), .Y(n_896) );
OA21x2_ASAP7_75t_L g897 ( .A1(n_739), .A2(n_231), .B(n_304), .Y(n_897) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_684), .A2(n_83), .B1(n_85), .B2(n_86), .Y(n_898) );
INVx6_ASAP7_75t_L g899 ( .A(n_704), .Y(n_899) );
NAND2xp33_ASAP7_75t_L g900 ( .A(n_704), .B(n_215), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_749), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_732), .A2(n_86), .B1(n_87), .B2(n_88), .Y(n_902) );
AOI21xp5_ASAP7_75t_L g903 ( .A1(n_730), .A2(n_238), .B(n_299), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_668), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_741), .Y(n_905) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_724), .A2(n_88), .B1(n_89), .B2(n_90), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_708), .B(n_91), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_704), .Y(n_908) );
AND2x4_ASAP7_75t_L g909 ( .A(n_724), .B(n_92), .Y(n_909) );
A2O1A1Ixp33_ASAP7_75t_L g910 ( .A1(n_692), .A2(n_92), .B(n_93), .C(n_95), .Y(n_910) );
AO21x1_ASAP7_75t_L g911 ( .A1(n_702), .A2(n_242), .B(n_298), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g912 ( .A1(n_707), .A2(n_95), .B1(n_96), .B2(n_97), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_729), .B(n_96), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g914 ( .A(n_729), .B(n_97), .Y(n_914) );
INVxp67_ASAP7_75t_L g915 ( .A(n_771), .Y(n_915) );
OR2x6_ASAP7_75t_L g916 ( .A(n_690), .B(n_99), .Y(n_916) );
NAND2xp5_ASAP7_75t_SL g917 ( .A(n_777), .B(n_99), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_676), .Y(n_918) );
AOI21xp5_ASAP7_75t_L g919 ( .A1(n_677), .A2(n_245), .B(n_295), .Y(n_919) );
BUFx8_ASAP7_75t_SL g920 ( .A(n_666), .Y(n_920) );
INVx4_ASAP7_75t_L g921 ( .A(n_690), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_701), .B(n_100), .Y(n_922) );
AOI21xp5_ASAP7_75t_SL g923 ( .A1(n_780), .A2(n_301), .B(n_240), .Y(n_923) );
NOR2xp33_ASAP7_75t_SL g924 ( .A(n_724), .B(n_216), .Y(n_924) );
NAND3x1_ASAP7_75t_L g925 ( .A(n_731), .B(n_102), .C(n_104), .Y(n_925) );
O2A1O1Ixp33_ASAP7_75t_SL g926 ( .A1(n_758), .A2(n_229), .B(n_289), .C(n_287), .Y(n_926) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_701), .B(n_102), .Y(n_927) );
INVx4_ASAP7_75t_SL g928 ( .A(n_690), .Y(n_928) );
OAI21xp5_ASAP7_75t_L g929 ( .A1(n_670), .A2(n_104), .B(n_105), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_676), .Y(n_930) );
BUFx2_ASAP7_75t_SL g931 ( .A(n_690), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_701), .B(n_105), .Y(n_932) );
NAND2xp5_ASAP7_75t_SL g933 ( .A(n_777), .B(n_106), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_676), .B(n_106), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_676), .B(n_107), .Y(n_935) );
OAI21x1_ASAP7_75t_SL g936 ( .A1(n_676), .A2(n_107), .B(n_108), .Y(n_936) );
BUFx5_ASAP7_75t_L g937 ( .A(n_705), .Y(n_937) );
INVx2_ASAP7_75t_L g938 ( .A(n_676), .Y(n_938) );
INVx2_ASAP7_75t_SL g939 ( .A(n_690), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_892), .B(n_108), .Y(n_940) );
BUFx12f_ASAP7_75t_L g941 ( .A(n_845), .Y(n_941) );
AO21x2_ASAP7_75t_L g942 ( .A1(n_801), .A2(n_250), .B(n_285), .Y(n_942) );
OAI21xp5_ASAP7_75t_L g943 ( .A1(n_929), .A2(n_109), .B(n_110), .Y(n_943) );
INVx1_ASAP7_75t_SL g944 ( .A(n_886), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_791), .Y(n_945) );
AO31x2_ASAP7_75t_L g946 ( .A1(n_810), .A2(n_110), .A3(n_112), .B(n_113), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_918), .Y(n_947) );
INVx2_ASAP7_75t_SL g948 ( .A(n_859), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_930), .Y(n_949) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_804), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_901), .B(n_112), .Y(n_951) );
HB1xp67_ASAP7_75t_L g952 ( .A(n_915), .Y(n_952) );
INVx4_ASAP7_75t_L g953 ( .A(n_928), .Y(n_953) );
OR2x2_ASAP7_75t_L g954 ( .A(n_812), .B(n_114), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_891), .B(n_114), .Y(n_955) );
INVx2_ASAP7_75t_L g956 ( .A(n_938), .Y(n_956) );
AOI21xp5_ASAP7_75t_L g957 ( .A1(n_893), .A2(n_253), .B(n_279), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_800), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_851), .B(n_115), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_807), .Y(n_960) );
AOI21x1_ASAP7_75t_L g961 ( .A1(n_919), .A2(n_219), .B(n_278), .Y(n_961) );
AND2x4_ASAP7_75t_L g962 ( .A(n_825), .B(n_115), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_871), .B(n_116), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_808), .Y(n_964) );
OAI21xp5_ASAP7_75t_L g965 ( .A1(n_929), .A2(n_116), .B(n_118), .Y(n_965) );
OA21x2_ASAP7_75t_L g966 ( .A1(n_823), .A2(n_824), .B(n_833), .Y(n_966) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_870), .B(n_118), .Y(n_967) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_881), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_798), .Y(n_969) );
INVx3_ASAP7_75t_L g970 ( .A(n_856), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_795), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_844), .B(n_119), .Y(n_972) );
AO31x2_ASAP7_75t_L g973 ( .A1(n_890), .A2(n_120), .A3(n_121), .B(n_122), .Y(n_973) );
NOR2xp33_ASAP7_75t_L g974 ( .A(n_879), .B(n_120), .Y(n_974) );
NAND3xp33_ASAP7_75t_L g975 ( .A(n_865), .B(n_121), .C(n_124), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_934), .Y(n_976) );
INVx2_ASAP7_75t_L g977 ( .A(n_818), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_935), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_821), .Y(n_979) );
AO21x2_ASAP7_75t_L g980 ( .A1(n_809), .A2(n_267), .B(n_263), .Y(n_980) );
OAI21xp5_ASAP7_75t_L g981 ( .A1(n_828), .A2(n_124), .B(n_125), .Y(n_981) );
HB1xp67_ASAP7_75t_L g982 ( .A(n_916), .Y(n_982) );
AO21x2_ASAP7_75t_L g983 ( .A1(n_788), .A2(n_258), .B(n_257), .Y(n_983) );
A2O1A1Ixp33_ASAP7_75t_L g984 ( .A1(n_819), .A2(n_125), .B(n_126), .C(n_127), .Y(n_984) );
AND2x4_ASAP7_75t_L g985 ( .A(n_855), .B(n_126), .Y(n_985) );
OR2x2_ASAP7_75t_L g986 ( .A(n_803), .B(n_127), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_838), .Y(n_987) );
BUFx8_ASAP7_75t_L g988 ( .A(n_816), .Y(n_988) );
AND2x4_ASAP7_75t_L g989 ( .A(n_862), .B(n_129), .Y(n_989) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_916), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_816), .A2(n_130), .B1(n_131), .B2(n_132), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_839), .A2(n_131), .B1(n_134), .B2(n_135), .Y(n_992) );
AOI21xp5_ASAP7_75t_L g993 ( .A1(n_837), .A2(n_857), .B(n_789), .Y(n_993) );
BUFx3_ASAP7_75t_L g994 ( .A(n_860), .Y(n_994) );
UNKNOWN g995 ( );
AND2x6_ASAP7_75t_L g996 ( .A(n_875), .B(n_136), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_794), .Y(n_997) );
BUFx10_ASAP7_75t_L g998 ( .A(n_916), .Y(n_998) );
CKINVDCx11_ASAP7_75t_R g999 ( .A(n_854), .Y(n_999) );
NOR2xp33_ASAP7_75t_L g1000 ( .A(n_846), .B(n_137), .Y(n_1000) );
AOI21xp5_ASAP7_75t_L g1001 ( .A1(n_926), .A2(n_137), .B(n_138), .Y(n_1001) );
INVx3_ASAP7_75t_SL g1002 ( .A(n_928), .Y(n_1002) );
NAND2x1p5_ASAP7_75t_L g1003 ( .A(n_921), .B(n_856), .Y(n_1003) );
BUFx2_ASAP7_75t_L g1004 ( .A(n_846), .Y(n_1004) );
BUFx6f_ASAP7_75t_L g1005 ( .A(n_882), .Y(n_1005) );
BUFx2_ASAP7_75t_L g1006 ( .A(n_921), .Y(n_1006) );
CKINVDCx5p33_ASAP7_75t_R g1007 ( .A(n_920), .Y(n_1007) );
INVx2_ASAP7_75t_SL g1008 ( .A(n_939), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_878), .B(n_868), .Y(n_1009) );
AO31x2_ASAP7_75t_L g1010 ( .A1(n_836), .A2(n_911), .A3(n_790), .B(n_858), .Y(n_1010) );
INVx3_ASAP7_75t_L g1011 ( .A(n_856), .Y(n_1011) );
NOR2xp33_ASAP7_75t_L g1012 ( .A(n_894), .B(n_872), .Y(n_1012) );
INVx2_ASAP7_75t_L g1013 ( .A(n_877), .Y(n_1013) );
OR2x6_ASAP7_75t_L g1014 ( .A(n_931), .B(n_875), .Y(n_1014) );
OR2x6_ASAP7_75t_L g1015 ( .A(n_820), .B(n_787), .Y(n_1015) );
AOI21xp5_ASAP7_75t_L g1016 ( .A1(n_885), .A2(n_887), .B(n_869), .Y(n_1016) );
AND2x4_ASAP7_75t_L g1017 ( .A(n_822), .B(n_861), .Y(n_1017) );
AO21x2_ASAP7_75t_L g1018 ( .A1(n_828), .A2(n_834), .B(n_853), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_794), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_806), .Y(n_1020) );
AO31x2_ASAP7_75t_L g1021 ( .A1(n_910), .A2(n_813), .A3(n_884), .B(n_914), .Y(n_1021) );
OAI21x1_ASAP7_75t_L g1022 ( .A1(n_908), .A2(n_913), .B(n_903), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_831), .Y(n_1023) );
BUFx2_ASAP7_75t_L g1024 ( .A(n_820), .Y(n_1024) );
OAI21xp5_ASAP7_75t_L g1025 ( .A1(n_811), .A2(n_850), .B(n_842), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_895), .Y(n_1026) );
BUFx8_ASAP7_75t_L g1027 ( .A(n_880), .Y(n_1027) );
AND2x4_ASAP7_75t_L g1028 ( .A(n_822), .B(n_861), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_866), .Y(n_1029) );
AOI21xp5_ASAP7_75t_L g1030 ( .A1(n_852), .A2(n_863), .B(n_864), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_909), .A2(n_912), .B1(n_830), .B2(n_861), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_922), .Y(n_1032) );
AO21x2_ASAP7_75t_L g1033 ( .A1(n_936), .A2(n_912), .B(n_849), .Y(n_1033) );
INVxp67_ASAP7_75t_L g1034 ( .A(n_817), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_932), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_867), .B(n_905), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_792), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_832), .B(n_793), .Y(n_1038) );
OAI21x1_ASAP7_75t_SL g1039 ( .A1(n_840), .A2(n_843), .B(n_797), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_835), .Y(n_1040) );
CKINVDCx11_ASAP7_75t_R g1041 ( .A(n_815), .Y(n_1041) );
HB1xp67_ASAP7_75t_L g1042 ( .A(n_927), .Y(n_1042) );
INVx1_ASAP7_75t_SL g1043 ( .A(n_830), .Y(n_1043) );
AO21x2_ASAP7_75t_L g1044 ( .A1(n_900), .A2(n_896), .B(n_889), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_799), .Y(n_1045) );
AO31x2_ASAP7_75t_L g1046 ( .A1(n_906), .A2(n_898), .A3(n_876), .B(n_805), .Y(n_1046) );
AOI21xp5_ASAP7_75t_L g1047 ( .A1(n_843), .A2(n_826), .B(n_897), .Y(n_1047) );
INVx2_ASAP7_75t_SL g1048 ( .A(n_814), .Y(n_1048) );
INVx3_ASAP7_75t_L g1049 ( .A(n_873), .Y(n_1049) );
INVx8_ASAP7_75t_L g1050 ( .A(n_882), .Y(n_1050) );
AOI21xp5_ASAP7_75t_L g1051 ( .A1(n_924), .A2(n_888), .B(n_923), .Y(n_1051) );
AOI21x1_ASAP7_75t_L g1052 ( .A1(n_907), .A2(n_904), .B(n_917), .Y(n_1052) );
OA21x2_ASAP7_75t_L g1053 ( .A1(n_785), .A2(n_902), .B(n_933), .Y(n_1053) );
NOR2xp33_ASAP7_75t_L g1054 ( .A(n_883), .B(n_847), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_848), .B(n_827), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_841), .B(n_925), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_827), .B(n_848), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_848), .Y(n_1058) );
INVx4_ASAP7_75t_L g1059 ( .A(n_899), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_899), .B(n_937), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_937), .Y(n_1061) );
INVx3_ASAP7_75t_L g1062 ( .A(n_937), .Y(n_1062) );
OAI21xp5_ASAP7_75t_L g1063 ( .A1(n_929), .A2(n_675), .B(n_670), .Y(n_1063) );
AOI21xp5_ASAP7_75t_L g1064 ( .A1(n_786), .A2(n_580), .B(n_670), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_791), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_791), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_791), .Y(n_1067) );
AOI21xp5_ASAP7_75t_L g1068 ( .A1(n_786), .A2(n_580), .B(n_670), .Y(n_1068) );
OA21x2_ASAP7_75t_L g1069 ( .A1(n_796), .A2(n_760), .B(n_802), .Y(n_1069) );
BUFx2_ASAP7_75t_L g1070 ( .A(n_825), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_901), .B(n_572), .Y(n_1071) );
AO31x2_ASAP7_75t_L g1072 ( .A1(n_874), .A2(n_810), .A3(n_776), .B(n_755), .Y(n_1072) );
OAI21xp5_ASAP7_75t_L g1073 ( .A1(n_929), .A2(n_675), .B(n_670), .Y(n_1073) );
BUFx2_ASAP7_75t_L g1074 ( .A(n_825), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_901), .B(n_572), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_791), .Y(n_1076) );
OAI21x1_ASAP7_75t_SL g1077 ( .A1(n_834), .A2(n_840), .B(n_828), .Y(n_1077) );
OR2x2_ASAP7_75t_L g1078 ( .A(n_804), .B(n_661), .Y(n_1078) );
OR2x6_ASAP7_75t_L g1079 ( .A(n_931), .B(n_690), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_791), .Y(n_1080) );
INVx1_ASAP7_75t_SL g1081 ( .A(n_886), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_791), .Y(n_1082) );
OAI21x1_ASAP7_75t_SL g1083 ( .A1(n_834), .A2(n_840), .B(n_828), .Y(n_1083) );
NAND2x1p5_ASAP7_75t_L g1084 ( .A(n_921), .B(n_690), .Y(n_1084) );
INVx2_ASAP7_75t_L g1085 ( .A(n_938), .Y(n_1085) );
AOI21xp5_ASAP7_75t_L g1086 ( .A1(n_786), .A2(n_580), .B(n_670), .Y(n_1086) );
AOI22xp5_ASAP7_75t_L g1087 ( .A1(n_901), .A2(n_594), .B1(n_575), .B2(n_619), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_791), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1058), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1045), .Y(n_1090) );
OAI33xp33_ASAP7_75t_L g1091 ( .A1(n_991), .A2(n_1040), .A3(n_997), .B1(n_1019), .B2(n_1056), .B3(n_1029), .Y(n_1091) );
INVx2_ASAP7_75t_L g1092 ( .A(n_1069), .Y(n_1092) );
INVx3_ASAP7_75t_L g1093 ( .A(n_1050), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1055), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_956), .B(n_1085), .Y(n_1095) );
AO21x2_ASAP7_75t_L g1096 ( .A1(n_1047), .A2(n_993), .B(n_1057), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g1097 ( .A(n_950), .Y(n_1097) );
BUFx3_ASAP7_75t_L g1098 ( .A(n_1006), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_1087), .B(n_1071), .Y(n_1099) );
INVxp67_ASAP7_75t_L g1100 ( .A(n_952), .Y(n_1100) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_1015), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_945), .Y(n_1102) );
INVx3_ASAP7_75t_L g1103 ( .A(n_1050), .Y(n_1103) );
AND2x4_ASAP7_75t_L g1104 ( .A(n_1017), .B(n_1028), .Y(n_1104) );
INVx3_ASAP7_75t_L g1105 ( .A(n_1050), .Y(n_1105) );
OR2x6_ASAP7_75t_L g1106 ( .A(n_1014), .B(n_1015), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_958), .B(n_960), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_947), .Y(n_1108) );
HB1xp67_ASAP7_75t_L g1109 ( .A(n_1015), .Y(n_1109) );
OR2x2_ASAP7_75t_L g1110 ( .A(n_1078), .B(n_1087), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_949), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_964), .B(n_971), .Y(n_1112) );
INVx3_ASAP7_75t_L g1113 ( .A(n_1017), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_969), .B(n_1065), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1066), .Y(n_1115) );
INVx3_ASAP7_75t_L g1116 ( .A(n_1028), .Y(n_1116) );
OR2x6_ASAP7_75t_L g1117 ( .A(n_1014), .B(n_1024), .Y(n_1117) );
INVx3_ASAP7_75t_L g1118 ( .A(n_1005), .Y(n_1118) );
BUFx2_ASAP7_75t_L g1119 ( .A(n_996), .Y(n_1119) );
OR2x6_ASAP7_75t_L g1120 ( .A(n_1014), .B(n_985), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_1054), .A2(n_1042), .B1(n_996), .B2(n_995), .Y(n_1121) );
OR2x2_ASAP7_75t_L g1122 ( .A(n_944), .B(n_1081), .Y(n_1122) );
AO21x2_ASAP7_75t_L g1123 ( .A1(n_1077), .A2(n_1083), .B(n_1039), .Y(n_1123) );
HB1xp67_ASAP7_75t_L g1124 ( .A(n_944), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1067), .Y(n_1125) );
BUFx3_ASAP7_75t_L g1126 ( .A(n_1084), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_996), .A2(n_985), .B1(n_989), .B2(n_982), .Y(n_1127) );
AO21x2_ASAP7_75t_L g1128 ( .A1(n_1063), .A2(n_1073), .B(n_975), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1076), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1080), .Y(n_1130) );
OR2x2_ASAP7_75t_L g1131 ( .A(n_1081), .B(n_951), .Y(n_1131) );
HB1xp67_ASAP7_75t_SL g1132 ( .A(n_988), .Y(n_1132) );
BUFx2_ASAP7_75t_L g1133 ( .A(n_996), .Y(n_1133) );
HB1xp67_ASAP7_75t_L g1134 ( .A(n_1070), .Y(n_1134) );
AO21x2_ASAP7_75t_L g1135 ( .A1(n_1063), .A2(n_1073), .B(n_975), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1082), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1088), .Y(n_1137) );
INVx2_ASAP7_75t_L g1138 ( .A(n_977), .Y(n_1138) );
OR2x2_ASAP7_75t_L g1139 ( .A(n_951), .B(n_955), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g1140 ( .A(n_1074), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_979), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1013), .B(n_1026), .Y(n_1142) );
INVx4_ASAP7_75t_L g1143 ( .A(n_953), .Y(n_1143) );
OR2x2_ASAP7_75t_L g1144 ( .A(n_1075), .B(n_1032), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_987), .B(n_1009), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_989), .Y(n_1146) );
INVx3_ASAP7_75t_L g1147 ( .A(n_1003), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_940), .Y(n_1148) );
INVxp67_ASAP7_75t_SL g1149 ( .A(n_990), .Y(n_1149) );
BUFx2_ASAP7_75t_L g1150 ( .A(n_1043), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1151 ( .A(n_1035), .B(n_940), .Y(n_1151) );
OAI21x1_ASAP7_75t_L g1152 ( .A1(n_1064), .A2(n_1086), .B(n_1068), .Y(n_1152) );
AND2x4_ASAP7_75t_L g1153 ( .A(n_970), .B(n_1011), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_972), .Y(n_1154) );
BUFx3_ASAP7_75t_L g1155 ( .A(n_1079), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_946), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_959), .Y(n_1157) );
OR2x6_ASAP7_75t_L g1158 ( .A(n_1031), .B(n_943), .Y(n_1158) );
AO31x2_ASAP7_75t_L g1159 ( .A1(n_1031), .A2(n_1001), .A3(n_1016), .B(n_1030), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_943), .B(n_965), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_963), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_965), .B(n_1020), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_962), .Y(n_1163) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1072), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_962), .Y(n_1165) );
INVx2_ASAP7_75t_L g1166 ( .A(n_1072), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1023), .B(n_976), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1034), .B(n_978), .Y(n_1168) );
INVxp67_ASAP7_75t_L g1169 ( .A(n_1079), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_954), .Y(n_1170) );
HB1xp67_ASAP7_75t_L g1171 ( .A(n_968), .Y(n_1171) );
BUFx3_ASAP7_75t_L g1172 ( .A(n_1079), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_986), .Y(n_1173) );
AO21x1_ASAP7_75t_SL g1174 ( .A1(n_981), .A2(n_1061), .B(n_1060), .Y(n_1174) );
INVx3_ASAP7_75t_L g1175 ( .A(n_970), .Y(n_1175) );
BUFx2_ASAP7_75t_L g1176 ( .A(n_1043), .Y(n_1176) );
HB1xp67_ASAP7_75t_L g1177 ( .A(n_948), .Y(n_1177) );
HB1xp67_ASAP7_75t_L g1178 ( .A(n_1008), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1037), .B(n_1038), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1046), .B(n_1036), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_981), .B(n_1025), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_946), .Y(n_1182) );
INVx1_ASAP7_75t_SL g1183 ( .A(n_1004), .Y(n_1183) );
INVx3_ASAP7_75t_L g1184 ( .A(n_1011), .Y(n_1184) );
AO21x2_ASAP7_75t_L g1185 ( .A1(n_1018), .A2(n_1025), .B(n_1033), .Y(n_1185) );
AO21x2_ASAP7_75t_L g1186 ( .A1(n_1018), .A2(n_1033), .B(n_942), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1046), .B(n_946), .Y(n_1187) );
HB1xp67_ASAP7_75t_L g1188 ( .A(n_1048), .Y(n_1188) );
AOI21x1_ASAP7_75t_L g1189 ( .A1(n_966), .A2(n_1051), .B(n_961), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1046), .B(n_991), .Y(n_1190) );
OR2x6_ASAP7_75t_L g1191 ( .A(n_953), .B(n_1062), .Y(n_1191) );
INVxp33_ASAP7_75t_L g1192 ( .A(n_999), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_973), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_973), .Y(n_1194) );
AO21x2_ASAP7_75t_L g1195 ( .A1(n_980), .A2(n_1044), .B(n_1022), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_973), .B(n_984), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1052), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1010), .Y(n_1198) );
OR2x6_ASAP7_75t_L g1199 ( .A(n_1049), .B(n_1059), .Y(n_1199) );
BUFx3_ASAP7_75t_L g1200 ( .A(n_1002), .Y(n_1200) );
INVx2_ASAP7_75t_SL g1201 ( .A(n_988), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1010), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_998), .Y(n_1203) );
BUFx2_ASAP7_75t_L g1204 ( .A(n_1098), .Y(n_1204) );
INVx2_ASAP7_75t_L g1205 ( .A(n_1092), .Y(n_1205) );
INVxp67_ASAP7_75t_L g1206 ( .A(n_1098), .Y(n_1206) );
BUFx2_ASAP7_75t_L g1207 ( .A(n_1119), .Y(n_1207) );
INVx2_ASAP7_75t_L g1208 ( .A(n_1092), .Y(n_1208) );
HB1xp67_ASAP7_75t_L g1209 ( .A(n_1097), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1114), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1114), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1111), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1111), .Y(n_1213) );
OR2x2_ASAP7_75t_L g1214 ( .A(n_1094), .B(n_1021), .Y(n_1214) );
BUFx2_ASAP7_75t_L g1215 ( .A(n_1119), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1216 ( .A(n_1180), .B(n_1021), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1167), .B(n_998), .Y(n_1217) );
NAND2xp5_ASAP7_75t_SL g1218 ( .A(n_1133), .B(n_1000), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1167), .B(n_992), .Y(n_1219) );
INVxp67_ASAP7_75t_SL g1220 ( .A(n_1133), .Y(n_1220) );
OR2x2_ASAP7_75t_L g1221 ( .A(n_1180), .B(n_1021), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1110), .B(n_1012), .Y(n_1222) );
AND2x4_ASAP7_75t_L g1223 ( .A(n_1089), .B(n_1059), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1190), .B(n_1010), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1190), .B(n_983), .Y(n_1225) );
BUFx6f_ASAP7_75t_L g1226 ( .A(n_1191), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1187), .B(n_1053), .Y(n_1227) );
HB1xp67_ASAP7_75t_L g1228 ( .A(n_1122), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1110), .B(n_967), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1187), .B(n_1053), .Y(n_1230) );
BUFx2_ASAP7_75t_L g1231 ( .A(n_1120), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1115), .Y(n_1232) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1131), .B(n_994), .Y(n_1233) );
OR2x2_ASAP7_75t_L g1234 ( .A(n_1131), .B(n_974), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1181), .B(n_957), .Y(n_1235) );
CKINVDCx16_ASAP7_75t_R g1236 ( .A(n_1132), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1115), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1181), .B(n_1041), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1239 ( .A(n_1122), .B(n_1007), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g1240 ( .A(n_1124), .Y(n_1240) );
INVx1_ASAP7_75t_SL g1241 ( .A(n_1126), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1144), .B(n_1027), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1125), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1138), .B(n_941), .Y(n_1244) );
INVxp67_ASAP7_75t_SL g1245 ( .A(n_1127), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_1090), .B(n_1027), .Y(n_1246) );
HB1xp67_ASAP7_75t_L g1247 ( .A(n_1134), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1144), .B(n_1099), .Y(n_1248) );
BUFx2_ASAP7_75t_L g1249 ( .A(n_1104), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1107), .B(n_1090), .Y(n_1250) );
INVxp67_ASAP7_75t_L g1251 ( .A(n_1177), .Y(n_1251) );
INVx3_ASAP7_75t_L g1252 ( .A(n_1191), .Y(n_1252) );
OR2x2_ASAP7_75t_L g1253 ( .A(n_1151), .B(n_1139), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1125), .Y(n_1254) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_1121), .A2(n_1158), .B1(n_1160), .B2(n_1091), .Y(n_1255) );
BUFx2_ASAP7_75t_L g1256 ( .A(n_1120), .Y(n_1256) );
INVxp67_ASAP7_75t_SL g1257 ( .A(n_1150), .Y(n_1257) );
HB1xp67_ASAP7_75t_L g1258 ( .A(n_1140), .Y(n_1258) );
INVx2_ASAP7_75t_SL g1259 ( .A(n_1104), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1112), .B(n_1129), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g1261 ( .A1(n_1158), .A2(n_1160), .B1(n_1120), .B2(n_1162), .Y(n_1261) );
INVxp67_ASAP7_75t_L g1262 ( .A(n_1126), .Y(n_1262) );
OR2x2_ASAP7_75t_SL g1263 ( .A(n_1101), .B(n_1109), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1102), .Y(n_1264) );
NAND2x1_ASAP7_75t_L g1265 ( .A(n_1120), .B(n_1106), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1112), .B(n_1095), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1108), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1130), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1136), .Y(n_1269) );
AND2x4_ASAP7_75t_L g1270 ( .A(n_1123), .B(n_1106), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1137), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1095), .B(n_1142), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1142), .B(n_1162), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1145), .B(n_1170), .Y(n_1274) );
BUFx2_ASAP7_75t_L g1275 ( .A(n_1150), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1198), .B(n_1202), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1141), .B(n_1173), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1198), .B(n_1202), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1151), .B(n_1148), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1158), .B(n_1193), .Y(n_1280) );
AND2x4_ASAP7_75t_L g1281 ( .A(n_1123), .B(n_1106), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1158), .B(n_1193), .Y(n_1282) );
AND2x4_ASAP7_75t_L g1283 ( .A(n_1123), .B(n_1106), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1194), .B(n_1128), .Y(n_1284) );
OR2x2_ASAP7_75t_L g1285 ( .A(n_1139), .B(n_1176), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1100), .B(n_1154), .Y(n_1286) );
AND2x4_ASAP7_75t_L g1287 ( .A(n_1104), .B(n_1113), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1194), .B(n_1128), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1128), .B(n_1135), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_1176), .B(n_1149), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1260), .B(n_1171), .Y(n_1291) );
INVx1_ASAP7_75t_SL g1292 ( .A(n_1241), .Y(n_1292) );
BUFx2_ASAP7_75t_SL g1293 ( .A(n_1226), .Y(n_1293) );
INVx2_ASAP7_75t_L g1294 ( .A(n_1205), .Y(n_1294) );
AND2x4_ASAP7_75t_L g1295 ( .A(n_1270), .B(n_1156), .Y(n_1295) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1205), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1260), .B(n_1168), .Y(n_1297) );
OR2x2_ASAP7_75t_L g1298 ( .A(n_1285), .B(n_1182), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1250), .B(n_1146), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1264), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1285), .B(n_1182), .Y(n_1301) );
OR2x2_ASAP7_75t_L g1302 ( .A(n_1228), .B(n_1185), .Y(n_1302) );
NAND2xp67_ASAP7_75t_L g1303 ( .A(n_1238), .B(n_1196), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1224), .B(n_1185), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1305 ( .A(n_1253), .B(n_1185), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_1250), .B(n_1163), .Y(n_1306) );
INVx2_ASAP7_75t_L g1307 ( .A(n_1208), .Y(n_1307) );
AND2x4_ASAP7_75t_L g1308 ( .A(n_1270), .B(n_1197), .Y(n_1308) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1253), .B(n_1164), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1272), .B(n_1165), .Y(n_1310) );
OR2x2_ASAP7_75t_L g1311 ( .A(n_1273), .B(n_1166), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1273), .B(n_1166), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1227), .B(n_1135), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1267), .Y(n_1314) );
HB1xp67_ASAP7_75t_L g1315 ( .A(n_1204), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1227), .B(n_1135), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1230), .B(n_1096), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1230), .B(n_1096), .Y(n_1318) );
AND2x4_ASAP7_75t_SL g1319 ( .A(n_1287), .B(n_1143), .Y(n_1319) );
NAND2xp5_ASAP7_75t_L g1320 ( .A(n_1272), .B(n_1157), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1280), .B(n_1096), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1280), .B(n_1197), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1282), .B(n_1186), .Y(n_1323) );
OAI22xp5_ASAP7_75t_L g1324 ( .A1(n_1261), .A2(n_1117), .B1(n_1155), .B2(n_1172), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1210), .B(n_1179), .Y(n_1325) );
BUFx3_ASAP7_75t_L g1326 ( .A(n_1223), .Y(n_1326) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1268), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1269), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1282), .B(n_1186), .Y(n_1329) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1271), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1284), .B(n_1186), .Y(n_1331) );
OR2x2_ASAP7_75t_L g1332 ( .A(n_1214), .B(n_1159), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1284), .B(n_1196), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1288), .B(n_1174), .Y(n_1334) );
NOR2xp33_ASAP7_75t_L g1335 ( .A(n_1242), .B(n_1183), .Y(n_1335) );
AND2x4_ASAP7_75t_SL g1336 ( .A(n_1287), .B(n_1143), .Y(n_1336) );
AND2x4_ASAP7_75t_SL g1337 ( .A(n_1287), .B(n_1143), .Y(n_1337) );
OR2x2_ASAP7_75t_L g1338 ( .A(n_1214), .B(n_1159), .Y(n_1338) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_1290), .B(n_1275), .Y(n_1339) );
HB1xp67_ASAP7_75t_L g1340 ( .A(n_1209), .Y(n_1340) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1212), .Y(n_1341) );
AND2x4_ASAP7_75t_SL g1342 ( .A(n_1226), .B(n_1117), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1288), .B(n_1174), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1213), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1276), .B(n_1152), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1276), .B(n_1152), .Y(n_1346) );
INVxp67_ASAP7_75t_SL g1347 ( .A(n_1290), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1278), .B(n_1195), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1349 ( .A(n_1275), .B(n_1159), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1225), .B(n_1195), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_1245), .A2(n_1117), .B1(n_1155), .B2(n_1172), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1211), .B(n_1161), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1300), .Y(n_1353) );
HB1xp67_ASAP7_75t_L g1354 ( .A(n_1340), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1333), .B(n_1312), .Y(n_1355) );
OR2x2_ASAP7_75t_L g1356 ( .A(n_1291), .B(n_1240), .Y(n_1356) );
NAND2x1_ASAP7_75t_SL g1357 ( .A(n_1315), .B(n_1238), .Y(n_1357) );
NOR2xp33_ASAP7_75t_L g1358 ( .A(n_1292), .B(n_1229), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1312), .B(n_1247), .Y(n_1359) );
NOR2x1p5_ASAP7_75t_SL g1360 ( .A(n_1349), .B(n_1189), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1333), .B(n_1216), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1304), .B(n_1221), .Y(n_1362) );
INVx2_ASAP7_75t_L g1363 ( .A(n_1294), .Y(n_1363) );
OR2x2_ASAP7_75t_L g1364 ( .A(n_1311), .B(n_1266), .Y(n_1364) );
INVx1_ASAP7_75t_SL g1365 ( .A(n_1319), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g1366 ( .A(n_1347), .B(n_1258), .Y(n_1366) );
OR2x2_ASAP7_75t_L g1367 ( .A(n_1311), .B(n_1233), .Y(n_1367) );
NAND2xp5_ASAP7_75t_L g1368 ( .A(n_1320), .B(n_1248), .Y(n_1368) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1314), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1304), .B(n_1221), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1297), .B(n_1255), .Y(n_1371) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1327), .Y(n_1372) );
INVx1_ASAP7_75t_SL g1373 ( .A(n_1319), .Y(n_1373) );
INVxp67_ASAP7_75t_L g1374 ( .A(n_1339), .Y(n_1374) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1328), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_1335), .A2(n_1222), .B1(n_1234), .B2(n_1233), .Y(n_1376) );
OR2x6_ASAP7_75t_L g1377 ( .A(n_1326), .B(n_1265), .Y(n_1377) );
NAND2x1_ASAP7_75t_L g1378 ( .A(n_1308), .B(n_1207), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1330), .Y(n_1379) );
OR2x2_ASAP7_75t_L g1380 ( .A(n_1339), .B(n_1309), .Y(n_1380) );
AND2x4_ASAP7_75t_L g1381 ( .A(n_1295), .B(n_1281), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1334), .B(n_1257), .Y(n_1382) );
NOR2xp33_ASAP7_75t_L g1383 ( .A(n_1303), .B(n_1234), .Y(n_1383) );
INVxp67_ASAP7_75t_L g1384 ( .A(n_1326), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1334), .B(n_1206), .Y(n_1385) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1341), .Y(n_1386) );
OR2x2_ASAP7_75t_L g1387 ( .A(n_1309), .B(n_1286), .Y(n_1387) );
HB1xp67_ASAP7_75t_L g1388 ( .A(n_1294), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1344), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1352), .Y(n_1390) );
OR2x2_ASAP7_75t_L g1391 ( .A(n_1298), .B(n_1207), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1392 ( .A(n_1306), .B(n_1232), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1313), .B(n_1289), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1299), .B(n_1237), .Y(n_1394) );
INVx2_ASAP7_75t_L g1395 ( .A(n_1296), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1313), .B(n_1289), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1310), .B(n_1243), .Y(n_1397) );
AND2x2_ASAP7_75t_SL g1398 ( .A(n_1336), .B(n_1215), .Y(n_1398) );
OR2x2_ASAP7_75t_L g1399 ( .A(n_1298), .B(n_1215), .Y(n_1399) );
HB1xp67_ASAP7_75t_L g1400 ( .A(n_1296), .Y(n_1400) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1301), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1316), .B(n_1281), .Y(n_1402) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1301), .Y(n_1403) );
OR2x2_ASAP7_75t_L g1404 ( .A(n_1305), .B(n_1279), .Y(n_1404) );
OAI222xp33_ASAP7_75t_L g1405 ( .A1(n_1343), .A2(n_1218), .B1(n_1246), .B2(n_1249), .C1(n_1231), .C2(n_1256), .Y(n_1405) );
HB1xp67_ASAP7_75t_L g1406 ( .A(n_1307), .Y(n_1406) );
INVxp67_ASAP7_75t_L g1407 ( .A(n_1325), .Y(n_1407) );
NAND2xp5_ASAP7_75t_L g1408 ( .A(n_1316), .B(n_1254), .Y(n_1408) );
OR2x2_ASAP7_75t_L g1409 ( .A(n_1305), .B(n_1251), .Y(n_1409) );
NOR2xp33_ASAP7_75t_L g1410 ( .A(n_1407), .B(n_1236), .Y(n_1410) );
NAND2xp5_ASAP7_75t_L g1411 ( .A(n_1401), .B(n_1403), .Y(n_1411) );
INVx2_ASAP7_75t_L g1412 ( .A(n_1363), .Y(n_1412) );
INVx2_ASAP7_75t_L g1413 ( .A(n_1363), .Y(n_1413) );
AND2x4_ASAP7_75t_L g1414 ( .A(n_1381), .B(n_1402), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1354), .Y(n_1415) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1390), .B(n_1331), .Y(n_1416) );
OAI211xp5_ASAP7_75t_L g1417 ( .A1(n_1357), .A2(n_1351), .B(n_1218), .C(n_1169), .Y(n_1417) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1393), .B(n_1331), .Y(n_1418) );
AND2x2_ASAP7_75t_L g1419 ( .A(n_1355), .B(n_1323), .Y(n_1419) );
INVx2_ASAP7_75t_SL g1420 ( .A(n_1398), .Y(n_1420) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1354), .Y(n_1421) );
HB1xp67_ASAP7_75t_L g1422 ( .A(n_1388), .Y(n_1422) );
AND2x4_ASAP7_75t_L g1423 ( .A(n_1381), .B(n_1295), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1355), .B(n_1323), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1353), .Y(n_1425) );
NOR3xp33_ASAP7_75t_L g1426 ( .A(n_1405), .B(n_1239), .C(n_1244), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1393), .B(n_1329), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1396), .B(n_1317), .Y(n_1428) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1369), .Y(n_1429) );
NAND2x1p5_ASAP7_75t_L g1430 ( .A(n_1398), .B(n_1226), .Y(n_1430) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1372), .Y(n_1431) );
INVx1_ASAP7_75t_SL g1432 ( .A(n_1365), .Y(n_1432) );
INVx2_ASAP7_75t_L g1433 ( .A(n_1395), .Y(n_1433) );
INVx2_ASAP7_75t_L g1434 ( .A(n_1395), .Y(n_1434) );
AOI22xp5_ASAP7_75t_L g1435 ( .A1(n_1383), .A2(n_1343), .B1(n_1324), .B2(n_1329), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1396), .B(n_1321), .Y(n_1436) );
HB1xp67_ASAP7_75t_L g1437 ( .A(n_1388), .Y(n_1437) );
NAND2xp5_ASAP7_75t_L g1438 ( .A(n_1362), .B(n_1317), .Y(n_1438) );
AND2x4_ASAP7_75t_L g1439 ( .A(n_1381), .B(n_1402), .Y(n_1439) );
NAND2x1_ASAP7_75t_L g1440 ( .A(n_1377), .B(n_1283), .Y(n_1440) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1400), .Y(n_1441) );
NAND2xp5_ASAP7_75t_L g1442 ( .A(n_1362), .B(n_1318), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1370), .B(n_1318), .Y(n_1443) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1400), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1375), .Y(n_1445) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1379), .Y(n_1446) );
NAND2xp5_ASAP7_75t_L g1447 ( .A(n_1370), .B(n_1348), .Y(n_1447) );
OR2x2_ASAP7_75t_L g1448 ( .A(n_1380), .B(n_1302), .Y(n_1448) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1406), .Y(n_1449) );
OAI22xp33_ASAP7_75t_L g1450 ( .A1(n_1420), .A2(n_1373), .B1(n_1377), .B2(n_1378), .Y(n_1450) );
AOI21xp5_ASAP7_75t_L g1451 ( .A1(n_1440), .A2(n_1377), .B(n_1337), .Y(n_1451) );
HB1xp67_ASAP7_75t_L g1452 ( .A(n_1422), .Y(n_1452) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1415), .Y(n_1453) );
OA21x2_ASAP7_75t_L g1454 ( .A1(n_1435), .A2(n_1384), .B(n_1371), .Y(n_1454) );
AOI22xp33_ASAP7_75t_L g1455 ( .A1(n_1426), .A2(n_1358), .B1(n_1383), .B2(n_1376), .Y(n_1455) );
INVxp67_ASAP7_75t_L g1456 ( .A(n_1437), .Y(n_1456) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1421), .Y(n_1457) );
INVx2_ASAP7_75t_L g1458 ( .A(n_1412), .Y(n_1458) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1448), .Y(n_1459) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1414), .B(n_1359), .Y(n_1460) );
AOI222xp33_ASAP7_75t_L g1461 ( .A1(n_1410), .A2(n_1376), .B1(n_1358), .B2(n_1374), .C1(n_1368), .C2(n_1366), .Y(n_1461) );
NOR2xp33_ASAP7_75t_L g1462 ( .A(n_1432), .B(n_1239), .Y(n_1462) );
AND2x4_ASAP7_75t_L g1463 ( .A(n_1420), .B(n_1385), .Y(n_1463) );
O2A1O1Ixp33_ASAP7_75t_SL g1464 ( .A1(n_1440), .A2(n_1417), .B(n_1201), .C(n_1303), .Y(n_1464) );
AOI321xp33_ASAP7_75t_SL g1465 ( .A1(n_1418), .A2(n_1192), .A3(n_1356), .B1(n_1201), .B2(n_1246), .C(n_1361), .Y(n_1465) );
INVx2_ASAP7_75t_SL g1466 ( .A(n_1414), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1448), .Y(n_1467) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1425), .Y(n_1468) );
AOI221xp5_ASAP7_75t_L g1469 ( .A1(n_1429), .A2(n_1386), .B1(n_1389), .B2(n_1397), .C(n_1392), .Y(n_1469) );
AOI22xp5_ASAP7_75t_L g1470 ( .A1(n_1416), .A2(n_1382), .B1(n_1244), .B2(n_1408), .Y(n_1470) );
OR2x2_ASAP7_75t_L g1471 ( .A(n_1438), .B(n_1387), .Y(n_1471) );
AOI21xp5_ASAP7_75t_L g1472 ( .A1(n_1430), .A2(n_1337), .B(n_1336), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1414), .B(n_1321), .Y(n_1473) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1431), .Y(n_1474) );
OAI21xp5_ASAP7_75t_L g1475 ( .A1(n_1430), .A2(n_1178), .B(n_1262), .Y(n_1475) );
OAI21xp5_ASAP7_75t_L g1476 ( .A1(n_1430), .A2(n_1188), .B(n_1409), .Y(n_1476) );
A2O1A1Ixp33_ASAP7_75t_L g1477 ( .A1(n_1451), .A2(n_1423), .B(n_1439), .C(n_1200), .Y(n_1477) );
AOI221x1_ASAP7_75t_L g1478 ( .A1(n_1462), .A2(n_1445), .B1(n_1446), .B2(n_1449), .C(n_1444), .Y(n_1478) );
XOR2x2_ASAP7_75t_L g1479 ( .A(n_1462), .B(n_1200), .Y(n_1479) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1459), .Y(n_1480) );
AOI21xp5_ASAP7_75t_L g1481 ( .A1(n_1464), .A2(n_1423), .B(n_1439), .Y(n_1481) );
NAND2xp5_ASAP7_75t_L g1482 ( .A(n_1455), .B(n_1419), .Y(n_1482) );
AOI22xp5_ASAP7_75t_L g1483 ( .A1(n_1455), .A2(n_1423), .B1(n_1439), .B2(n_1411), .Y(n_1483) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1467), .Y(n_1484) );
AOI21xp5_ASAP7_75t_L g1485 ( .A1(n_1450), .A2(n_1444), .B(n_1441), .Y(n_1485) );
OAI21xp5_ASAP7_75t_L g1486 ( .A1(n_1450), .A2(n_1217), .B(n_1277), .Y(n_1486) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1468), .Y(n_1487) );
AOI21xp33_ASAP7_75t_L g1488 ( .A1(n_1461), .A2(n_1203), .B(n_1274), .Y(n_1488) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1474), .Y(n_1489) );
OAI21xp33_ASAP7_75t_SL g1490 ( .A1(n_1466), .A2(n_1424), .B(n_1436), .Y(n_1490) );
AOI22xp33_ASAP7_75t_L g1491 ( .A1(n_1463), .A2(n_1283), .B1(n_1231), .B2(n_1256), .Y(n_1491) );
AOI322xp5_ASAP7_75t_L g1492 ( .A1(n_1465), .A2(n_1424), .A3(n_1427), .B1(n_1436), .B2(n_1428), .C1(n_1443), .C2(n_1442), .Y(n_1492) );
OAI21xp33_ASAP7_75t_SL g1493 ( .A1(n_1460), .A2(n_1447), .B(n_1449), .Y(n_1493) );
AOI221xp5_ASAP7_75t_L g1494 ( .A1(n_1469), .A2(n_1441), .B1(n_1394), .B2(n_1364), .C(n_1413), .Y(n_1494) );
OAI322xp33_ASAP7_75t_L g1495 ( .A1(n_1456), .A2(n_1367), .A3(n_1399), .B1(n_1391), .B2(n_1404), .C1(n_1349), .C2(n_1332), .Y(n_1495) );
OAI211xp5_ASAP7_75t_L g1496 ( .A1(n_1472), .A2(n_1219), .B(n_1259), .C(n_1220), .Y(n_1496) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1473), .B(n_1345), .Y(n_1497) );
NOR2x1_ASAP7_75t_L g1498 ( .A(n_1475), .B(n_1476), .Y(n_1498) );
NAND3xp33_ASAP7_75t_SL g1499 ( .A(n_1456), .B(n_1332), .C(n_1338), .Y(n_1499) );
NOR2xp33_ASAP7_75t_L g1500 ( .A(n_1463), .B(n_1412), .Y(n_1500) );
AOI22xp33_ASAP7_75t_L g1501 ( .A1(n_1454), .A2(n_1283), .B1(n_1295), .B2(n_1350), .Y(n_1501) );
OAI221xp5_ASAP7_75t_L g1502 ( .A1(n_1454), .A2(n_1117), .B1(n_1338), .B2(n_1413), .C(n_1433), .Y(n_1502) );
NAND2xp5_ASAP7_75t_L g1503 ( .A(n_1452), .B(n_1433), .Y(n_1503) );
AOI211xp5_ASAP7_75t_SL g1504 ( .A1(n_1470), .A2(n_1252), .B(n_1235), .C(n_1147), .Y(n_1504) );
NOR2xp33_ASAP7_75t_L g1505 ( .A(n_1471), .B(n_1434), .Y(n_1505) );
NAND3xp33_ASAP7_75t_L g1506 ( .A(n_1453), .B(n_1434), .C(n_1302), .Y(n_1506) );
OAI21xp33_ASAP7_75t_L g1507 ( .A1(n_1457), .A2(n_1360), .B(n_1458), .Y(n_1507) );
NOR3xp33_ASAP7_75t_L g1508 ( .A(n_1486), .B(n_1498), .C(n_1496), .Y(n_1508) );
AOI221xp5_ASAP7_75t_L g1509 ( .A1(n_1488), .A2(n_1482), .B1(n_1494), .B2(n_1495), .C(n_1486), .Y(n_1509) );
A2O1A1Ixp33_ASAP7_75t_L g1510 ( .A1(n_1492), .A2(n_1481), .B(n_1490), .C(n_1493), .Y(n_1510) );
AOI211xp5_ASAP7_75t_L g1511 ( .A1(n_1477), .A2(n_1502), .B(n_1507), .C(n_1485), .Y(n_1511) );
NAND4xp25_ASAP7_75t_L g1512 ( .A(n_1504), .B(n_1483), .C(n_1501), .D(n_1478), .Y(n_1512) );
AOI221xp5_ASAP7_75t_L g1513 ( .A1(n_1499), .A2(n_1480), .B1(n_1484), .B2(n_1489), .C(n_1487), .Y(n_1513) );
NOR3xp33_ASAP7_75t_L g1514 ( .A(n_1506), .B(n_1503), .C(n_1147), .Y(n_1514) );
OAI21xp5_ASAP7_75t_SL g1515 ( .A1(n_1491), .A2(n_1500), .B(n_1342), .Y(n_1515) );
OAI211xp5_ASAP7_75t_SL g1516 ( .A1(n_1479), .A2(n_1505), .B(n_1252), .C(n_1147), .Y(n_1516) );
NOR3xp33_ASAP7_75t_L g1517 ( .A(n_1508), .B(n_1093), .C(n_1103), .Y(n_1517) );
NOR3xp33_ASAP7_75t_L g1518 ( .A(n_1510), .B(n_1093), .C(n_1103), .Y(n_1518) );
NOR3xp33_ASAP7_75t_L g1519 ( .A(n_1512), .B(n_1093), .C(n_1103), .Y(n_1519) );
NAND2xp5_ASAP7_75t_L g1520 ( .A(n_1509), .B(n_1497), .Y(n_1520) );
NAND3x1_ASAP7_75t_L g1521 ( .A(n_1513), .B(n_1252), .C(n_1116), .Y(n_1521) );
NOR2xp33_ASAP7_75t_L g1522 ( .A(n_1515), .B(n_1263), .Y(n_1522) );
NOR3xp33_ASAP7_75t_L g1523 ( .A(n_1516), .B(n_1105), .C(n_1175), .Y(n_1523) );
NAND5xp2_ASAP7_75t_L g1524 ( .A(n_1518), .B(n_1511), .C(n_1514), .D(n_1235), .E(n_1346), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1519), .B(n_1322), .Y(n_1525) );
AND2x4_ASAP7_75t_L g1526 ( .A(n_1517), .B(n_1308), .Y(n_1526) );
NOR3xp33_ASAP7_75t_L g1527 ( .A(n_1520), .B(n_1105), .C(n_1175), .Y(n_1527) );
OR2x6_ASAP7_75t_L g1528 ( .A(n_1521), .B(n_1105), .Y(n_1528) );
INVx2_ASAP7_75t_L g1529 ( .A(n_1526), .Y(n_1529) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1527), .Y(n_1530) );
INVx2_ASAP7_75t_L g1531 ( .A(n_1525), .Y(n_1531) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1524), .Y(n_1532) );
BUFx2_ASAP7_75t_SL g1533 ( .A(n_1529), .Y(n_1533) );
OAI22xp5_ASAP7_75t_L g1534 ( .A1(n_1532), .A2(n_1522), .B1(n_1528), .B2(n_1523), .Y(n_1534) );
AOI22xp33_ASAP7_75t_L g1535 ( .A1(n_1533), .A2(n_1530), .B1(n_1531), .B2(n_1223), .Y(n_1535) );
OAI22xp5_ASAP7_75t_L g1536 ( .A1(n_1534), .A2(n_1263), .B1(n_1293), .B2(n_1199), .Y(n_1536) );
AOI21xp5_ASAP7_75t_L g1537 ( .A1(n_1535), .A2(n_1199), .B(n_1153), .Y(n_1537) );
NAND2xp5_ASAP7_75t_L g1538 ( .A(n_1537), .B(n_1536), .Y(n_1538) );
OR2x6_ASAP7_75t_L g1539 ( .A(n_1538), .B(n_1175), .Y(n_1539) );
AOI21xp5_ASAP7_75t_L g1540 ( .A1(n_1539), .A2(n_1184), .B(n_1118), .Y(n_1540) );
endmodule