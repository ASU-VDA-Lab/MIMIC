module fake_netlist_6_687_n_1732 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1732);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1732;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_15),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_12),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_60),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_36),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_48),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_9),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_14),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_91),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_83),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_57),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_127),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_67),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_40),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_119),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_8),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_65),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_64),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_66),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_33),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_44),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_23),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_45),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_75),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_31),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_85),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_2),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_106),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_72),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_6),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_125),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_95),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_146),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_133),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_39),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_41),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_144),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_21),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_108),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_31),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_150),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_14),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_28),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_1),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_112),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_19),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_118),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_105),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_78),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_23),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_104),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_129),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_161),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_70),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_102),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_107),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_131),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_136),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_30),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_15),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_139),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_163),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_79),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_58),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_1),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_49),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_53),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_156),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_73),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_141),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_74),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_117),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_12),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_142),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_30),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_24),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_69),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_55),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_71),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_51),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_77),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_149),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_88),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_4),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_24),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_93),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_33),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_97),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_53),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_22),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_103),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_137),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_43),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_113),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_114),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_47),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_134),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_100),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_86),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_21),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_87),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_96),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_128),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_61),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_48),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_152),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_120),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_5),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_27),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_9),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_140),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_29),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_126),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_147),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_81),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_47),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_92),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_40),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_80),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_68),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_76),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_51),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_143),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_158),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_109),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_99),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_121),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_2),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_16),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_42),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_110),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_7),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_52),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_45),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_39),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_34),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_13),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_46),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_20),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_124),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_43),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_98),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_34),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_49),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_56),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_17),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_82),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_41),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_19),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_28),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_52),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_27),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_123),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_197),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_181),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_282),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_198),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_282),
.Y(n_333)
);

NOR2xp67_ASAP7_75t_L g334 ( 
.A(n_253),
.B(n_0),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_237),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_200),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_203),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_282),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_289),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_287),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_204),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_208),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_212),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_206),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_253),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_289),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_216),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_224),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_289),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_177),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_0),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_293),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_225),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_324),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_253),
.Y(n_358)
);

NAND2xp33_ASAP7_75t_R g359 ( 
.A(n_268),
.B(n_3),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_310),
.Y(n_360)
);

INVxp33_ASAP7_75t_SL g361 ( 
.A(n_167),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_294),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_259),
.B(n_3),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_258),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_235),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_258),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_243),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_167),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_310),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_278),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_226),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_314),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_187),
.B(n_4),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_314),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_227),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_314),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_324),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_314),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_165),
.B(n_5),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_314),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_228),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_238),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_238),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_295),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_295),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_278),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_170),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_230),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_236),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_217),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_242),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_171),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_190),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_213),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_244),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_245),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_247),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_261),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_214),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_265),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_218),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_272),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_169),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_276),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_246),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_327),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_393),
.B(n_270),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_329),
.B(n_270),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_388),
.B(n_217),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_336),
.B(n_268),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_330),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_337),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_370),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_341),
.B(n_221),
.Y(n_422)
);

NOR2x1_ASAP7_75t_L g423 ( 
.A(n_334),
.B(n_268),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_342),
.Y(n_424)
);

NOR2x1_ASAP7_75t_L g425 ( 
.A(n_331),
.B(n_186),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_371),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_343),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_348),
.Y(n_428)
);

AND2x2_ASAP7_75t_SL g429 ( 
.A(n_353),
.B(n_186),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_406),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g431 ( 
.A1(n_345),
.A2(n_222),
.B(n_210),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_333),
.B(n_168),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_333),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_349),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_357),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_388),
.B(n_166),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_338),
.B(n_339),
.Y(n_437)
);

INVx6_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_328),
.Y(n_439)
);

OAI21x1_ASAP7_75t_L g440 ( 
.A1(n_345),
.A2(n_222),
.B(n_210),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_338),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_356),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_373),
.B(n_229),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_346),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_346),
.B(n_168),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_347),
.Y(n_446)
);

OA21x2_ASAP7_75t_L g447 ( 
.A1(n_347),
.A2(n_351),
.B(n_350),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_332),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_350),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_377),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_R g451 ( 
.A(n_366),
.B(n_313),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_351),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_335),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_355),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_390),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_360),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_360),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_352),
.B(n_166),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_363),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_363),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_374),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_369),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_374),
.B(n_172),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_391),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_375),
.B(n_166),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_376),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_376),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_359),
.A2(n_180),
.B1(n_291),
.B2(n_207),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_398),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_399),
.B(n_264),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_378),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_378),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_380),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_382),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_400),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_436),
.B(n_401),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_417),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_429),
.A2(n_438),
.B1(n_412),
.B2(n_423),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_411),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_416),
.B(n_403),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_409),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_409),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_L g488 ( 
.A(n_423),
.B(n_185),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_429),
.A2(n_364),
.B1(n_344),
.B2(n_381),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_429),
.B(n_264),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_411),
.Y(n_491)
);

AO22x2_ASAP7_75t_L g492 ( 
.A1(n_467),
.A2(n_460),
.B1(n_300),
.B2(n_267),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_417),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_422),
.B(n_405),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_438),
.A2(n_361),
.B1(n_358),
.B2(n_308),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_443),
.B(n_407),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_472),
.B(n_267),
.Y(n_497)
);

INVx4_ASAP7_75t_SL g498 ( 
.A(n_438),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_418),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_438),
.B(n_365),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_409),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_438),
.B(n_383),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_420),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_418),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_421),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_412),
.B(n_234),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_432),
.B(n_320),
.Y(n_507)
);

AND2x6_ASAP7_75t_L g508 ( 
.A(n_436),
.B(n_300),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_410),
.B(n_394),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_451),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_414),
.B(n_367),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_421),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_415),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_414),
.A2(n_249),
.B1(n_302),
.B2(n_303),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_415),
.Y(n_515)
);

AND2x6_ASAP7_75t_L g516 ( 
.A(n_425),
.B(n_185),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_432),
.B(n_318),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_447),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_445),
.B(n_173),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_433),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_415),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_426),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_435),
.B(n_392),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_433),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_419),
.B(n_372),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_465),
.A2(n_322),
.B1(n_305),
.B2(n_325),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_431),
.B(n_389),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_447),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_441),
.B(n_179),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_441),
.B(n_192),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_424),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_459),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_456),
.A2(n_211),
.B1(n_260),
.B2(n_257),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_411),
.Y(n_534)
);

AND2x6_ASAP7_75t_L g535 ( 
.A(n_425),
.B(n_185),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_427),
.B(n_340),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_464),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_480),
.B(n_384),
.Y(n_538)
);

AND2x2_ASAP7_75t_SL g539 ( 
.A(n_470),
.B(n_185),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_426),
.Y(n_540)
);

NOR2x1p5_ASAP7_75t_L g541 ( 
.A(n_428),
.B(n_169),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_447),
.A2(n_262),
.B1(n_301),
.B2(n_219),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_435),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_426),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_459),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_434),
.B(n_219),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_447),
.A2(n_219),
.B1(n_326),
.B2(n_408),
.Y(n_547)
);

BUFx10_ASAP7_75t_L g548 ( 
.A(n_442),
.Y(n_548)
);

AND2x6_ASAP7_75t_L g549 ( 
.A(n_413),
.B(n_219),
.Y(n_549)
);

BUFx4f_ASAP7_75t_L g550 ( 
.A(n_459),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_444),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_431),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_480),
.A2(n_219),
.B1(n_326),
.B2(n_408),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_430),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_457),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_440),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_440),
.B(n_404),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_444),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_446),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_446),
.B(n_196),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_457),
.B(n_395),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_450),
.B(n_326),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_466),
.A2(n_354),
.B1(n_362),
.B2(n_292),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_459),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_444),
.Y(n_565)
);

OR2x6_ASAP7_75t_L g566 ( 
.A(n_471),
.B(n_395),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_459),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_411),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_449),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_470),
.B(n_273),
.C(n_239),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_449),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_SL g572 ( 
.A(n_479),
.B(n_164),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_453),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_453),
.B(n_201),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_413),
.B(n_326),
.Y(n_575)
);

NAND3xp33_ASAP7_75t_L g576 ( 
.A(n_455),
.B(n_240),
.C(n_269),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_455),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_458),
.B(n_202),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_461),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_L g580 ( 
.A(n_411),
.B(n_326),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_461),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_462),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_437),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_463),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_439),
.Y(n_585)
);

OAI22xp33_ASAP7_75t_L g586 ( 
.A1(n_464),
.A2(n_232),
.B1(n_233),
.B2(n_309),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_411),
.B(n_205),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_469),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_437),
.B(n_317),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_459),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_468),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_462),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_475),
.A2(n_404),
.B1(n_402),
.B2(n_397),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_475),
.B(n_384),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_462),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_476),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_477),
.B(n_385),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_477),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_473),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_478),
.B(n_220),
.Y(n_600)
);

AND2x6_ASAP7_75t_L g601 ( 
.A(n_478),
.B(n_231),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_468),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_468),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_468),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_452),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_452),
.B(n_209),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_448),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_452),
.A2(n_402),
.B1(n_397),
.B2(n_396),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_473),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_468),
.B(n_241),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_468),
.B(n_174),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_473),
.B(n_250),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_474),
.A2(n_396),
.B1(n_275),
.B2(n_274),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_L g614 ( 
.A(n_474),
.B(n_251),
.Y(n_614)
);

AND2x6_ASAP7_75t_L g615 ( 
.A(n_474),
.B(n_252),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_474),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_474),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_474),
.Y(n_618)
);

BUFx10_ASAP7_75t_L g619 ( 
.A(n_454),
.Y(n_619)
);

BUFx10_ASAP7_75t_L g620 ( 
.A(n_422),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_557),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_523),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_490),
.A2(n_255),
.B1(n_256),
.B2(n_271),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_557),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_507),
.B(n_175),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_583),
.B(n_279),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_483),
.B(n_284),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_583),
.B(n_296),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_485),
.B(n_494),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_527),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_506),
.B(n_175),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_527),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_510),
.B(n_531),
.Y(n_633)
);

NOR2x1p5_ASAP7_75t_L g634 ( 
.A(n_496),
.B(n_182),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_527),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_490),
.A2(n_297),
.B1(n_176),
.B2(n_292),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_557),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_517),
.B(n_176),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_594),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_525),
.B(n_178),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_486),
.Y(n_641)
);

NOR3xp33_ASAP7_75t_L g642 ( 
.A(n_572),
.B(n_195),
.C(n_199),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_594),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_L g644 ( 
.A(n_508),
.B(n_183),
.Y(n_644)
);

INVxp67_ASAP7_75t_SL g645 ( 
.A(n_590),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_550),
.A2(n_304),
.B(n_280),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_531),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_539),
.B(n_183),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_486),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_555),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_481),
.B(n_184),
.Y(n_651)
);

NAND3xp33_ASAP7_75t_L g652 ( 
.A(n_489),
.B(n_248),
.C(n_263),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_561),
.B(n_555),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_487),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_498),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_539),
.B(n_184),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_547),
.B(n_188),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_531),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_519),
.B(n_188),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_597),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_597),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_543),
.B(n_387),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_487),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_518),
.B(n_194),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_538),
.Y(n_665)
);

INVxp67_ASAP7_75t_SL g666 ( 
.A(n_590),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_492),
.A2(n_288),
.B1(n_194),
.B2(n_280),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_503),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_518),
.B(n_277),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_550),
.A2(n_290),
.B(n_277),
.Y(n_670)
);

NOR3xp33_ASAP7_75t_L g671 ( 
.A(n_572),
.B(n_215),
.C(n_312),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_497),
.A2(n_387),
.B(n_386),
.C(n_223),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_501),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_528),
.A2(n_290),
.B(n_286),
.C(n_288),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_589),
.B(n_182),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_620),
.B(n_299),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_528),
.A2(n_299),
.B(n_286),
.C(n_298),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_508),
.B(n_304),
.Y(n_678)
);

O2A1O1Ixp5_ASAP7_75t_L g679 ( 
.A1(n_497),
.A2(n_386),
.B(n_254),
.C(n_298),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_620),
.B(n_254),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_508),
.B(n_321),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_508),
.A2(n_254),
.B1(n_189),
.B2(n_306),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_508),
.B(n_316),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_482),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_508),
.B(n_319),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_537),
.B(n_323),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_493),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_499),
.B(n_504),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_620),
.B(n_323),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_505),
.B(n_311),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_512),
.Y(n_691)
);

BUFx8_ASAP7_75t_L g692 ( 
.A(n_585),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_601),
.A2(n_281),
.B1(n_306),
.B2(n_285),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_513),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_498),
.B(n_552),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_554),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_513),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_552),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_520),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_524),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_570),
.B(n_307),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_511),
.Y(n_702)
);

AND2x6_ASAP7_75t_L g703 ( 
.A(n_556),
.B(n_59),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_502),
.B(n_285),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_546),
.B(n_281),
.Y(n_705)
);

NOR2xp67_ASAP7_75t_L g706 ( 
.A(n_563),
.B(n_509),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_546),
.B(n_193),
.Y(n_707)
);

INVx8_ASAP7_75t_L g708 ( 
.A(n_566),
.Y(n_708)
);

AND2x6_ASAP7_75t_SL g709 ( 
.A(n_536),
.B(n_283),
.Y(n_709)
);

AND2x2_ASAP7_75t_SL g710 ( 
.A(n_488),
.B(n_122),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_SL g711 ( 
.A(n_548),
.B(n_266),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_562),
.B(n_191),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_515),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_562),
.B(n_191),
.Y(n_714)
);

NOR3x1_ASAP7_75t_L g715 ( 
.A(n_533),
.B(n_189),
.C(n_7),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_515),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_559),
.B(n_162),
.Y(n_717)
);

OAI21xp33_ASAP7_75t_L g718 ( 
.A1(n_495),
.A2(n_6),
.B(n_8),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_521),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_569),
.B(n_571),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_566),
.B(n_10),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_511),
.B(n_10),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_521),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_548),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_573),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_577),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_579),
.B(n_159),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_566),
.B(n_11),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_581),
.B(n_157),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_566),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_606),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_584),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_607),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_606),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_522),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_588),
.B(n_596),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_548),
.B(n_11),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_500),
.B(n_16),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_500),
.B(n_17),
.Y(n_739)
);

INVxp67_ASAP7_75t_SL g740 ( 
.A(n_603),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_598),
.B(n_155),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_542),
.B(n_611),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_586),
.B(n_18),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_500),
.B(n_18),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_492),
.A2(n_153),
.B1(n_138),
.B2(n_132),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_500),
.B(n_20),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_492),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_498),
.B(n_111),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_619),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_526),
.B(n_576),
.C(n_514),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_541),
.A2(n_101),
.B1(n_89),
.B2(n_84),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_619),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_619),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_605),
.B(n_22),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_522),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_551),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_608),
.B(n_25),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_556),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_551),
.Y(n_759)
);

INVx8_ASAP7_75t_L g760 ( 
.A(n_601),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_558),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_529),
.B(n_25),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_616),
.B(n_63),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_540),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_617),
.B(n_62),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_534),
.B(n_26),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_601),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_767)
);

BUFx8_ASAP7_75t_L g768 ( 
.A(n_612),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_540),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_613),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_600),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_530),
.B(n_578),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_617),
.B(n_35),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_560),
.B(n_37),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_558),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_574),
.B(n_37),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_603),
.B(n_618),
.Y(n_777)
);

INVxp33_ASAP7_75t_L g778 ( 
.A(n_600),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_742),
.A2(n_575),
.B(n_565),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_653),
.B(n_593),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_621),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_650),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_627),
.A2(n_575),
.B(n_488),
.C(n_610),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_629),
.B(n_602),
.Y(n_784)
);

INVx5_ASAP7_75t_L g785 ( 
.A(n_703),
.Y(n_785)
);

BUFx4f_ASAP7_75t_L g786 ( 
.A(n_708),
.Y(n_786)
);

AOI21x1_ASAP7_75t_L g787 ( 
.A1(n_777),
.A2(n_587),
.B(n_610),
.Y(n_787)
);

AOI21x1_ASAP7_75t_L g788 ( 
.A1(n_664),
.A2(n_587),
.B(n_609),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_630),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_640),
.B(n_564),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_624),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_637),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_632),
.A2(n_564),
.B(n_532),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_632),
.A2(n_564),
.B(n_532),
.Y(n_794)
);

AOI21x1_ASAP7_75t_L g795 ( 
.A1(n_669),
.A2(n_565),
.B(n_609),
.Y(n_795)
);

A2O1A1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_772),
.A2(n_614),
.B(n_534),
.C(n_592),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_772),
.B(n_582),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_710),
.A2(n_553),
.B1(n_599),
.B2(n_595),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_635),
.A2(n_545),
.B(n_532),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_635),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_698),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_710),
.A2(n_592),
.B1(n_599),
.B2(n_595),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_686),
.Y(n_803)
);

NOR2xp67_ASAP7_75t_L g804 ( 
.A(n_647),
.B(n_582),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_625),
.B(n_601),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_637),
.A2(n_544),
.B(n_601),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_645),
.A2(n_545),
.B(n_567),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_622),
.B(n_544),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_666),
.A2(n_567),
.B(n_545),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_696),
.Y(n_810)
);

BUFx12f_ASAP7_75t_L g811 ( 
.A(n_692),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_767),
.A2(n_747),
.B1(n_734),
.B2(n_627),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_740),
.A2(n_567),
.B(n_591),
.Y(n_813)
);

BUFx8_ASAP7_75t_L g814 ( 
.A(n_753),
.Y(n_814)
);

AOI21xp33_ASAP7_75t_L g815 ( 
.A1(n_701),
.A2(n_580),
.B(n_591),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_750),
.A2(n_568),
.B1(n_491),
.B2(n_484),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_684),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_R g818 ( 
.A(n_658),
.B(n_580),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_702),
.B(n_604),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_674),
.A2(n_516),
.B(n_535),
.Y(n_820)
);

OAI21xp33_ASAP7_75t_L g821 ( 
.A1(n_705),
.A2(n_568),
.B(n_491),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_631),
.B(n_491),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_623),
.A2(n_568),
.B1(n_491),
.B2(n_484),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_687),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_631),
.B(n_568),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_677),
.A2(n_535),
.B(n_516),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_639),
.B(n_484),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_641),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_643),
.B(n_484),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_758),
.A2(n_602),
.B(n_516),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_675),
.B(n_38),
.Y(n_831)
);

AOI21xp33_ASAP7_75t_L g832 ( 
.A1(n_701),
.A2(n_38),
.B(n_42),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_648),
.A2(n_656),
.B(n_766),
.C(n_718),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_758),
.A2(n_602),
.B(n_535),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_731),
.A2(n_535),
.B1(n_549),
.B2(n_612),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_SL g836 ( 
.A(n_711),
.B(n_549),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_698),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_662),
.B(n_44),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_689),
.B(n_46),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_672),
.A2(n_549),
.B(n_612),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_660),
.B(n_661),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_760),
.A2(n_549),
.B(n_615),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_649),
.A2(n_615),
.B(n_612),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_733),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_665),
.B(n_612),
.Y(n_845)
);

AO21x1_ASAP7_75t_L g846 ( 
.A1(n_648),
.A2(n_615),
.B(n_50),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_651),
.A2(n_50),
.B1(n_54),
.B2(n_656),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_668),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_651),
.B(n_638),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_676),
.B(n_689),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_676),
.B(n_778),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_691),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_704),
.B(n_680),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_733),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_706),
.B(n_659),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_699),
.B(n_700),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_707),
.A2(n_714),
.B(n_712),
.C(n_774),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_712),
.A2(n_714),
.B(n_774),
.C(n_776),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_725),
.B(n_726),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_732),
.B(n_626),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_SL g861 ( 
.A(n_633),
.B(n_724),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_695),
.A2(n_657),
.B(n_628),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_688),
.B(n_720),
.Y(n_863)
);

BUFx4f_ASAP7_75t_L g864 ( 
.A(n_708),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_736),
.B(n_722),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_771),
.B(n_730),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_649),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_654),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_634),
.B(n_737),
.Y(n_869)
);

OAI22xp33_ASAP7_75t_L g870 ( 
.A1(n_667),
.A2(n_751),
.B1(n_743),
.B2(n_745),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_728),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_654),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_760),
.A2(n_644),
.B(n_655),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_703),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_738),
.A2(n_746),
.B(n_739),
.C(n_744),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_663),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_760),
.A2(n_655),
.B(n_695),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_708),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_673),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_757),
.A2(n_770),
.B(n_762),
.C(n_636),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_SL g881 ( 
.A(n_703),
.B(n_721),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_703),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_678),
.A2(n_681),
.B(n_685),
.Y(n_883)
);

AOI21x1_ASAP7_75t_L g884 ( 
.A1(n_756),
.A2(n_775),
.B(n_761),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_SL g885 ( 
.A1(n_763),
.A2(n_748),
.B(n_729),
.C(n_727),
.Y(n_885)
);

OAI321xp33_ASAP7_75t_L g886 ( 
.A1(n_652),
.A2(n_721),
.A3(n_682),
.B1(n_746),
.B2(n_744),
.C(n_739),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_738),
.A2(n_754),
.B(n_679),
.C(n_690),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_703),
.Y(n_888)
);

O2A1O1Ixp5_ASAP7_75t_L g889 ( 
.A1(n_683),
.A2(n_773),
.B(n_741),
.C(n_717),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_748),
.A2(n_765),
.B(n_759),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_769),
.B(n_716),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_694),
.A2(n_719),
.B(n_764),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_692),
.Y(n_893)
);

OAI21xp33_ASAP7_75t_L g894 ( 
.A1(n_693),
.A2(n_642),
.B(n_671),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_697),
.A2(n_735),
.B(n_764),
.Y(n_895)
);

NAND2x1p5_ASAP7_75t_L g896 ( 
.A(n_763),
.B(n_723),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_646),
.B(n_670),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_697),
.A2(n_735),
.B(n_713),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_769),
.B(n_723),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_755),
.A2(n_754),
.B(n_749),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_749),
.B(n_752),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_715),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_768),
.B(n_752),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_768),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_709),
.Y(n_905)
);

BUFx8_ASAP7_75t_L g906 ( 
.A(n_753),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_698),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_621),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_637),
.Y(n_909)
);

CKINVDCx10_ASAP7_75t_R g910 ( 
.A(n_692),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_698),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_621),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_629),
.B(n_772),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_742),
.A2(n_632),
.B(n_630),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_629),
.B(n_494),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_629),
.B(n_772),
.Y(n_916)
);

AOI21x1_ASAP7_75t_L g917 ( 
.A1(n_777),
.A2(n_490),
.B(n_664),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_742),
.A2(n_632),
.B(n_630),
.Y(n_918)
);

BUFx4f_ASAP7_75t_L g919 ( 
.A(n_708),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_647),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_650),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_742),
.A2(n_632),
.B(n_630),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_629),
.B(n_772),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_629),
.A2(n_772),
.B(n_705),
.C(n_712),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_627),
.A2(n_490),
.B(n_656),
.C(n_648),
.Y(n_925)
);

AO22x1_ASAP7_75t_L g926 ( 
.A1(n_701),
.A2(n_715),
.B1(n_721),
.B2(n_629),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_650),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_629),
.A2(n_772),
.B(n_705),
.C(n_712),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_627),
.A2(n_490),
.B(n_656),
.C(n_648),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_698),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_653),
.B(n_622),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_742),
.A2(n_632),
.B(n_630),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_629),
.B(n_772),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_742),
.A2(n_632),
.B(n_630),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_629),
.B(n_772),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_621),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_686),
.B(n_537),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_629),
.A2(n_772),
.B(n_705),
.C(n_712),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_742),
.A2(n_632),
.B(n_630),
.Y(n_939)
);

AOI21x1_ASAP7_75t_L g940 ( 
.A1(n_777),
.A2(n_490),
.B(n_664),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_702),
.B(n_639),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_627),
.A2(n_539),
.B1(n_629),
.B2(n_490),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_630),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_629),
.B(n_772),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_742),
.A2(n_632),
.B(n_630),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_629),
.B(n_772),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_629),
.B(n_494),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_801),
.Y(n_948)
);

OAI21x1_ASAP7_75t_SL g949 ( 
.A1(n_846),
.A2(n_833),
.B(n_925),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_858),
.A2(n_857),
.B(n_924),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_913),
.B(n_923),
.Y(n_951)
);

BUFx12f_ASAP7_75t_L g952 ( 
.A(n_811),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_883),
.A2(n_897),
.B(n_933),
.Y(n_953)
);

OAI21x1_ASAP7_75t_L g954 ( 
.A1(n_917),
.A2(n_940),
.B(n_914),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_914),
.A2(n_945),
.B(n_890),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_935),
.A2(n_946),
.B(n_944),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_810),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_915),
.A2(n_947),
.B1(n_942),
.B2(n_865),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_854),
.Y(n_959)
);

AO21x1_ASAP7_75t_L g960 ( 
.A1(n_929),
.A2(n_839),
.B(n_870),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_789),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_945),
.A2(n_884),
.B(n_918),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_844),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_863),
.A2(n_797),
.B(n_885),
.Y(n_964)
);

INVx5_ASAP7_75t_L g965 ( 
.A(n_801),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_800),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_850),
.B(n_790),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_922),
.A2(n_934),
.B(n_932),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_939),
.A2(n_787),
.B(n_873),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_931),
.B(n_780),
.Y(n_970)
);

AOI21x1_ASAP7_75t_L g971 ( 
.A1(n_822),
.A2(n_825),
.B(n_784),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_893),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_851),
.B(n_937),
.Y(n_973)
);

INVx5_ASAP7_75t_L g974 ( 
.A(n_801),
.Y(n_974)
);

OAI22x1_ASAP7_75t_L g975 ( 
.A1(n_902),
.A2(n_847),
.B1(n_853),
.B2(n_866),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_849),
.B(n_860),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_837),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_782),
.Y(n_978)
);

AO22x1_ASAP7_75t_L g979 ( 
.A1(n_905),
.A2(n_920),
.B1(n_869),
.B2(n_803),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_805),
.A2(n_813),
.B(n_809),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_871),
.B(n_838),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_808),
.B(n_841),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_841),
.B(n_856),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_785),
.A2(n_875),
.B1(n_812),
.B2(n_874),
.Y(n_984)
);

NAND2x1p5_ASAP7_75t_L g985 ( 
.A(n_785),
.B(n_874),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_941),
.B(n_921),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_SL g987 ( 
.A(n_861),
.B(n_878),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_SL g988 ( 
.A1(n_874),
.A2(n_888),
.B(n_882),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_785),
.B(n_881),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_927),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_862),
.A2(n_802),
.B(n_796),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_817),
.B(n_824),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_SL g993 ( 
.A1(n_882),
.A2(n_888),
.B(n_785),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_807),
.A2(n_830),
.B(n_834),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_779),
.A2(n_889),
.B(n_816),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_848),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_852),
.B(n_941),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_859),
.B(n_855),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_879),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_831),
.B(n_926),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_804),
.B(n_861),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_880),
.A2(n_832),
.B(n_886),
.C(n_894),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_779),
.A2(n_896),
.B(n_806),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_812),
.A2(n_888),
.B1(n_882),
.B2(n_887),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_781),
.B(n_791),
.Y(n_1005)
);

NAND2x1_ASAP7_75t_L g1006 ( 
.A(n_837),
.B(n_907),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_878),
.B(n_908),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_910),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_912),
.B(n_936),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_896),
.A2(n_806),
.B(n_892),
.Y(n_1010)
);

AOI21x1_ASAP7_75t_L g1011 ( 
.A1(n_891),
.A2(n_793),
.B(n_794),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_901),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_943),
.Y(n_1013)
);

O2A1O1Ixp5_ASAP7_75t_L g1014 ( 
.A1(n_815),
.A2(n_900),
.B(n_862),
.C(n_840),
.Y(n_1014)
);

AOI21xp33_ASAP7_75t_L g1015 ( 
.A1(n_886),
.A2(n_881),
.B(n_845),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_895),
.A2(n_898),
.B(n_877),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_814),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_819),
.B(n_827),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_903),
.B(n_829),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_820),
.A2(n_826),
.B(n_799),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_820),
.A2(n_826),
.B(n_840),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_899),
.A2(n_842),
.B(n_823),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_786),
.B(n_864),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_837),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_815),
.A2(n_821),
.B(n_783),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_792),
.B(n_909),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_786),
.B(n_919),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_907),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_899),
.A2(n_823),
.B(n_798),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_SL g1030 ( 
.A1(n_827),
.A2(n_819),
.B(n_836),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_792),
.B(n_909),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_814),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_872),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_907),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_828),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_911),
.B(n_930),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_864),
.B(n_919),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_835),
.A2(n_868),
.B(n_876),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_911),
.A2(n_930),
.B1(n_867),
.B2(n_904),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_SL g1040 ( 
.A1(n_832),
.A2(n_836),
.B(n_911),
.Y(n_1040)
);

AOI21x1_ASAP7_75t_L g1041 ( 
.A1(n_930),
.A2(n_818),
.B(n_906),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_906),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_SL g1043 ( 
.A1(n_924),
.A2(n_938),
.B(n_928),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_858),
.A2(n_857),
.B(n_924),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_795),
.A2(n_788),
.B(n_843),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_913),
.A2(n_916),
.B(n_933),
.C(n_923),
.Y(n_1046)
);

NAND2x1p5_ASAP7_75t_L g1047 ( 
.A(n_785),
.B(n_874),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_801),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_913),
.B(n_916),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_795),
.A2(n_788),
.B(n_843),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_795),
.A2(n_788),
.B(n_843),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_858),
.A2(n_857),
.B(n_924),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_858),
.A2(n_857),
.B(n_924),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_795),
.A2(n_788),
.B(n_843),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_795),
.A2(n_788),
.B(n_843),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_913),
.A2(n_916),
.B(n_933),
.C(n_923),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_810),
.Y(n_1057)
);

AOI21x1_ASAP7_75t_L g1058 ( 
.A1(n_883),
.A2(n_825),
.B(n_822),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_795),
.A2(n_788),
.B(n_843),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_883),
.A2(n_632),
.B(n_630),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_913),
.B(n_916),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_850),
.B(n_653),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_789),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_795),
.A2(n_788),
.B(n_843),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_795),
.A2(n_788),
.B(n_843),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_883),
.A2(n_632),
.B(n_630),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_883),
.A2(n_632),
.B(n_630),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_913),
.B(n_916),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_913),
.B(n_916),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_795),
.A2(n_788),
.B(n_843),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_913),
.B(n_916),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_801),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_913),
.B(n_916),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_913),
.B(n_916),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_795),
.A2(n_788),
.B(n_843),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_883),
.A2(n_632),
.B(n_630),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_795),
.A2(n_788),
.B(n_843),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_913),
.A2(n_916),
.B(n_933),
.C(n_923),
.Y(n_1078)
);

AO21x2_ASAP7_75t_L g1079 ( 
.A1(n_815),
.A2(n_858),
.B(n_883),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_913),
.B(n_916),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_795),
.A2(n_788),
.B(n_843),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_913),
.B(n_916),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_879),
.Y(n_1083)
);

NAND2x1_ASAP7_75t_L g1084 ( 
.A(n_801),
.B(n_630),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_913),
.A2(n_916),
.B(n_933),
.C(n_923),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_957),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_963),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_1057),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1061),
.A2(n_1082),
.B1(n_1049),
.B2(n_1068),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_950),
.A2(n_1052),
.B(n_1044),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_985),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1061),
.B(n_1082),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_996),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_1023),
.B(n_1027),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_980),
.A2(n_1025),
.B(n_1053),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_970),
.B(n_973),
.Y(n_1096)
);

NAND2x1_ASAP7_75t_L g1097 ( 
.A(n_993),
.B(n_988),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_990),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_951),
.A2(n_1069),
.B1(n_1071),
.B2(n_1073),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_1074),
.B(n_1080),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1013),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_985),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_959),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_956),
.B(n_1046),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_978),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1062),
.B(n_981),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1037),
.B(n_1007),
.Y(n_1107)
);

NOR2xp67_ASAP7_75t_L g1108 ( 
.A(n_1019),
.B(n_978),
.Y(n_1108)
);

AOI221x1_ASAP7_75t_L g1109 ( 
.A1(n_1002),
.A2(n_958),
.B1(n_1015),
.B2(n_984),
.C(n_1004),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1000),
.B(n_986),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_L g1111 ( 
.A(n_1002),
.B(n_967),
.C(n_1056),
.Y(n_1111)
);

INVx3_ASAP7_75t_SL g1112 ( 
.A(n_1017),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1046),
.A2(n_1085),
.B1(n_1056),
.B2(n_1078),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_997),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_952),
.Y(n_1115)
);

OA21x2_ASAP7_75t_L g1116 ( 
.A1(n_991),
.A2(n_1014),
.B(n_1020),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_1047),
.Y(n_1117)
);

OR2x6_ASAP7_75t_L g1118 ( 
.A(n_993),
.B(n_988),
.Y(n_1118)
);

BUFx2_ASAP7_75t_SL g1119 ( 
.A(n_965),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1005),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_972),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_960),
.A2(n_1001),
.B1(n_987),
.B2(n_975),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_976),
.B(n_982),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_977),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1060),
.A2(n_1076),
.B(n_1066),
.Y(n_1125)
);

CKINVDCx16_ASAP7_75t_R g1126 ( 
.A(n_952),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_999),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_965),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_983),
.A2(n_992),
.B1(n_1009),
.B2(n_989),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_972),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1033),
.B(n_1018),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_998),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1008),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1035),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_979),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1047),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_1007),
.B(n_1041),
.Y(n_1137)
);

BUFx10_ASAP7_75t_L g1138 ( 
.A(n_1042),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_977),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1012),
.B(n_1007),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_999),
.B(n_1083),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_977),
.Y(n_1142)
);

OR2x2_ASAP7_75t_L g1143 ( 
.A(n_961),
.B(n_966),
.Y(n_1143)
);

BUFx4f_ASAP7_75t_L g1144 ( 
.A(n_1048),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_965),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1048),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_1063),
.B(n_1034),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1031),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_1048),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_948),
.B(n_1028),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1026),
.Y(n_1151)
);

INVx4_ASAP7_75t_L g1152 ( 
.A(n_965),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1017),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1026),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1039),
.A2(n_1032),
.B1(n_1079),
.B2(n_1036),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1032),
.A2(n_1079),
.B1(n_1084),
.B2(n_1034),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_949),
.A2(n_1040),
.B1(n_1038),
.B2(n_1028),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_948),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_948),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_974),
.A2(n_1024),
.B1(n_1048),
.B2(n_1072),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_1024),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1028),
.B(n_1072),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1072),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_SL g1164 ( 
.A(n_974),
.B(n_1072),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_974),
.Y(n_1165)
);

BUFx12f_ASAP7_75t_L g1166 ( 
.A(n_1006),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1067),
.A2(n_994),
.B(n_968),
.Y(n_1167)
);

CKINVDCx11_ASAP7_75t_R g1168 ( 
.A(n_1030),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_1022),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1029),
.A2(n_971),
.B1(n_1021),
.B2(n_1022),
.Y(n_1170)
);

BUFx12f_ASAP7_75t_L g1171 ( 
.A(n_1058),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_955),
.B(n_1003),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_955),
.B(n_1003),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_954),
.B(n_962),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1010),
.Y(n_1175)
);

OAI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1011),
.A2(n_995),
.B1(n_968),
.B2(n_1016),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1016),
.B(n_969),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1045),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1050),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1050),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1051),
.B(n_1054),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1051),
.A2(n_1054),
.B(n_1055),
.C(n_1059),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1081),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_SL g1184 ( 
.A(n_1077),
.B(n_1064),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1070),
.B(n_1075),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1061),
.A2(n_916),
.B1(n_923),
.B2(n_913),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_977),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1061),
.B(n_1082),
.Y(n_1189)
);

INVx6_ASAP7_75t_L g1190 ( 
.A(n_965),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1061),
.A2(n_916),
.B1(n_923),
.B2(n_913),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_973),
.B(n_915),
.Y(n_1192)
);

INVx6_ASAP7_75t_L g1193 ( 
.A(n_965),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_953),
.A2(n_964),
.B(n_1043),
.Y(n_1194)
);

BUFx4_ASAP7_75t_R g1195 ( 
.A(n_987),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1005),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_957),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_957),
.Y(n_1198)
);

AO22x1_ASAP7_75t_L g1199 ( 
.A1(n_1061),
.A2(n_915),
.B1(n_947),
.B2(n_839),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_957),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1061),
.B(n_1082),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_996),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_953),
.A2(n_964),
.B(n_1043),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1005),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1005),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1061),
.B(n_1082),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1061),
.B(n_1082),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1061),
.A2(n_916),
.B1(n_923),
.B2(n_913),
.Y(n_1208)
);

BUFx10_ASAP7_75t_L g1209 ( 
.A(n_1042),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1061),
.B(n_1082),
.Y(n_1210)
);

BUFx12f_ASAP7_75t_L g1211 ( 
.A(n_952),
.Y(n_1211)
);

INVx3_ASAP7_75t_SL g1212 ( 
.A(n_1017),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1005),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1023),
.B(n_1027),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_973),
.B(n_1062),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_970),
.B(n_937),
.Y(n_1216)
);

OR2x6_ASAP7_75t_L g1217 ( 
.A(n_993),
.B(n_988),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1005),
.Y(n_1218)
);

BUFx2_ASAP7_75t_SL g1219 ( 
.A(n_978),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_952),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1090),
.A2(n_1192),
.B1(n_1122),
.B2(n_1089),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1093),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1144),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1143),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_1190),
.Y(n_1225)
);

CKINVDCx14_ASAP7_75t_R g1226 ( 
.A(n_1088),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1089),
.B(n_1099),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1118),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1134),
.Y(n_1229)
);

OAI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1092),
.A2(n_1206),
.B1(n_1189),
.B2(n_1207),
.Y(n_1230)
);

BUFx8_ASAP7_75t_SL g1231 ( 
.A(n_1211),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1118),
.Y(n_1232)
);

AO21x1_ASAP7_75t_SL g1233 ( 
.A1(n_1090),
.A2(n_1104),
.B(n_1157),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1101),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1086),
.Y(n_1235)
);

OAI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1092),
.A2(n_1189),
.B1(n_1210),
.B2(n_1201),
.Y(n_1236)
);

INVx4_ASAP7_75t_L g1237 ( 
.A(n_1190),
.Y(n_1237)
);

BUFx2_ASAP7_75t_R g1238 ( 
.A(n_1112),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1099),
.B(n_1201),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1097),
.B(n_1175),
.Y(n_1240)
);

CKINVDCx11_ASAP7_75t_R g1241 ( 
.A(n_1212),
.Y(n_1241)
);

NAND2x1p5_ASAP7_75t_L g1242 ( 
.A(n_1178),
.B(n_1179),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1147),
.Y(n_1243)
);

CKINVDCx11_ASAP7_75t_R g1244 ( 
.A(n_1126),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1197),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1215),
.A2(n_1096),
.B1(n_1110),
.B2(n_1191),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1193),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1120),
.Y(n_1248)
);

AO21x2_ASAP7_75t_L g1249 ( 
.A1(n_1167),
.A2(n_1176),
.B(n_1203),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1196),
.Y(n_1250)
);

BUFx2_ASAP7_75t_SL g1251 ( 
.A(n_1108),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_1128),
.Y(n_1252)
);

INVxp33_ASAP7_75t_L g1253 ( 
.A(n_1106),
.Y(n_1253)
);

CKINVDCx11_ASAP7_75t_R g1254 ( 
.A(n_1153),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1206),
.B(n_1207),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1135),
.A2(n_1210),
.B1(n_1195),
.B2(n_1208),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1103),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1204),
.Y(n_1258)
);

BUFx10_ASAP7_75t_L g1259 ( 
.A(n_1133),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1205),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1132),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1123),
.B(n_1100),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1197),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1199),
.B(n_1187),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1187),
.A2(n_1208),
.B1(n_1191),
.B2(n_1111),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1118),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1137),
.B(n_1107),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1213),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1216),
.A2(n_1168),
.B1(n_1129),
.B2(n_1113),
.Y(n_1269)
);

AOI222xp33_ASAP7_75t_L g1270 ( 
.A1(n_1218),
.A2(n_1114),
.B1(n_1113),
.B2(n_1129),
.C1(n_1104),
.C2(n_1214),
.Y(n_1270)
);

INVx11_ASAP7_75t_L g1271 ( 
.A(n_1166),
.Y(n_1271)
);

CKINVDCx11_ASAP7_75t_R g1272 ( 
.A(n_1130),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1114),
.A2(n_1140),
.B1(n_1219),
.B2(n_1164),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1131),
.B(n_1094),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1115),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1148),
.B(n_1127),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1202),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1171),
.A2(n_1098),
.B1(n_1214),
.B2(n_1107),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1194),
.A2(n_1203),
.B(n_1125),
.Y(n_1279)
);

INVx6_ASAP7_75t_L g1280 ( 
.A(n_1152),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1200),
.A2(n_1198),
.B1(n_1137),
.B2(n_1202),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1141),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1116),
.B(n_1173),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1151),
.B(n_1154),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1144),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1182),
.A2(n_1185),
.B(n_1186),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1200),
.A2(n_1155),
.B1(n_1156),
.B2(n_1105),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1131),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1172),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1217),
.A2(n_1087),
.B1(n_1164),
.B2(n_1121),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1158),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1138),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1162),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1170),
.A2(n_1138),
.B1(n_1209),
.B2(n_1116),
.Y(n_1294)
);

CKINVDCx14_ASAP7_75t_R g1295 ( 
.A(n_1220),
.Y(n_1295)
);

AOI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1177),
.A2(n_1173),
.B(n_1183),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1159),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1217),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1209),
.A2(n_1217),
.B1(n_1150),
.B2(n_1117),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1091),
.Y(n_1300)
);

INVx3_ASAP7_75t_L g1301 ( 
.A(n_1091),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1181),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1161),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1161),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1119),
.A2(n_1160),
.B1(n_1145),
.B2(n_1102),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1117),
.B(n_1136),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1174),
.A2(n_1160),
.B(n_1136),
.Y(n_1307)
);

AOI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1177),
.A2(n_1169),
.B(n_1145),
.Y(n_1308)
);

INVx5_ASAP7_75t_SL g1309 ( 
.A(n_1124),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1146),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1139),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1184),
.A2(n_1165),
.B(n_1180),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1142),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1146),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1149),
.A2(n_1124),
.B1(n_1163),
.B2(n_1188),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1163),
.B(n_1188),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1126),
.Y(n_1317)
);

OAI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1092),
.A2(n_711),
.B1(n_629),
.B2(n_913),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1090),
.A2(n_711),
.B1(n_850),
.B2(n_839),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1090),
.A2(n_915),
.B1(n_947),
.B2(n_839),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1143),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1143),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_1108),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1090),
.A2(n_915),
.B1(n_947),
.B2(n_839),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1143),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1143),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1089),
.B(n_1099),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1143),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1109),
.A2(n_995),
.B(n_1095),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1109),
.A2(n_995),
.B(n_1095),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1143),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1261),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1289),
.B(n_1302),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1298),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1261),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1227),
.B(n_1327),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1289),
.B(n_1302),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1222),
.Y(n_1338)
);

NAND2x1_ASAP7_75t_L g1339 ( 
.A(n_1228),
.B(n_1232),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1296),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1296),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1298),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1293),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1283),
.Y(n_1344)
);

AO21x1_ASAP7_75t_SL g1345 ( 
.A1(n_1265),
.A2(n_1269),
.B(n_1264),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1262),
.B(n_1255),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1283),
.B(n_1239),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1293),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1257),
.Y(n_1349)
);

INVxp67_ASAP7_75t_L g1350 ( 
.A(n_1277),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1262),
.B(n_1288),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1239),
.B(n_1233),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1228),
.B(n_1232),
.Y(n_1353)
);

INVx4_ASAP7_75t_L g1354 ( 
.A(n_1298),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1274),
.B(n_1230),
.Y(n_1355)
);

INVxp67_ASAP7_75t_SL g1356 ( 
.A(n_1282),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1308),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1253),
.B(n_1226),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1319),
.A2(n_1324),
.B1(n_1320),
.B2(n_1221),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1313),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1286),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1233),
.B(n_1284),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1313),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1284),
.B(n_1276),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1286),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1276),
.B(n_1270),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1312),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1312),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1228),
.B(n_1232),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1312),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1307),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1307),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1245),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1329),
.B(n_1330),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1329),
.B(n_1330),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1236),
.B(n_1318),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1242),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1242),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1253),
.B(n_1246),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1248),
.B(n_1250),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1291),
.B(n_1297),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1287),
.B(n_1279),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1242),
.Y(n_1383)
);

NAND2x1p5_ASAP7_75t_L g1384 ( 
.A(n_1266),
.B(n_1252),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1240),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1266),
.B(n_1224),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1258),
.B(n_1260),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1294),
.A2(n_1229),
.B(n_1268),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1266),
.B(n_1331),
.Y(n_1389)
);

INVx4_ASAP7_75t_L g1390 ( 
.A(n_1280),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1249),
.A2(n_1290),
.B(n_1310),
.Y(n_1391)
);

BUFx4f_ASAP7_75t_L g1392 ( 
.A(n_1223),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1267),
.B(n_1300),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1226),
.B(n_1263),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1256),
.B(n_1328),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1311),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1241),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1234),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1326),
.B(n_1321),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1299),
.A2(n_1314),
.B(n_1243),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_1322),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1344),
.B(n_1325),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1361),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1344),
.B(n_1303),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1344),
.B(n_1304),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1347),
.B(n_1340),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1347),
.B(n_1281),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1340),
.B(n_1323),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1359),
.A2(n_1278),
.B1(n_1267),
.B2(n_1273),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1378),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1341),
.B(n_1251),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1374),
.B(n_1316),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1374),
.B(n_1316),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1375),
.B(n_1352),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1356),
.B(n_1305),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1335),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1375),
.B(n_1267),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1336),
.B(n_1306),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1352),
.B(n_1306),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1355),
.B(n_1301),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1336),
.B(n_1301),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1339),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1357),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1376),
.B(n_1301),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1345),
.A2(n_1244),
.B1(n_1272),
.B2(n_1317),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1345),
.A2(n_1244),
.B1(n_1272),
.B2(n_1317),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1367),
.B(n_1292),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1333),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1337),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1365),
.B(n_1292),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1395),
.A2(n_1238),
.B1(n_1315),
.B2(n_1295),
.Y(n_1431)
);

AOI21xp33_ASAP7_75t_L g1432 ( 
.A1(n_1382),
.A2(n_1225),
.B(n_1247),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1362),
.B(n_1309),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1367),
.B(n_1235),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1362),
.B(n_1309),
.Y(n_1435)
);

NOR2x1_ASAP7_75t_L g1436 ( 
.A(n_1385),
.B(n_1237),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_L g1437 ( 
.A(n_1432),
.B(n_1382),
.C(n_1379),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1402),
.B(n_1338),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1432),
.B(n_1379),
.C(n_1400),
.Y(n_1439)
);

AND4x1_ASAP7_75t_L g1440 ( 
.A(n_1425),
.B(n_1358),
.C(n_1394),
.D(n_1366),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_SL g1441 ( 
.A(n_1425),
.B(n_1353),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_R g1442 ( 
.A(n_1426),
.B(n_1397),
.Y(n_1442)
);

AND2x2_ASAP7_75t_SL g1443 ( 
.A(n_1426),
.B(n_1334),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1402),
.B(n_1401),
.Y(n_1444)
);

AOI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1424),
.A2(n_1350),
.B1(n_1396),
.B2(n_1349),
.C(n_1401),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1431),
.A2(n_1295),
.B1(n_1346),
.B2(n_1373),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1409),
.A2(n_1392),
.B1(n_1366),
.B2(n_1351),
.Y(n_1447)
);

AND2x2_ASAP7_75t_SL g1448 ( 
.A(n_1415),
.B(n_1334),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1431),
.A2(n_1342),
.B1(n_1334),
.B2(n_1354),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1414),
.B(n_1368),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1414),
.B(n_1368),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1424),
.B(n_1235),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1428),
.B(n_1332),
.Y(n_1453)
);

NAND3xp33_ASAP7_75t_L g1454 ( 
.A(n_1420),
.B(n_1400),
.C(n_1389),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1429),
.B(n_1332),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1429),
.B(n_1343),
.Y(n_1456)
);

NAND2xp33_ASAP7_75t_SL g1457 ( 
.A(n_1415),
.B(n_1334),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1404),
.B(n_1348),
.Y(n_1458)
);

NAND3xp33_ASAP7_75t_L g1459 ( 
.A(n_1420),
.B(n_1411),
.C(n_1409),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1414),
.B(n_1370),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1412),
.B(n_1370),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1412),
.B(n_1391),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1412),
.B(n_1391),
.Y(n_1463)
);

NOR3xp33_ASAP7_75t_L g1464 ( 
.A(n_1411),
.B(n_1390),
.C(n_1339),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1404),
.B(n_1405),
.Y(n_1465)
);

AOI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1416),
.A2(n_1396),
.B1(n_1360),
.B2(n_1363),
.C(n_1387),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1413),
.B(n_1391),
.Y(n_1467)
);

OAI221xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1407),
.A2(n_1399),
.B1(n_1389),
.B2(n_1386),
.C(n_1380),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1413),
.B(n_1371),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_1427),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1405),
.B(n_1364),
.Y(n_1471)
);

NAND3xp33_ASAP7_75t_L g1472 ( 
.A(n_1411),
.B(n_1400),
.C(n_1388),
.Y(n_1472)
);

OAI221xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1407),
.A2(n_1399),
.B1(n_1337),
.B2(n_1378),
.C(n_1372),
.Y(n_1473)
);

AOI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1416),
.A2(n_1364),
.B1(n_1381),
.B2(n_1398),
.C(n_1377),
.Y(n_1474)
);

AOI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1405),
.A2(n_1407),
.B1(n_1418),
.B2(n_1430),
.C(n_1421),
.Y(n_1475)
);

OA211x2_ASAP7_75t_L g1476 ( 
.A1(n_1421),
.A2(n_1384),
.B(n_1392),
.C(n_1390),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1423),
.Y(n_1477)
);

OAI21xp33_ASAP7_75t_L g1478 ( 
.A1(n_1434),
.A2(n_1383),
.B(n_1377),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1419),
.A2(n_1369),
.B1(n_1353),
.B2(n_1393),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1462),
.B(n_1406),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1477),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1438),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1464),
.B(n_1422),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1475),
.B(n_1430),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1477),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1443),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1470),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1450),
.B(n_1417),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1462),
.B(n_1406),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_L g1490 ( 
.A(n_1459),
.B(n_1408),
.C(n_1434),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1469),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1469),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1461),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1450),
.B(n_1417),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1451),
.B(n_1417),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1463),
.B(n_1467),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1460),
.B(n_1419),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1461),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1460),
.B(n_1422),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1463),
.B(n_1422),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1467),
.B(n_1406),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1445),
.B(n_1408),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1448),
.B(n_1419),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1444),
.B(n_1427),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1456),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1465),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1457),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1453),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1455),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1448),
.B(n_1410),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1458),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1452),
.B(n_1254),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1454),
.B(n_1422),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1437),
.B(n_1427),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1471),
.B(n_1479),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1472),
.Y(n_1516)
);

NOR2xp67_ASAP7_75t_L g1517 ( 
.A(n_1516),
.B(n_1439),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1500),
.B(n_1443),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1505),
.B(n_1466),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1512),
.B(n_1241),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1491),
.Y(n_1521)
);

NOR2x1_ASAP7_75t_L g1522 ( 
.A(n_1507),
.B(n_1436),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1516),
.B(n_1473),
.Y(n_1523)
);

O2A1O1Ixp5_ASAP7_75t_L g1524 ( 
.A1(n_1516),
.A2(n_1441),
.B(n_1457),
.C(n_1468),
.Y(n_1524)
);

NOR2x1_ASAP7_75t_L g1525 ( 
.A(n_1507),
.B(n_1441),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1500),
.B(n_1410),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1514),
.B(n_1408),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1490),
.B(n_1440),
.C(n_1449),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1481),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1481),
.Y(n_1530)
);

AND2x4_ASAP7_75t_SL g1531 ( 
.A(n_1510),
.B(n_1433),
.Y(n_1531)
);

INVxp67_ASAP7_75t_L g1532 ( 
.A(n_1508),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1485),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_1514),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1505),
.B(n_1474),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1502),
.A2(n_1440),
.B(n_1447),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1485),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1487),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1483),
.B(n_1500),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1500),
.B(n_1410),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1487),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1499),
.B(n_1403),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1492),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1499),
.B(n_1403),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1492),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1499),
.B(n_1486),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1493),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1484),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1493),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1482),
.B(n_1254),
.Y(n_1550)
);

AND4x1_ASAP7_75t_L g1551 ( 
.A(n_1510),
.B(n_1442),
.C(n_1433),
.D(n_1435),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1509),
.B(n_1511),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1498),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1486),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1509),
.B(n_1478),
.Y(n_1555)
);

OAI21xp33_ASAP7_75t_L g1556 ( 
.A1(n_1536),
.A2(n_1528),
.B(n_1523),
.Y(n_1556)
);

NOR2x1_ASAP7_75t_L g1557 ( 
.A(n_1525),
.B(n_1486),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1518),
.B(n_1499),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1529),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1529),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1518),
.B(n_1546),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1546),
.B(n_1513),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1521),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1530),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1554),
.B(n_1513),
.Y(n_1565)
);

OAI21xp33_ASAP7_75t_L g1566 ( 
.A1(n_1523),
.A2(n_1513),
.B(n_1515),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1554),
.B(n_1513),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1551),
.B(n_1483),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1517),
.A2(n_1446),
.B(n_1483),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1530),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1527),
.B(n_1496),
.Y(n_1571)
);

NAND2x1_ASAP7_75t_L g1572 ( 
.A(n_1522),
.B(n_1483),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1519),
.B(n_1515),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1539),
.B(n_1503),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1539),
.B(n_1503),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1533),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1527),
.B(n_1496),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1537),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1539),
.B(n_1497),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1526),
.B(n_1540),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1534),
.B(n_1480),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1538),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1526),
.B(n_1497),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1540),
.B(n_1488),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1532),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1538),
.Y(n_1586)
);

AND2x4_ASAP7_75t_L g1587 ( 
.A(n_1531),
.B(n_1488),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1541),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1541),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1547),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1542),
.B(n_1544),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1547),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1555),
.B(n_1480),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1524),
.B(n_1511),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1552),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1535),
.B(n_1489),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1549),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1531),
.B(n_1494),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1557),
.B(n_1542),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1574),
.B(n_1544),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1556),
.A2(n_1548),
.B1(n_1550),
.B2(n_1476),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1572),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1559),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1561),
.B(n_1521),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1572),
.A2(n_1568),
.B(n_1569),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1561),
.B(n_1549),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1565),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1559),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1596),
.B(n_1553),
.Y(n_1609)
);

INVx4_ASAP7_75t_L g1610 ( 
.A(n_1585),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1588),
.Y(n_1611)
);

OR2x6_ASAP7_75t_L g1612 ( 
.A(n_1565),
.B(n_1390),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1560),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1573),
.B(n_1543),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1594),
.A2(n_1489),
.B1(n_1501),
.B2(n_1506),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1560),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1564),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1574),
.B(n_1553),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1564),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1570),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1566),
.B(n_1595),
.Y(n_1621)
);

NOR2x1_ASAP7_75t_L g1622 ( 
.A(n_1567),
.B(n_1520),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1575),
.B(n_1545),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1567),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1579),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1596),
.B(n_1501),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1570),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1593),
.B(n_1504),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1587),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1576),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1575),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1580),
.B(n_1494),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1593),
.B(n_1504),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1579),
.B(n_1495),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1605),
.A2(n_1578),
.B(n_1576),
.Y(n_1635)
);

OAI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1605),
.A2(n_1562),
.B(n_1578),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1622),
.A2(n_1562),
.B1(n_1580),
.B2(n_1587),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1610),
.B(n_1583),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1610),
.B(n_1583),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1610),
.B(n_1584),
.Y(n_1640)
);

OAI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1621),
.A2(n_1581),
.B1(n_1577),
.B2(n_1571),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1603),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_SL g1643 ( 
.A1(n_1601),
.A2(n_1558),
.B(n_1581),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1608),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1613),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_SL g1646 ( 
.A1(n_1615),
.A2(n_1558),
.B(n_1587),
.Y(n_1646)
);

NAND3xp33_ASAP7_75t_L g1647 ( 
.A(n_1624),
.B(n_1586),
.C(n_1582),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1631),
.A2(n_1598),
.B1(n_1584),
.B2(n_1476),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1607),
.B(n_1591),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1616),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1614),
.B(n_1231),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1607),
.B(n_1591),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1631),
.B(n_1598),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1628),
.B(n_1231),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1611),
.Y(n_1655)
);

OAI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1629),
.A2(n_1577),
.B1(n_1571),
.B2(n_1598),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1629),
.A2(n_1586),
.B1(n_1582),
.B2(n_1589),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1602),
.A2(n_1589),
.B1(n_1592),
.B2(n_1590),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1599),
.B(n_1590),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1628),
.B(n_1275),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_1659),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1653),
.B(n_1625),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1637),
.B(n_1625),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1638),
.B(n_1623),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1639),
.B(n_1623),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1640),
.B(n_1623),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1655),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1655),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1649),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1647),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1636),
.B(n_1600),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1642),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1654),
.B(n_1275),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1660),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1648),
.B(n_1600),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1644),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1658),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1651),
.B(n_1600),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1641),
.A2(n_1599),
.B1(n_1612),
.B2(n_1602),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1652),
.Y(n_1680)
);

NAND4xp25_ASAP7_75t_L g1681 ( 
.A(n_1679),
.B(n_1643),
.C(n_1646),
.D(n_1635),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1678),
.B(n_1641),
.Y(n_1682)
);

OAI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1670),
.A2(n_1656),
.B(n_1611),
.Y(n_1683)
);

NOR3x1_ASAP7_75t_L g1684 ( 
.A(n_1664),
.B(n_1650),
.C(n_1645),
.Y(n_1684)
);

NOR3xp33_ASAP7_75t_L g1685 ( 
.A(n_1674),
.B(n_1657),
.C(n_1630),
.Y(n_1685)
);

OAI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1670),
.A2(n_1612),
.B1(n_1609),
.B2(n_1620),
.C(n_1627),
.Y(n_1686)
);

NOR3xp33_ASAP7_75t_L g1687 ( 
.A(n_1670),
.B(n_1619),
.C(n_1617),
.Y(n_1687)
);

O2A1O1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1677),
.A2(n_1599),
.B(n_1609),
.C(n_1612),
.Y(n_1688)
);

NOR2x1_ASAP7_75t_L g1689 ( 
.A(n_1667),
.B(n_1612),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1661),
.A2(n_1606),
.B1(n_1618),
.B2(n_1604),
.C(n_1592),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1661),
.A2(n_1633),
.B(n_1606),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1667),
.A2(n_1633),
.B(n_1618),
.Y(n_1692)
);

NOR3xp33_ASAP7_75t_L g1693 ( 
.A(n_1681),
.B(n_1673),
.C(n_1680),
.Y(n_1693)
);

NAND3x1_ASAP7_75t_L g1694 ( 
.A(n_1687),
.B(n_1668),
.C(n_1678),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1692),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1683),
.Y(n_1696)
);

NOR3xp33_ASAP7_75t_L g1697 ( 
.A(n_1682),
.B(n_1668),
.C(n_1669),
.Y(n_1697)
);

NAND3xp33_ASAP7_75t_L g1698 ( 
.A(n_1685),
.B(n_1667),
.C(n_1669),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1691),
.B(n_1662),
.Y(n_1699)
);

NAND4xp75_ASAP7_75t_L g1700 ( 
.A(n_1684),
.B(n_1671),
.C(n_1663),
.D(n_1675),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1686),
.B(n_1665),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_SL g1702 ( 
.A(n_1697),
.B(n_1688),
.C(n_1671),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1698),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1694),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1696),
.B(n_1662),
.Y(n_1705)
);

NAND4xp75_ASAP7_75t_L g1706 ( 
.A(n_1695),
.B(n_1689),
.C(n_1690),
.D(n_1663),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_L g1707 ( 
.A(n_1704),
.B(n_1700),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1705),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1703),
.A2(n_1701),
.B1(n_1693),
.B2(n_1675),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1706),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1702),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1704),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1712),
.B(n_1699),
.Y(n_1713)
);

NOR4xp25_ASAP7_75t_L g1714 ( 
.A(n_1711),
.B(n_1676),
.C(n_1672),
.D(n_1666),
.Y(n_1714)
);

AOI211xp5_ASAP7_75t_L g1715 ( 
.A1(n_1710),
.A2(n_1676),
.B(n_1672),
.C(n_1626),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1707),
.B(n_1672),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1709),
.B(n_1604),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1713),
.B(n_1708),
.Y(n_1718)
);

XNOR2x1_ASAP7_75t_L g1719 ( 
.A(n_1717),
.B(n_1259),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1716),
.Y(n_1720)
);

XNOR2xp5_ASAP7_75t_L g1721 ( 
.A(n_1719),
.B(n_1715),
.Y(n_1721)
);

NOR2x1p5_ASAP7_75t_L g1722 ( 
.A(n_1721),
.B(n_1718),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1722),
.Y(n_1723)
);

AO21x2_ASAP7_75t_L g1724 ( 
.A1(n_1722),
.A2(n_1714),
.B(n_1720),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1724),
.A2(n_1626),
.B(n_1597),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1724),
.B(n_1259),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1726),
.A2(n_1723),
.B1(n_1259),
.B2(n_1634),
.Y(n_1727)
);

OR2x6_ASAP7_75t_L g1728 ( 
.A(n_1725),
.B(n_1271),
.Y(n_1728)
);

OAI21x1_ASAP7_75t_L g1729 ( 
.A1(n_1727),
.A2(n_1563),
.B(n_1632),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1729),
.A2(n_1728),
.B1(n_1634),
.B2(n_1597),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1730),
.A2(n_1563),
.B1(n_1634),
.B2(n_1632),
.C(n_1285),
.Y(n_1731)
);

AOI211xp5_ASAP7_75t_L g1732 ( 
.A1(n_1731),
.A2(n_1271),
.B(n_1285),
.C(n_1223),
.Y(n_1732)
);


endmodule