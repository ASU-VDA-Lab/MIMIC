module fake_netlist_1_12654_n_34 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g9 ( .A(n_1), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_2), .Y(n_10) );
NAND2xp5_ASAP7_75t_SL g11 ( .A(n_4), .B(n_0), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_3), .B(n_4), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g13 ( .A(n_6), .B(n_1), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_3), .B(n_1), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
OAI21xp33_ASAP7_75t_L g17 ( .A1(n_10), .A2(n_0), .B(n_2), .Y(n_17) );
OAI21x1_ASAP7_75t_L g18 ( .A1(n_9), .A2(n_0), .B(n_2), .Y(n_18) );
AOI21xp33_ASAP7_75t_L g19 ( .A1(n_10), .A2(n_6), .B(n_7), .Y(n_19) );
OR2x2_ASAP7_75t_L g20 ( .A(n_16), .B(n_7), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_9), .A2(n_8), .B(n_12), .Y(n_21) );
AOI221x1_ASAP7_75t_L g22 ( .A1(n_9), .A2(n_8), .B1(n_16), .B2(n_15), .C(n_14), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_18), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_20), .B(n_14), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_18), .Y(n_25) );
INVx2_ASAP7_75t_SL g26 ( .A(n_23), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
AOI221x1_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_17), .B1(n_21), .B2(n_19), .C(n_13), .Y(n_28) );
AOI221xp5_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_24), .B1(n_20), .B2(n_11), .C(n_15), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
NOR3xp33_ASAP7_75t_L g31 ( .A(n_29), .B(n_27), .C(n_26), .Y(n_31) );
OAI22xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_22), .B1(n_26), .B2(n_30), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_30), .B(n_26), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_32), .B(n_33), .Y(n_34) );
endmodule