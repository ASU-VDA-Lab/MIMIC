module fake_aes_11193_n_1312 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_356, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_355, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1312);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_355;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1312;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_411;
wire n_860;
wire n_1208;
wire n_1201;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1205;
wire n_923;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_994;
wire n_930;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_1062;
wire n_1271;
wire n_708;
wire n_907;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_1299;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1130;
wire n_584;
wire n_1042;
wire n_912;
wire n_1043;
wire n_1283;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_401;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1275;
wire n_955;
wire n_1093;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_275), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_270), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_26), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_290), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_31), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_192), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_235), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_225), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_352), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_296), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_311), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_349), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_228), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_37), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_76), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_284), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_114), .Y(n_375) );
INVxp33_ASAP7_75t_L g376 ( .A(n_149), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_102), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_339), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_122), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_133), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_16), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_351), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_334), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_158), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_0), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_315), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_268), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_244), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_306), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_3), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_251), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_347), .Y(n_392) );
CKINVDCx16_ASAP7_75t_R g393 ( .A(n_61), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_137), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_229), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_317), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_92), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_285), .Y(n_398) );
INVx2_ASAP7_75t_SL g399 ( .A(n_341), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_278), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_15), .Y(n_401) );
NOR2xp67_ASAP7_75t_L g402 ( .A(n_274), .B(n_118), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_32), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_71), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_280), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_345), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_17), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_22), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_291), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_241), .Y(n_410) );
INVxp33_ASAP7_75t_L g411 ( .A(n_245), .Y(n_411) );
BUFx8_ASAP7_75t_SL g412 ( .A(n_95), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_354), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_226), .Y(n_414) );
CKINVDCx14_ASAP7_75t_R g415 ( .A(n_106), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_353), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_346), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_292), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_338), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_30), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_128), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_282), .Y(n_422) );
BUFx10_ASAP7_75t_L g423 ( .A(n_82), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_7), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_86), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_131), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_44), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_37), .Y(n_428) );
INVxp33_ASAP7_75t_SL g429 ( .A(n_329), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_227), .Y(n_430) );
NOR2xp67_ASAP7_75t_L g431 ( .A(n_243), .B(n_257), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_10), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_115), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_259), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_276), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_117), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_90), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_304), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_97), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_2), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_211), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_233), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_113), .Y(n_443) );
NOR2xp67_ASAP7_75t_L g444 ( .A(n_12), .B(n_121), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_6), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_336), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_252), .Y(n_447) );
BUFx3_ASAP7_75t_L g448 ( .A(n_221), .Y(n_448) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_318), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_298), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_11), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_101), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_325), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_283), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_273), .Y(n_455) );
INVxp33_ASAP7_75t_SL g456 ( .A(n_24), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_335), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_147), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_342), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_288), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_189), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_302), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_156), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_134), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_301), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_332), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_344), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_232), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_9), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_289), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_89), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_55), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_159), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_355), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_72), .Y(n_475) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_56), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_79), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_168), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_320), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_333), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_21), .Y(n_481) );
NOR2xp67_ASAP7_75t_L g482 ( .A(n_17), .B(n_129), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_33), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_126), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_340), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_150), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_194), .Y(n_487) );
BUFx3_ASAP7_75t_L g488 ( .A(n_21), .Y(n_488) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_209), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_269), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_294), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_357), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_271), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_94), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_350), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_312), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_161), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_63), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_224), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_116), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_157), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_337), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_190), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_127), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_356), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_78), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_34), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_255), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_246), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_253), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_203), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_53), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_348), .Y(n_513) );
INVx2_ASAP7_75t_SL g514 ( .A(n_43), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_50), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_167), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_70), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_343), .Y(n_518) );
BUFx5_ASAP7_75t_L g519 ( .A(n_146), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_439), .B(n_0), .Y(n_520) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_366), .A2(n_46), .B(n_45), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_519), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_391), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_519), .Y(n_524) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_449), .Y(n_525) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_363), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_514), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_370), .B(n_1), .Y(n_528) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_449), .Y(n_529) );
BUFx3_ASAP7_75t_L g530 ( .A(n_389), .Y(n_530) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_449), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_399), .B(n_1), .Y(n_532) );
INVx5_ASAP7_75t_L g533 ( .A(n_465), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_372), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_465), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_363), .Y(n_536) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_367), .A2(n_48), .B(n_47), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_427), .B(n_2), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_382), .B(n_3), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_393), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_540) );
BUFx2_ASAP7_75t_L g541 ( .A(n_488), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_423), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_519), .Y(n_543) );
INVx3_ASAP7_75t_L g544 ( .A(n_423), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_376), .B(n_4), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_381), .Y(n_546) );
CKINVDCx6p67_ASAP7_75t_R g547 ( .A(n_458), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_538), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_538), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_542), .B(n_411), .Y(n_550) );
OR2x6_ASAP7_75t_L g551 ( .A(n_520), .B(n_424), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_530), .B(n_404), .Y(n_552) );
INVxp33_ASAP7_75t_L g553 ( .A(n_526), .Y(n_553) );
AND2x6_ASAP7_75t_L g554 ( .A(n_520), .B(n_368), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_536), .B(n_547), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_522), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_542), .B(n_360), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_522), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_524), .Y(n_559) );
BUFx4f_ASAP7_75t_L g560 ( .A(n_547), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_538), .Y(n_561) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_525), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_530), .B(n_471), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_527), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_542), .B(n_362), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_524), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_534), .B(n_377), .Y(n_567) );
AND3x2_ASAP7_75t_L g568 ( .A(n_520), .B(n_489), .C(n_374), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_546), .B(n_378), .Y(n_569) );
NAND2x1p5_ASAP7_75t_L g570 ( .A(n_544), .B(n_440), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_543), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_554), .B(n_523), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_564), .Y(n_573) );
BUFx5_ASAP7_75t_L g574 ( .A(n_554), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_553), .A2(n_545), .B1(n_456), .B2(n_540), .C(n_541), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_570), .B(n_528), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_554), .B(n_544), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_554), .B(n_544), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_551), .B(n_528), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_551), .B(n_528), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_551), .B(n_545), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_560), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_548), .B(n_532), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_555), .A2(n_388), .B1(n_466), .B2(n_359), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_552), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_549), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_552), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_556), .Y(n_588) );
BUFx3_ASAP7_75t_L g589 ( .A(n_560), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_561), .B(n_539), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_550), .A2(n_518), .B1(n_385), .B2(n_401), .Y(n_591) );
OR2x6_ASAP7_75t_L g592 ( .A(n_567), .B(n_451), .Y(n_592) );
INVxp67_ASAP7_75t_L g593 ( .A(n_563), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_558), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_567), .B(n_361), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_569), .A2(n_543), .B1(n_507), .B2(n_429), .Y(n_596) );
AND2x2_ASAP7_75t_SL g597 ( .A(n_569), .B(n_537), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_568), .B(n_415), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_557), .B(n_468), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_563), .B(n_364), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_565), .B(n_365), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_559), .B(n_369), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_566), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_571), .A2(n_537), .B(n_521), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_562), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_562), .B(n_403), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_562), .B(n_371), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_560), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_556), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_570), .B(n_373), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g611 ( .A1(n_583), .A2(n_489), .B(n_374), .C(n_432), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_585), .B(n_407), .Y(n_612) );
NOR2x1p5_ASAP7_75t_L g613 ( .A(n_589), .B(n_408), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_588), .Y(n_614) );
NAND2x1_ASAP7_75t_L g615 ( .A(n_594), .B(n_603), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_581), .B(n_420), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_585), .B(n_428), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_593), .A2(n_481), .B1(n_483), .B2(n_445), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_576), .A2(n_537), .B(n_521), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_579), .A2(n_521), .B(n_380), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_580), .A2(n_392), .B(n_379), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_609), .Y(n_622) );
AOI21x1_ASAP7_75t_L g623 ( .A1(n_604), .A2(n_431), .B(n_402), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_593), .A2(n_396), .B1(n_398), .B2(n_394), .Y(n_624) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_598), .A2(n_383), .B(n_375), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_595), .B(n_412), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_587), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_587), .B(n_384), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_591), .B(n_386), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_604), .A2(n_421), .B(n_418), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_592), .A2(n_430), .B1(n_433), .B2(n_426), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_574), .B(n_387), .Y(n_632) );
AND2x4_ASAP7_75t_L g633 ( .A(n_592), .B(n_444), .Y(n_633) );
BUFx12f_ASAP7_75t_L g634 ( .A(n_582), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_592), .B(n_395), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g636 ( .A1(n_586), .A2(n_482), .B(n_442), .C(n_452), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_590), .A2(n_454), .B(n_450), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_572), .A2(n_459), .B(n_455), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_597), .A2(n_461), .B(n_460), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_597), .A2(n_578), .B(n_577), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_600), .A2(n_464), .B(n_463), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_596), .B(n_397), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_573), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_610), .B(n_400), .Y(n_644) );
INVx2_ASAP7_75t_SL g645 ( .A(n_606), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_602), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_607), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_574), .B(n_405), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_601), .A2(n_478), .B(n_472), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_596), .A2(n_485), .B(n_484), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_584), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_599), .A2(n_491), .B(n_490), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_575), .B(n_406), .Y(n_653) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_605), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_574), .B(n_608), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_574), .B(n_409), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_627), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_640), .A2(n_493), .B(n_492), .Y(n_658) );
AO31x2_ASAP7_75t_L g659 ( .A1(n_620), .A2(n_498), .A3(n_499), .B(n_496), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_643), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_650), .B(n_574), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_619), .A2(n_502), .B(n_500), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_614), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_650), .B(n_612), .Y(n_664) );
OR2x6_ASAP7_75t_L g665 ( .A(n_634), .B(n_613), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_651), .A2(n_616), .B1(n_618), .B2(n_626), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_622), .Y(n_667) );
OAI21x1_ASAP7_75t_L g668 ( .A1(n_623), .A2(n_506), .B(n_505), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_617), .B(n_574), .Y(n_669) );
AND2x4_ASAP7_75t_L g670 ( .A(n_645), .B(n_390), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_646), .B(n_390), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_611), .A2(n_511), .B(n_513), .C(n_509), .Y(n_672) );
AND2x6_ASAP7_75t_L g673 ( .A(n_655), .B(n_516), .Y(n_673) );
OR2x6_ASAP7_75t_L g674 ( .A(n_633), .B(n_390), .Y(n_674) );
OAI21xp5_ASAP7_75t_L g675 ( .A1(n_639), .A2(n_413), .B(n_410), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_647), .B(n_448), .Y(n_676) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_654), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_633), .B(n_469), .Y(n_678) );
INVxp67_ASAP7_75t_L g679 ( .A(n_635), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_637), .A2(n_495), .B(n_474), .C(n_469), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_624), .B(n_469), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_631), .B(n_414), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_628), .B(n_416), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_630), .A2(n_419), .B(n_417), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_653), .A2(n_425), .B1(n_434), .B2(n_422), .Y(n_685) );
AO21x2_ASAP7_75t_L g686 ( .A1(n_636), .A2(n_638), .B(n_641), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_642), .Y(n_687) );
INVx3_ASAP7_75t_L g688 ( .A(n_654), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_652), .A2(n_437), .B1(n_438), .B2(n_436), .C(n_435), .Y(n_689) );
AOI21xp5_ASAP7_75t_SL g690 ( .A1(n_654), .A2(n_476), .B(n_465), .Y(n_690) );
OAI21x1_ASAP7_75t_L g691 ( .A1(n_615), .A2(n_519), .B(n_476), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_629), .Y(n_692) );
AOI31xp67_ASAP7_75t_L g693 ( .A1(n_632), .A2(n_648), .A3(n_519), .B(n_476), .Y(n_693) );
NAND3x1_ASAP7_75t_L g694 ( .A(n_644), .B(n_5), .C(n_7), .Y(n_694) );
OAI21x1_ASAP7_75t_SL g695 ( .A1(n_621), .A2(n_519), .B(n_8), .Y(n_695) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_649), .Y(n_696) );
OAI21x1_ASAP7_75t_L g697 ( .A1(n_656), .A2(n_51), .B(n_49), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_625), .A2(n_443), .B(n_441), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_627), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_643), .Y(n_700) );
AO31x2_ASAP7_75t_L g701 ( .A1(n_620), .A2(n_529), .A3(n_531), .B(n_525), .Y(n_701) );
OAI21x1_ASAP7_75t_L g702 ( .A1(n_619), .A2(n_54), .B(n_52), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_651), .A2(n_447), .B1(n_453), .B2(n_446), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_627), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_627), .B(n_457), .Y(n_705) );
BUFx12f_ASAP7_75t_L g706 ( .A(n_634), .Y(n_706) );
OAI21x1_ASAP7_75t_L g707 ( .A1(n_619), .A2(n_58), .B(n_57), .Y(n_707) );
AOI221x1_ASAP7_75t_L g708 ( .A1(n_620), .A2(n_531), .B1(n_535), .B2(n_529), .C(n_525), .Y(n_708) );
OAI21x1_ASAP7_75t_L g709 ( .A1(n_702), .A2(n_529), .B(n_525), .Y(n_709) );
OA21x2_ASAP7_75t_L g710 ( .A1(n_708), .A2(n_467), .B(n_462), .Y(n_710) );
OAI21x1_ASAP7_75t_L g711 ( .A1(n_707), .A2(n_531), .B(n_529), .Y(n_711) );
OAI21x1_ASAP7_75t_L g712 ( .A1(n_691), .A2(n_535), .B(n_531), .Y(n_712) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_677), .Y(n_713) );
OR2x6_ASAP7_75t_L g714 ( .A(n_706), .B(n_8), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_677), .B(n_664), .Y(n_715) );
OAI21x1_ASAP7_75t_L g716 ( .A1(n_662), .A2(n_535), .B(n_533), .Y(n_716) );
OAI21x1_ASAP7_75t_L g717 ( .A1(n_668), .A2(n_535), .B(n_533), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_660), .Y(n_718) );
AO21x2_ASAP7_75t_L g719 ( .A1(n_695), .A2(n_533), .B(n_60), .Y(n_719) );
OAI21x1_ASAP7_75t_SL g720 ( .A1(n_695), .A2(n_9), .B(n_10), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_669), .A2(n_533), .B(n_473), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_657), .Y(n_722) );
OAI21xp5_ASAP7_75t_L g723 ( .A1(n_672), .A2(n_475), .B(n_470), .Y(n_723) );
AO21x2_ASAP7_75t_L g724 ( .A1(n_658), .A2(n_533), .B(n_62), .Y(n_724) );
OA21x2_ASAP7_75t_L g725 ( .A1(n_697), .A2(n_479), .B(n_477), .Y(n_725) );
OAI21x1_ASAP7_75t_L g726 ( .A1(n_671), .A2(n_64), .B(n_59), .Y(n_726) );
OAI21x1_ASAP7_75t_L g727 ( .A1(n_661), .A2(n_66), .B(n_65), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_686), .A2(n_486), .B(n_480), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_687), .A2(n_494), .B(n_497), .C(n_487), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_700), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_696), .A2(n_503), .B(n_501), .Y(n_731) );
BUFx2_ASAP7_75t_R g732 ( .A(n_705), .Y(n_732) );
OA21x2_ASAP7_75t_L g733 ( .A1(n_680), .A2(n_508), .B(n_504), .Y(n_733) );
OA21x2_ASAP7_75t_L g734 ( .A1(n_701), .A2(n_512), .B(n_510), .Y(n_734) );
BUFx8_ASAP7_75t_L g735 ( .A(n_678), .Y(n_735) );
INVx2_ASAP7_75t_SL g736 ( .A(n_665), .Y(n_736) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_688), .Y(n_737) );
OAI21x1_ASAP7_75t_L g738 ( .A1(n_690), .A2(n_68), .B(n_67), .Y(n_738) );
NAND2xp33_ASAP7_75t_L g739 ( .A(n_673), .B(n_515), .Y(n_739) );
BUFx2_ASAP7_75t_L g740 ( .A(n_674), .Y(n_740) );
OA21x2_ASAP7_75t_L g741 ( .A1(n_701), .A2(n_517), .B(n_73), .Y(n_741) );
BUFx2_ASAP7_75t_L g742 ( .A(n_674), .Y(n_742) );
OAI21x1_ASAP7_75t_L g743 ( .A1(n_667), .A2(n_74), .B(n_69), .Y(n_743) );
BUFx2_ASAP7_75t_L g744 ( .A(n_665), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_663), .Y(n_745) );
AO21x2_ASAP7_75t_L g746 ( .A1(n_675), .A2(n_77), .B(n_75), .Y(n_746) );
INVx3_ASAP7_75t_L g747 ( .A(n_699), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_704), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_659), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_681), .A2(n_11), .B(n_12), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_679), .B(n_13), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_659), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_693), .Y(n_753) );
OAI21xp5_ASAP7_75t_L g754 ( .A1(n_684), .A2(n_13), .B(n_14), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_694), .Y(n_755) );
NAND3xp33_ASAP7_75t_L g756 ( .A(n_666), .B(n_14), .C(n_15), .Y(n_756) );
OAI21x1_ASAP7_75t_L g757 ( .A1(n_683), .A2(n_81), .B(n_80), .Y(n_757) );
NAND2x1_ASAP7_75t_L g758 ( .A(n_673), .B(n_83), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_670), .Y(n_759) );
AOI21x1_ASAP7_75t_L g760 ( .A1(n_676), .A2(n_85), .B(n_84), .Y(n_760) );
AO31x2_ASAP7_75t_L g761 ( .A1(n_682), .A2(n_19), .A3(n_16), .B(n_18), .Y(n_761) );
OAI21x1_ASAP7_75t_L g762 ( .A1(n_698), .A2(n_88), .B(n_87), .Y(n_762) );
AND2x4_ASAP7_75t_L g763 ( .A(n_676), .B(n_18), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_673), .Y(n_764) );
BUFx3_ASAP7_75t_L g765 ( .A(n_692), .Y(n_765) );
OAI21x1_ASAP7_75t_L g766 ( .A1(n_685), .A2(n_93), .B(n_91), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_703), .Y(n_767) );
OR2x2_ASAP7_75t_L g768 ( .A(n_689), .B(n_19), .Y(n_768) );
A2O1A1Ixp33_ASAP7_75t_L g769 ( .A1(n_664), .A2(n_23), .B(n_20), .C(n_22), .Y(n_769) );
OAI21x1_ASAP7_75t_L g770 ( .A1(n_702), .A2(n_98), .B(n_96), .Y(n_770) );
AO31x2_ASAP7_75t_L g771 ( .A1(n_708), .A2(n_24), .A3(n_20), .B(n_23), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_660), .Y(n_772) );
OAI21x1_ASAP7_75t_L g773 ( .A1(n_702), .A2(n_100), .B(n_99), .Y(n_773) );
OR3x4_ASAP7_75t_SL g774 ( .A(n_665), .B(n_25), .C(n_26), .Y(n_774) );
OA21x2_ASAP7_75t_L g775 ( .A1(n_708), .A2(n_104), .B(n_103), .Y(n_775) );
OA21x2_ASAP7_75t_L g776 ( .A1(n_708), .A2(n_107), .B(n_105), .Y(n_776) );
AO21x2_ASAP7_75t_L g777 ( .A1(n_753), .A2(n_25), .B(n_27), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_718), .Y(n_778) );
NAND3x1_ASAP7_75t_L g779 ( .A(n_755), .B(n_27), .C(n_28), .Y(n_779) );
AO21x2_ASAP7_75t_L g780 ( .A1(n_753), .A2(n_28), .B(n_29), .Y(n_780) );
OR2x2_ASAP7_75t_L g781 ( .A(n_722), .B(n_29), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_745), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_755), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_718), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_730), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_772), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_772), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_745), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_744), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_748), .Y(n_790) );
AOI21x1_ASAP7_75t_L g791 ( .A1(n_752), .A2(n_33), .B(n_34), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_747), .Y(n_792) );
OR2x6_ASAP7_75t_L g793 ( .A(n_736), .B(n_35), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_747), .Y(n_794) );
BUFx2_ASAP7_75t_L g795 ( .A(n_735), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_761), .Y(n_796) );
OAI222xp33_ASAP7_75t_L g797 ( .A1(n_714), .A2(n_35), .B1(n_36), .B2(n_38), .C1(n_39), .C2(n_40), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_761), .Y(n_798) );
OA21x2_ASAP7_75t_L g799 ( .A1(n_752), .A2(n_109), .B(n_108), .Y(n_799) );
CKINVDCx6p67_ASAP7_75t_R g800 ( .A(n_714), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_749), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_713), .Y(n_802) );
INVx5_ASAP7_75t_L g803 ( .A(n_713), .Y(n_803) );
INVx4_ASAP7_75t_L g804 ( .A(n_713), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_761), .Y(n_805) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_715), .Y(n_806) );
BUFx2_ASAP7_75t_L g807 ( .A(n_735), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_771), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_771), .Y(n_809) );
INVx3_ASAP7_75t_L g810 ( .A(n_737), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_763), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_767), .B(n_36), .Y(n_812) );
INVx2_ASAP7_75t_SL g813 ( .A(n_765), .Y(n_813) );
OAI21x1_ASAP7_75t_L g814 ( .A1(n_709), .A2(n_111), .B(n_110), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_763), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_751), .Y(n_816) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_764), .Y(n_817) );
AO21x2_ASAP7_75t_L g818 ( .A1(n_711), .A2(n_38), .B(n_39), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_764), .Y(n_819) );
INVx3_ASAP7_75t_L g820 ( .A(n_737), .Y(n_820) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_740), .Y(n_821) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_742), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_768), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_720), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_759), .Y(n_825) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_771), .Y(n_826) );
AOI21x1_ASAP7_75t_L g827 ( .A1(n_741), .A2(n_40), .B(n_41), .Y(n_827) );
INVx2_ASAP7_75t_SL g828 ( .A(n_737), .Y(n_828) );
BUFx2_ASAP7_75t_SL g829 ( .A(n_767), .Y(n_829) );
AOI21x1_ASAP7_75t_L g830 ( .A1(n_741), .A2(n_41), .B(n_42), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_769), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_756), .Y(n_832) );
INVx2_ASAP7_75t_SL g833 ( .A(n_758), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_750), .Y(n_834) );
OAI21x1_ASAP7_75t_L g835 ( .A1(n_712), .A2(n_119), .B(n_112), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_754), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_760), .Y(n_837) );
NOR2x1_ASAP7_75t_L g838 ( .A(n_739), .B(n_42), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_733), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_717), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_733), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_732), .Y(n_842) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_734), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_719), .Y(n_844) );
AO21x2_ASAP7_75t_L g845 ( .A1(n_724), .A2(n_43), .B(n_44), .Y(n_845) );
INVx3_ASAP7_75t_L g846 ( .A(n_766), .Y(n_846) );
AND2x4_ASAP7_75t_L g847 ( .A(n_757), .B(n_120), .Y(n_847) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_734), .Y(n_848) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_725), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_743), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_729), .B(n_123), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_716), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g853 ( .A(n_774), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_746), .A2(n_124), .B1(n_125), .B2(n_130), .Y(n_854) );
OR2x2_ASAP7_75t_L g855 ( .A(n_723), .B(n_132), .Y(n_855) );
AO21x2_ASAP7_75t_L g856 ( .A1(n_724), .A2(n_135), .B(n_136), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_725), .B(n_138), .Y(n_857) );
CKINVDCx8_ASAP7_75t_R g858 ( .A(n_710), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_728), .A2(n_139), .B1(n_140), .B2(n_141), .Y(n_859) );
INVx3_ASAP7_75t_L g860 ( .A(n_762), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_726), .Y(n_861) );
INVx3_ASAP7_75t_L g862 ( .A(n_746), .Y(n_862) );
OAI21xp5_ASAP7_75t_L g863 ( .A1(n_721), .A2(n_142), .B(n_143), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_727), .Y(n_864) );
INVx2_ASAP7_75t_L g865 ( .A(n_738), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_770), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_773), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_710), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_731), .B(n_144), .Y(n_869) );
BUFx2_ASAP7_75t_SL g870 ( .A(n_775), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_775), .B(n_145), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_776), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_776), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_718), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_718), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_722), .B(n_148), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_718), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_718), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_730), .Y(n_879) );
INVx2_ASAP7_75t_SL g880 ( .A(n_795), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_782), .B(n_151), .Y(n_881) );
NAND2xp5_ASAP7_75t_SL g882 ( .A(n_858), .B(n_152), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_816), .B(n_153), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_790), .B(n_154), .Y(n_884) );
AOI221xp5_ASAP7_75t_L g885 ( .A1(n_823), .A2(n_155), .B1(n_160), .B2(n_162), .C(n_163), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_793), .B(n_164), .Y(n_886) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_800), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_782), .B(n_165), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_778), .Y(n_889) );
BUFx2_ASAP7_75t_L g890 ( .A(n_804), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_793), .B(n_166), .Y(n_891) );
OR2x2_ASAP7_75t_L g892 ( .A(n_788), .B(n_358), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_784), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_786), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_787), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_812), .A2(n_169), .B1(n_170), .B2(n_171), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_793), .B(n_172), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_874), .B(n_173), .Y(n_898) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_801), .Y(n_899) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_806), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_785), .B(n_174), .Y(n_901) );
BUFx2_ASAP7_75t_L g902 ( .A(n_804), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_875), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_879), .B(n_175), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_781), .B(n_176), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_878), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_825), .B(n_177), .Y(n_907) );
BUFx2_ASAP7_75t_L g908 ( .A(n_803), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_877), .B(n_178), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_777), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_777), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_811), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_815), .B(n_179), .Y(n_913) );
AND2x2_ASAP7_75t_L g914 ( .A(n_812), .B(n_180), .Y(n_914) );
OR2x2_ASAP7_75t_L g915 ( .A(n_821), .B(n_181), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_829), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_792), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_876), .B(n_182), .Y(n_918) );
OR2x2_ASAP7_75t_L g919 ( .A(n_821), .B(n_183), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_794), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_780), .Y(n_921) );
INVx2_ASAP7_75t_L g922 ( .A(n_780), .Y(n_922) );
NAND2xp5_ASAP7_75t_SL g923 ( .A(n_849), .B(n_184), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_802), .Y(n_924) );
HB1xp67_ASAP7_75t_L g925 ( .A(n_806), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_822), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_822), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_817), .Y(n_928) );
INVx2_ASAP7_75t_L g929 ( .A(n_791), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_836), .B(n_185), .Y(n_930) );
NOR2xp33_ASAP7_75t_L g931 ( .A(n_797), .B(n_186), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_842), .B(n_187), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_817), .Y(n_933) );
AO21x2_ASAP7_75t_L g934 ( .A1(n_837), .A2(n_188), .B(n_191), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_813), .B(n_193), .Y(n_935) );
NOR2xp33_ASAP7_75t_L g936 ( .A(n_797), .B(n_195), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_807), .B(n_196), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_819), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_818), .Y(n_939) );
BUFx2_ASAP7_75t_L g940 ( .A(n_803), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_789), .B(n_197), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_819), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_789), .B(n_198), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_818), .Y(n_944) );
INVx2_ASAP7_75t_L g945 ( .A(n_803), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_834), .B(n_199), .Y(n_946) );
INVx2_ASAP7_75t_L g947 ( .A(n_803), .Y(n_947) );
INVx2_ASAP7_75t_SL g948 ( .A(n_828), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_853), .B(n_200), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_824), .B(n_201), .Y(n_950) );
INVx3_ASAP7_75t_L g951 ( .A(n_810), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_783), .Y(n_952) );
BUFx6f_ASAP7_75t_L g953 ( .A(n_810), .Y(n_953) );
INVx2_ASAP7_75t_SL g954 ( .A(n_820), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_783), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_796), .B(n_202), .Y(n_956) );
AND2x4_ASAP7_75t_L g957 ( .A(n_820), .B(n_204), .Y(n_957) );
HB1xp67_ASAP7_75t_L g958 ( .A(n_849), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_798), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_805), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_853), .B(n_205), .Y(n_961) );
INVx3_ASAP7_75t_L g962 ( .A(n_833), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_839), .Y(n_963) );
AND2x2_ASAP7_75t_L g964 ( .A(n_838), .B(n_206), .Y(n_964) );
INVx2_ASAP7_75t_SL g965 ( .A(n_855), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_831), .B(n_207), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_841), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_826), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_826), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_832), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_843), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_851), .B(n_208), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_845), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_869), .B(n_210), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_857), .B(n_212), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_845), .Y(n_976) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_843), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_848), .B(n_213), .Y(n_978) );
AOI221xp5_ASAP7_75t_L g979 ( .A1(n_859), .A2(n_214), .B1(n_215), .B2(n_216), .C(n_217), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_779), .Y(n_980) );
NOR2x1_ASAP7_75t_SL g981 ( .A(n_859), .B(n_218), .Y(n_981) );
INVx2_ASAP7_75t_L g982 ( .A(n_808), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_848), .B(n_219), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_809), .B(n_220), .Y(n_984) );
AND2x4_ASAP7_75t_L g985 ( .A(n_868), .B(n_222), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_827), .B(n_223), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_830), .B(n_230), .Y(n_987) );
INVx1_ASAP7_75t_SL g988 ( .A(n_847), .Y(n_988) );
BUFx6f_ASAP7_75t_L g989 ( .A(n_835), .Y(n_989) );
BUFx2_ASAP7_75t_L g990 ( .A(n_847), .Y(n_990) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_840), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_856), .B(n_231), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_856), .B(n_234), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_861), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_863), .B(n_236), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_846), .B(n_237), .Y(n_996) );
AO21x2_ASAP7_75t_L g997 ( .A1(n_871), .A2(n_238), .B(n_239), .Y(n_997) );
INVx2_ASAP7_75t_L g998 ( .A(n_799), .Y(n_998) );
OR2x2_ASAP7_75t_L g999 ( .A(n_844), .B(n_240), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_799), .Y(n_1000) );
NAND4xp25_ASAP7_75t_SL g1001 ( .A(n_854), .B(n_242), .C(n_247), .D(n_248), .Y(n_1001) );
BUFx3_ASAP7_75t_L g1002 ( .A(n_814), .Y(n_1002) );
INVx3_ASAP7_75t_L g1003 ( .A(n_846), .Y(n_1003) );
INVx2_ASAP7_75t_L g1004 ( .A(n_852), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_863), .B(n_249), .Y(n_1005) );
BUFx6f_ASAP7_75t_L g1006 ( .A(n_860), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_866), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_867), .Y(n_1008) );
CKINVDCx16_ASAP7_75t_R g1009 ( .A(n_870), .Y(n_1009) );
NOR2xp33_ASAP7_75t_L g1010 ( .A(n_862), .B(n_250), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_872), .Y(n_1011) );
INVx4_ASAP7_75t_L g1012 ( .A(n_908), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1011), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_963), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_889), .B(n_873), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_926), .B(n_862), .Y(n_1016) );
HB1xp67_ASAP7_75t_L g1017 ( .A(n_899), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_927), .B(n_864), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_967), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_899), .Y(n_1020) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_890), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_959), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_902), .B(n_865), .Y(n_1023) );
BUFx2_ASAP7_75t_L g1024 ( .A(n_940), .Y(n_1024) );
INVx2_ASAP7_75t_L g1025 ( .A(n_893), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_894), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_895), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_903), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_906), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_952), .B(n_854), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_917), .Y(n_1031) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_900), .Y(n_1032) );
INVx3_ASAP7_75t_L g1033 ( .A(n_962), .Y(n_1033) );
AND2x4_ASAP7_75t_L g1034 ( .A(n_990), .B(n_860), .Y(n_1034) );
BUFx2_ASAP7_75t_L g1035 ( .A(n_945), .Y(n_1035) );
OR2x2_ASAP7_75t_L g1036 ( .A(n_920), .B(n_850), .Y(n_1036) );
INVxp67_ASAP7_75t_L g1037 ( .A(n_880), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_912), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_916), .B(n_850), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_928), .Y(n_1040) );
AND2x4_ASAP7_75t_L g1041 ( .A(n_988), .B(n_871), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_970), .B(n_254), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_955), .B(n_256), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_965), .B(n_258), .Y(n_1044) );
INVx2_ASAP7_75t_L g1045 ( .A(n_924), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_948), .B(n_260), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_900), .B(n_261), .Y(n_1047) );
INVx2_ASAP7_75t_L g1048 ( .A(n_933), .Y(n_1048) );
INVx2_ASAP7_75t_SL g1049 ( .A(n_887), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_925), .B(n_262), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_938), .Y(n_1051) );
INVxp67_ASAP7_75t_L g1052 ( .A(n_886), .Y(n_1052) );
AND2x4_ASAP7_75t_SL g1053 ( .A(n_887), .B(n_263), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_960), .Y(n_1054) );
INVx2_ASAP7_75t_L g1055 ( .A(n_942), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_925), .B(n_264), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_994), .Y(n_1057) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_947), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_980), .B(n_265), .Y(n_1059) );
AND2x4_ASAP7_75t_L g1060 ( .A(n_988), .B(n_266), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_941), .B(n_267), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_943), .B(n_272), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_968), .Y(n_1063) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_971), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_969), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_971), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_954), .B(n_277), .Y(n_1067) );
NOR2xp33_ASAP7_75t_L g1068 ( .A(n_949), .B(n_279), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_977), .Y(n_1069) );
OR2x2_ASAP7_75t_L g1070 ( .A(n_977), .B(n_281), .Y(n_1070) );
AOI22xp5_ASAP7_75t_L g1071 ( .A1(n_931), .A2(n_286), .B1(n_287), .B2(n_293), .Y(n_1071) );
AND2x4_ASAP7_75t_L g1072 ( .A(n_962), .B(n_295), .Y(n_1072) );
AND2x4_ASAP7_75t_L g1073 ( .A(n_1003), .B(n_297), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_883), .B(n_299), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_958), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_951), .B(n_300), .Y(n_1076) );
INVx3_ASAP7_75t_R g1077 ( .A(n_915), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_931), .A2(n_303), .B1(n_305), .B2(n_307), .Y(n_1078) );
BUFx6f_ASAP7_75t_L g1079 ( .A(n_953), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_905), .B(n_308), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_958), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_898), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_898), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_982), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_951), .B(n_309), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1007), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_973), .Y(n_1087) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_953), .Y(n_1088) );
AND2x4_ASAP7_75t_L g1089 ( .A(n_1003), .B(n_310), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_976), .Y(n_1090) );
INVxp67_ASAP7_75t_L g1091 ( .A(n_891), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_991), .Y(n_1092) );
AND2x4_ASAP7_75t_L g1093 ( .A(n_1006), .B(n_313), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_991), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1008), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_881), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_910), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_932), .B(n_314), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_937), .B(n_316), .Y(n_1099) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1004), .Y(n_1100) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_953), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_897), .B(n_319), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_961), .B(n_321), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_909), .B(n_322), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_914), .B(n_323), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_978), .B(n_324), .Y(n_1106) );
INVx2_ASAP7_75t_L g1107 ( .A(n_911), .Y(n_1107) );
INVx3_ASAP7_75t_SL g1108 ( .A(n_957), .Y(n_1108) );
INVx2_ASAP7_75t_L g1109 ( .A(n_921), .Y(n_1109) );
INVx3_ASAP7_75t_L g1110 ( .A(n_1009), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_881), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_936), .B(n_326), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_983), .B(n_327), .Y(n_1113) );
AND2x4_ASAP7_75t_L g1114 ( .A(n_1006), .B(n_328), .Y(n_1114) );
AND2x4_ASAP7_75t_L g1115 ( .A(n_1006), .B(n_330), .Y(n_1115) );
OR2x2_ASAP7_75t_L g1116 ( .A(n_919), .B(n_331), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_1017), .B(n_939), .Y(n_1117) );
HB1xp67_ASAP7_75t_L g1118 ( .A(n_1064), .Y(n_1118) );
INVxp33_ASAP7_75t_SL g1119 ( .A(n_1021), .Y(n_1119) );
INVx1_ASAP7_75t_SL g1120 ( .A(n_1024), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1026), .Y(n_1121) );
INVx2_ASAP7_75t_L g1122 ( .A(n_1020), .Y(n_1122) );
INVx2_ASAP7_75t_L g1123 ( .A(n_1012), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1124 ( .A(n_1058), .B(n_944), .Y(n_1124) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1012), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1035), .B(n_985), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_1013), .B(n_922), .Y(n_1127) );
INVx2_ASAP7_75t_SL g1128 ( .A(n_1049), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1110), .B(n_985), .Y(n_1129) );
NOR2xp67_ASAP7_75t_L g1130 ( .A(n_1110), .B(n_1001), .Y(n_1130) );
INVx2_ASAP7_75t_SL g1131 ( .A(n_1053), .Y(n_1131) );
OAI21xp33_ASAP7_75t_SL g1132 ( .A1(n_1033), .A2(n_882), .B(n_936), .Y(n_1132) );
HB1xp67_ASAP7_75t_L g1133 ( .A(n_1032), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1028), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1013), .B(n_929), .Y(n_1135) );
OR2x2_ASAP7_75t_L g1136 ( .A(n_1048), .B(n_956), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1029), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1052), .B(n_1010), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1091), .B(n_1010), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1025), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1027), .B(n_935), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_1014), .B(n_1000), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1031), .B(n_956), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1055), .B(n_975), .Y(n_1144) );
BUFx2_ASAP7_75t_SL g1145 ( .A(n_1072), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1040), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1051), .B(n_999), .Y(n_1147) );
HB1xp67_ASAP7_75t_L g1148 ( .A(n_1081), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1039), .B(n_1037), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1014), .B(n_998), .Y(n_1150) );
HB1xp67_ASAP7_75t_L g1151 ( .A(n_1092), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1038), .Y(n_1152) );
OR2x2_ASAP7_75t_L g1153 ( .A(n_1066), .B(n_888), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1019), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1019), .Y(n_1155) );
AND2x4_ASAP7_75t_L g1156 ( .A(n_1034), .B(n_1002), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1069), .B(n_1002), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1023), .B(n_964), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1075), .B(n_888), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1016), .B(n_913), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1063), .B(n_992), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1065), .B(n_993), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1057), .B(n_984), .Y(n_1163) );
NOR2xp33_ASAP7_75t_L g1164 ( .A(n_1108), .B(n_918), .Y(n_1164) );
NAND2x1p5_ASAP7_75t_L g1165 ( .A(n_1060), .B(n_882), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1022), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1022), .Y(n_1167) );
INVx2_ASAP7_75t_L g1168 ( .A(n_1045), .Y(n_1168) );
NAND3xp33_ASAP7_75t_L g1169 ( .A(n_1059), .B(n_885), .C(n_979), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1054), .Y(n_1170) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1054), .Y(n_1171) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1092), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1015), .Y(n_1173) );
AND2x4_ASAP7_75t_L g1174 ( .A(n_1034), .B(n_981), .Y(n_1174) );
AND2x4_ASAP7_75t_L g1175 ( .A(n_1018), .B(n_957), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1086), .Y(n_1176) );
AND2x4_ASAP7_75t_L g1177 ( .A(n_1094), .B(n_989), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1087), .B(n_984), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1033), .B(n_884), .Y(n_1179) );
INVx2_ASAP7_75t_L g1180 ( .A(n_1094), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1173), .B(n_1030), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1118), .Y(n_1182) );
INVxp67_ASAP7_75t_L g1183 ( .A(n_1133), .Y(n_1183) );
HB1xp67_ASAP7_75t_L g1184 ( .A(n_1118), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1121), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1120), .B(n_1036), .Y(n_1186) );
INVx2_ASAP7_75t_L g1187 ( .A(n_1124), .Y(n_1187) );
OAI21xp5_ASAP7_75t_L g1188 ( .A1(n_1130), .A2(n_896), .B(n_1072), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1134), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1120), .B(n_1082), .Y(n_1190) );
NOR2xp33_ASAP7_75t_L g1191 ( .A(n_1119), .B(n_1077), .Y(n_1191) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1149), .B(n_1084), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1158), .B(n_1088), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1126), .B(n_1101), .Y(n_1194) );
NAND3xp33_ASAP7_75t_L g1195 ( .A(n_1132), .B(n_979), .C(n_885), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1160), .B(n_1041), .Y(n_1196) );
NAND4xp25_ASAP7_75t_L g1197 ( .A(n_1169), .B(n_1068), .C(n_1112), .D(n_896), .Y(n_1197) );
HB1xp67_ASAP7_75t_L g1198 ( .A(n_1148), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1137), .Y(n_1199) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1117), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1152), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1151), .Y(n_1202) );
INVx3_ASAP7_75t_L g1203 ( .A(n_1123), .Y(n_1203) );
NOR2xp33_ASAP7_75t_L g1204 ( .A(n_1128), .B(n_1103), .Y(n_1204) );
OR2x2_ASAP7_75t_L g1205 ( .A(n_1151), .B(n_1084), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1206 ( .A(n_1140), .B(n_1095), .Y(n_1206) );
AOI221xp5_ASAP7_75t_L g1207 ( .A1(n_1146), .A2(n_1083), .B1(n_1087), .B2(n_1090), .C(n_1111), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1154), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1122), .B(n_1095), .Y(n_1209) );
HB1xp67_ASAP7_75t_L g1210 ( .A(n_1168), .Y(n_1210) );
INVx1_ASAP7_75t_SL g1211 ( .A(n_1145), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1155), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1143), .B(n_1096), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1176), .Y(n_1214) );
INVx2_ASAP7_75t_SL g1215 ( .A(n_1131), .Y(n_1215) );
INVx1_ASAP7_75t_SL g1216 ( .A(n_1125), .Y(n_1216) );
NAND2x1p5_ASAP7_75t_L g1217 ( .A(n_1174), .B(n_1060), .Y(n_1217) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1171), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1166), .B(n_1086), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g1220 ( .A1(n_1211), .A2(n_1164), .B1(n_1165), .B2(n_1129), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1182), .Y(n_1221) );
AOI22xp5_ASAP7_75t_SL g1222 ( .A1(n_1191), .A2(n_1174), .B1(n_1175), .B2(n_1165), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1184), .Y(n_1223) );
NAND3xp33_ASAP7_75t_L g1224 ( .A(n_1195), .B(n_1157), .C(n_1169), .Y(n_1224) );
AOI22xp5_ASAP7_75t_L g1225 ( .A1(n_1197), .A2(n_1138), .B1(n_1139), .B2(n_1144), .Y(n_1225) );
NOR2x1p5_ASAP7_75t_L g1226 ( .A(n_1195), .B(n_1161), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1205), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_1198), .B(n_1172), .Y(n_1228) );
OAI22xp5_ASAP7_75t_L g1229 ( .A1(n_1211), .A2(n_1175), .B1(n_1161), .B2(n_1162), .Y(n_1229) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1210), .Y(n_1230) );
NAND3xp33_ASAP7_75t_L g1231 ( .A(n_1202), .B(n_1157), .C(n_1135), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1206), .Y(n_1232) );
NAND3xp33_ASAP7_75t_L g1233 ( .A(n_1188), .B(n_1070), .C(n_1043), .Y(n_1233) );
NOR2xp33_ASAP7_75t_L g1234 ( .A(n_1215), .B(n_1162), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1185), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1207), .B(n_1180), .Y(n_1236) );
OR2x2_ASAP7_75t_L g1237 ( .A(n_1192), .B(n_1187), .Y(n_1237) );
INVx1_ASAP7_75t_SL g1238 ( .A(n_1186), .Y(n_1238) );
OAI22xp5_ASAP7_75t_L g1239 ( .A1(n_1217), .A2(n_1141), .B1(n_1167), .B2(n_1170), .Y(n_1239) );
NAND2xp33_ASAP7_75t_SL g1240 ( .A(n_1203), .B(n_1156), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1189), .Y(n_1241) );
INVxp67_ASAP7_75t_L g1242 ( .A(n_1190), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1199), .Y(n_1243) );
O2A1O1Ixp33_ASAP7_75t_L g1244 ( .A1(n_1224), .A2(n_1183), .B(n_1197), .C(n_1181), .Y(n_1244) );
INVx1_ASAP7_75t_SL g1245 ( .A(n_1238), .Y(n_1245) );
NOR4xp25_ASAP7_75t_L g1246 ( .A(n_1223), .B(n_1216), .C(n_1201), .D(n_1203), .Y(n_1246) );
NAND3xp33_ASAP7_75t_L g1247 ( .A(n_1222), .B(n_1214), .C(n_1212), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1227), .Y(n_1248) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_1229), .A2(n_1213), .B1(n_1216), .B2(n_1208), .C(n_1196), .Y(n_1249) );
AOI33xp33_ASAP7_75t_L g1250 ( .A1(n_1225), .A2(n_1193), .A3(n_1200), .B1(n_1194), .B2(n_1147), .B3(n_1218), .Y(n_1250) );
AOI211xp5_ASAP7_75t_SL g1251 ( .A1(n_1220), .A2(n_1204), .B(n_1061), .C(n_1062), .Y(n_1251) );
NOR2x1_ASAP7_75t_L g1252 ( .A(n_1226), .B(n_1001), .Y(n_1252) );
AOI221xp5_ASAP7_75t_L g1253 ( .A1(n_1234), .A2(n_1219), .B1(n_1163), .B2(n_1135), .C(n_1142), .Y(n_1253) );
OAI21xp33_ASAP7_75t_L g1254 ( .A1(n_1236), .A2(n_1217), .B(n_1209), .Y(n_1254) );
AOI21xp5_ASAP7_75t_L g1255 ( .A1(n_1240), .A2(n_1156), .B(n_1142), .Y(n_1255) );
OAI21xp5_ASAP7_75t_L g1256 ( .A1(n_1233), .A2(n_1071), .B(n_1102), .Y(n_1256) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_1233), .A2(n_1179), .B1(n_1153), .B2(n_1159), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1232), .B(n_1163), .Y(n_1258) );
NAND3xp33_ASAP7_75t_L g1259 ( .A(n_1231), .B(n_1090), .C(n_1177), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1244), .B(n_1242), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1250), .B(n_1235), .Y(n_1261) );
OAI221xp5_ASAP7_75t_L g1262 ( .A1(n_1246), .A2(n_1239), .B1(n_1228), .B2(n_1243), .C(n_1241), .Y(n_1262) );
OAI211xp5_ASAP7_75t_SL g1263 ( .A1(n_1252), .A2(n_1221), .B(n_1230), .C(n_1078), .Y(n_1263) );
AOI221xp5_ASAP7_75t_L g1264 ( .A1(n_1257), .A2(n_1237), .B1(n_1127), .B2(n_1177), .C(n_1178), .Y(n_1264) );
AOI222xp33_ASAP7_75t_L g1265 ( .A1(n_1245), .A2(n_1127), .B1(n_1178), .B2(n_1150), .C1(n_1044), .C2(n_1056), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1253), .B(n_1136), .Y(n_1266) );
OAI221xp5_ASAP7_75t_L g1267 ( .A1(n_1247), .A2(n_1116), .B1(n_1080), .B2(n_1150), .C(n_1105), .Y(n_1267) );
OAI211xp5_ASAP7_75t_L g1268 ( .A1(n_1254), .A2(n_1099), .B(n_1098), .C(n_972), .Y(n_1268) );
NOR2xp33_ASAP7_75t_L g1269 ( .A(n_1258), .B(n_1046), .Y(n_1269) );
BUFx2_ASAP7_75t_L g1270 ( .A(n_1249), .Y(n_1270) );
NAND4xp25_ASAP7_75t_L g1271 ( .A(n_1270), .B(n_1251), .C(n_1256), .D(n_1259), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1266), .Y(n_1272) );
AOI221xp5_ASAP7_75t_L g1273 ( .A1(n_1260), .A2(n_1248), .B1(n_1255), .B2(n_1050), .C(n_1047), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1261), .Y(n_1274) );
NAND4xp25_ASAP7_75t_L g1275 ( .A(n_1263), .B(n_974), .C(n_1074), .D(n_1113), .Y(n_1275) );
AOI21xp5_ASAP7_75t_L g1276 ( .A1(n_1262), .A2(n_923), .B(n_1089), .Y(n_1276) );
OAI21xp5_ASAP7_75t_L g1277 ( .A1(n_1268), .A2(n_1005), .B(n_995), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1269), .Y(n_1278) );
AOI211xp5_ASAP7_75t_L g1279 ( .A1(n_1274), .A2(n_1267), .B(n_1264), .C(n_1104), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1278), .B(n_1272), .Y(n_1280) );
INVx2_ASAP7_75t_L g1281 ( .A(n_1277), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1271), .B(n_1100), .Y(n_1282) );
NOR3x1_ASAP7_75t_L g1283 ( .A(n_1275), .B(n_1265), .C(n_923), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1273), .B(n_1042), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1280), .Y(n_1285) );
AOI221xp5_ASAP7_75t_L g1286 ( .A1(n_1281), .A2(n_1276), .B1(n_1041), .B2(n_1067), .C(n_966), .Y(n_1286) );
OAI221xp5_ASAP7_75t_L g1287 ( .A1(n_1279), .A2(n_950), .B1(n_946), .B2(n_930), .C(n_1106), .Y(n_1287) );
NAND4xp25_ASAP7_75t_SL g1288 ( .A(n_1282), .B(n_1076), .C(n_1085), .D(n_950), .Y(n_1288) );
OR2x2_ASAP7_75t_L g1289 ( .A(n_1284), .B(n_1097), .Y(n_1289) );
INVx1_ASAP7_75t_SL g1290 ( .A(n_1285), .Y(n_1290) );
BUFx2_ASAP7_75t_L g1291 ( .A(n_1289), .Y(n_1291) );
AND3x4_ASAP7_75t_L g1292 ( .A(n_1286), .B(n_1283), .C(n_1073), .Y(n_1292) );
XNOR2xp5_ASAP7_75t_L g1293 ( .A(n_1287), .B(n_1089), .Y(n_1293) );
INVx2_ASAP7_75t_L g1294 ( .A(n_1290), .Y(n_1294) );
HB1xp67_ASAP7_75t_L g1295 ( .A(n_1291), .Y(n_1295) );
XNOR2x1_ASAP7_75t_L g1296 ( .A(n_1292), .B(n_1288), .Y(n_1296) );
OAI22xp5_ASAP7_75t_L g1297 ( .A1(n_1294), .A2(n_1293), .B1(n_1073), .B2(n_1079), .Y(n_1297) );
OAI332xp33_ASAP7_75t_L g1298 ( .A1(n_1296), .A2(n_946), .A3(n_930), .B1(n_892), .B2(n_996), .B3(n_1097), .C1(n_1109), .C2(n_1107), .Y(n_1298) );
INVx2_ASAP7_75t_L g1299 ( .A(n_1295), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1299), .Y(n_1300) );
AOI21xp5_ASAP7_75t_L g1301 ( .A1(n_1297), .A2(n_996), .B(n_934), .Y(n_1301) );
OAI21x1_ASAP7_75t_SL g1302 ( .A1(n_1298), .A2(n_934), .B(n_1114), .Y(n_1302) );
HB1xp67_ASAP7_75t_L g1303 ( .A(n_1300), .Y(n_1303) );
AOI21xp5_ASAP7_75t_L g1304 ( .A1(n_1302), .A2(n_986), .B(n_987), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1305 ( .A(n_1301), .B(n_1079), .Y(n_1305) );
XNOR2xp5_ASAP7_75t_L g1306 ( .A(n_1303), .B(n_1115), .Y(n_1306) );
OAI21xp5_ASAP7_75t_L g1307 ( .A1(n_1305), .A2(n_907), .B(n_1114), .Y(n_1307) );
AO21x2_ASAP7_75t_L g1308 ( .A1(n_1304), .A2(n_904), .B(n_901), .Y(n_1308) );
AOI221xp5_ASAP7_75t_L g1309 ( .A1(n_1306), .A2(n_1115), .B1(n_1093), .B2(n_1079), .C(n_997), .Y(n_1309) );
AOI21xp5_ASAP7_75t_L g1310 ( .A1(n_1308), .A2(n_1093), .B(n_997), .Y(n_1310) );
OR2x6_ASAP7_75t_L g1311 ( .A(n_1307), .B(n_989), .Y(n_1311) );
AOI22xp33_ASAP7_75t_L g1312 ( .A1(n_1309), .A2(n_1311), .B1(n_1310), .B2(n_989), .Y(n_1312) );
endmodule