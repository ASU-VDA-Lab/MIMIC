module real_aes_7962_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_1066;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_1021;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_370;
wire n_1078;
wire n_384;
wire n_938;
wire n_744;
wire n_352;
wire n_935;
wire n_824;
wire n_875;
wire n_467;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_1053;
wire n_466;
wire n_636;
wire n_559;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_755;
wire n_532;
wire n_1025;
wire n_656;
wire n_746;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_455;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_1081;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_769;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_1041;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1003;
wire n_1000;
wire n_1028;
wire n_366;
wire n_727;
wire n_1014;
wire n_397;
wire n_749;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_899;
wire n_637;
wire n_526;
wire n_653;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_967;
wire n_719;
wire n_1045;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g491 ( .A1(n_0), .A2(n_260), .B1(n_492), .B2(n_494), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_1), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g1044 ( .A(n_2), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_3), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_4), .A2(n_48), .B1(n_678), .B2(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_5), .A2(n_321), .B1(n_570), .B2(n_1072), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_6), .A2(n_121), .B1(n_570), .B2(n_572), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_7), .Y(n_910) );
AO22x2_ASAP7_75t_L g375 ( .A1(n_8), .A2(n_209), .B1(n_376), .B2(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g1033 ( .A(n_8), .Y(n_1033) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_9), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_10), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_11), .A2(n_264), .B1(n_434), .B2(n_496), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_12), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_13), .A2(n_20), .B1(n_511), .B2(n_769), .Y(n_1077) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_14), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_15), .A2(n_226), .B1(n_579), .B2(n_580), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_16), .A2(n_141), .B1(n_631), .B2(n_680), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_17), .B(n_555), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_18), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_19), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_21), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_22), .A2(n_328), .B1(n_796), .B2(n_798), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_23), .A2(n_331), .B1(n_672), .B2(n_1002), .Y(n_1001) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_24), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_25), .Y(n_444) );
AOI222xp33_ASAP7_75t_L g707 ( .A1(n_26), .A2(n_50), .B1(n_313), .B2(n_504), .C1(n_708), .C2(n_709), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_27), .A2(n_108), .B1(n_484), .B2(n_924), .Y(n_923) );
CKINVDCx20_ASAP7_75t_R g947 ( .A(n_28), .Y(n_947) );
AO22x2_ASAP7_75t_L g379 ( .A1(n_29), .A2(n_94), .B1(n_376), .B2(n_380), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_30), .A2(n_344), .B1(n_880), .B2(n_899), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_31), .A2(n_195), .B1(n_574), .B2(n_980), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_32), .A2(n_228), .B1(n_451), .B2(n_484), .Y(n_704) );
INVx1_ASAP7_75t_L g723 ( .A(n_33), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_34), .A2(n_99), .B1(n_571), .B2(n_588), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_35), .A2(n_49), .B1(n_425), .B2(n_580), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_36), .A2(n_145), .B1(n_532), .B2(n_749), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_37), .A2(n_251), .B1(n_572), .B2(n_597), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_38), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g983 ( .A(n_39), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_40), .B(n_819), .Y(n_818) );
AOI22xp5_ASAP7_75t_SL g498 ( .A1(n_41), .A2(n_499), .B1(n_500), .B2(n_537), .Y(n_498) );
INVx1_ASAP7_75t_L g537 ( .A(n_41), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_42), .A2(n_268), .B1(n_402), .B2(n_407), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_43), .A2(n_203), .B1(n_402), .B2(n_479), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_44), .A2(n_306), .B1(n_640), .B2(n_734), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_45), .A2(n_225), .B1(n_531), .B2(n_532), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_46), .B(n_840), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_47), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_51), .A2(n_261), .B1(n_583), .B2(n_586), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_52), .B(n_555), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_53), .A2(n_291), .B1(n_751), .B2(n_752), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_54), .A2(n_546), .B1(n_589), .B2(n_590), .Y(n_545) );
INVx1_ASAP7_75t_L g589 ( .A(n_54), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_55), .A2(n_250), .B1(n_636), .B2(n_637), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g1047 ( .A(n_56), .Y(n_1047) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_57), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_58), .A2(n_273), .B1(n_583), .B2(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_59), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g982 ( .A(n_60), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_61), .A2(n_89), .B1(n_484), .B2(n_814), .Y(n_1051) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_62), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_63), .A2(n_84), .B1(n_796), .B2(n_953), .Y(n_952) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_64), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_65), .A2(n_231), .B1(n_509), .B2(n_787), .Y(n_968) );
AOI222xp33_ASAP7_75t_L g677 ( .A1(n_66), .A2(n_256), .B1(n_311), .B2(n_504), .C1(n_555), .C2(n_678), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g837 ( .A1(n_67), .A2(n_237), .B1(n_402), .B2(n_407), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_68), .A2(n_267), .B1(n_487), .B2(n_706), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_69), .A2(n_199), .B1(n_556), .B2(n_709), .Y(n_815) );
INVx1_ASAP7_75t_L g593 ( .A(n_70), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_71), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_72), .A2(n_115), .B1(n_518), .B2(n_521), .Y(n_771) );
AO22x2_ASAP7_75t_L g383 ( .A1(n_73), .A2(n_232), .B1(n_376), .B2(n_377), .Y(n_383) );
INVx1_ASAP7_75t_L g1030 ( .A(n_73), .Y(n_1030) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_74), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_75), .A2(n_76), .B1(n_496), .B2(n_706), .Y(n_1056) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_77), .A2(n_351), .B(n_359), .C(n_1035), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_78), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_79), .A2(n_92), .B1(n_581), .B2(n_603), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_80), .A2(n_214), .B1(n_403), .B2(n_407), .Y(n_474) );
OA22x2_ASAP7_75t_L g364 ( .A1(n_81), .A2(n_365), .B1(n_366), .B2(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_81), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_82), .A2(n_134), .B1(n_796), .B2(n_980), .Y(n_979) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_83), .Y(n_916) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_85), .A2(n_302), .B1(n_672), .B2(n_673), .C(n_674), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_86), .A2(n_128), .B1(n_507), .B2(n_509), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g1048 ( .A(n_87), .Y(n_1048) );
CKINVDCx20_ASAP7_75t_R g1042 ( .A(n_88), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_90), .A2(n_167), .B1(n_414), .B2(n_631), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g525 ( .A1(n_91), .A2(n_329), .B1(n_526), .B2(n_528), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_93), .A2(n_135), .B1(n_432), .B2(n_637), .Y(n_850) );
INVx1_ASAP7_75t_L g1034 ( .A(n_94), .Y(n_1034) );
AOI22xp33_ASAP7_75t_SL g513 ( .A1(n_95), .A2(n_151), .B1(n_414), .B2(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_96), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_97), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g918 ( .A(n_98), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_100), .A2(n_205), .B1(n_637), .B2(n_880), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_101), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_102), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_103), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g998 ( .A(n_104), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_105), .A2(n_263), .B1(n_487), .B2(n_847), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_106), .A2(n_283), .B1(n_667), .B2(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_107), .A2(n_117), .B1(n_875), .B2(n_876), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_109), .A2(n_280), .B1(n_453), .B2(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g912 ( .A(n_110), .Y(n_912) );
AOI22xp33_ASAP7_75t_SL g896 ( .A1(n_111), .A2(n_162), .B1(n_514), .B2(n_680), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_112), .B(n_967), .Y(n_966) );
AOI22xp33_ASAP7_75t_SL g900 ( .A1(n_113), .A2(n_275), .B1(n_496), .B2(n_798), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_114), .A2(n_305), .B1(n_403), .B2(n_514), .Y(n_1045) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_116), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_118), .A2(n_309), .B1(n_494), .B2(n_953), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_119), .A2(n_284), .B1(n_479), .B2(n_787), .Y(n_786) );
AOI22xp33_ASAP7_75t_SL g630 ( .A1(n_120), .A2(n_297), .B1(n_407), .B2(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g1000 ( .A1(n_122), .A2(n_179), .B1(n_709), .B2(n_787), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_123), .A2(n_303), .B1(n_535), .B2(n_574), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_124), .A2(n_174), .B1(n_629), .B2(n_1002), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_125), .A2(n_183), .B1(n_640), .B2(n_794), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_126), .A2(n_191), .B1(n_600), .B2(n_829), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_127), .Y(n_606) );
INVxp67_ASAP7_75t_L g1064 ( .A(n_129), .Y(n_1064) );
XNOR2x2_ASAP7_75t_L g1065 ( .A(n_129), .B(n_1066), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_130), .B(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_131), .A2(n_190), .B1(n_446), .B2(n_597), .Y(n_925) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_132), .Y(n_960) );
AND2x6_ASAP7_75t_L g353 ( .A(n_133), .B(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g1027 ( .A(n_133), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_136), .A2(n_219), .B1(n_570), .B2(n_873), .Y(n_872) );
AOI22xp33_ASAP7_75t_SL g768 ( .A1(n_137), .A2(n_252), .B1(n_509), .B2(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_138), .A2(n_160), .B1(n_487), .B2(n_599), .Y(n_1055) );
INVx1_ASAP7_75t_L g869 ( .A(n_139), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_140), .A2(n_240), .B1(n_603), .B2(n_1053), .Y(n_1052) );
CKINVDCx20_ASAP7_75t_R g937 ( .A(n_142), .Y(n_937) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_143), .A2(n_238), .B1(n_425), .B2(n_426), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_144), .A2(n_169), .B1(n_794), .B2(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_146), .A2(n_255), .B1(n_402), .B2(n_623), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_147), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_148), .A2(n_279), .B1(n_599), .B2(n_600), .Y(n_598) );
AOI222xp33_ASAP7_75t_L g1078 ( .A1(n_149), .A2(n_196), .B1(n_314), .B2(n_396), .C1(n_708), .C2(n_1053), .Y(n_1078) );
NAND2xp5_ASAP7_75t_SL g895 ( .A(n_150), .B(n_672), .Y(n_895) );
AO22x2_ASAP7_75t_L g385 ( .A1(n_152), .A2(n_222), .B1(n_376), .B2(n_380), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g1031 ( .A(n_152), .B(n_1032), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_153), .A2(n_181), .B1(n_432), .B2(n_668), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_154), .A2(n_164), .B1(n_574), .B2(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_155), .A2(n_236), .B1(n_442), .B2(n_532), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g986 ( .A(n_156), .Y(n_986) );
AOI211xp5_ASAP7_75t_L g962 ( .A1(n_157), .A2(n_396), .B(n_963), .C(n_969), .Y(n_962) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_158), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_159), .A2(n_327), .B1(n_583), .B2(n_586), .Y(n_799) );
AOI22xp33_ASAP7_75t_SL g892 ( .A1(n_161), .A2(n_246), .B1(n_407), .B2(n_556), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_163), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g939 ( .A(n_165), .Y(n_939) );
CKINVDCx20_ASAP7_75t_R g941 ( .A(n_166), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g972 ( .A(n_168), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_170), .Y(n_466) );
AOI22xp33_ASAP7_75t_SL g845 ( .A1(n_171), .A2(n_211), .B1(n_581), .B2(n_668), .Y(n_845) );
AOI22xp33_ASAP7_75t_SL g902 ( .A1(n_172), .A2(n_188), .B1(n_581), .B2(n_875), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_173), .A2(n_215), .B1(n_489), .B2(n_496), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_175), .A2(n_212), .B1(n_518), .B2(n_521), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_176), .A2(n_712), .B1(n_738), .B2(n_739), .Y(n_711) );
INVx1_ASAP7_75t_L g738 ( .A(n_176), .Y(n_738) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_177), .A2(n_332), .B1(n_426), .B2(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g505 ( .A(n_178), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_180), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_182), .Y(n_920) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_184), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_185), .A2(n_339), .B1(n_434), .B2(n_496), .Y(n_696) );
XOR2xp5_ASAP7_75t_L g1036 ( .A(n_186), .B(n_1037), .Y(n_1036) );
CKINVDCx20_ASAP7_75t_R g996 ( .A(n_187), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_189), .A2(n_266), .B1(n_431), .B2(n_434), .Y(n_430) );
AOI22xp33_ASAP7_75t_SL g849 ( .A1(n_192), .A2(n_274), .B1(n_425), .B2(n_636), .Y(n_849) );
AOI22xp33_ASAP7_75t_SL g898 ( .A1(n_193), .A2(n_325), .B1(n_574), .B2(n_899), .Y(n_898) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_194), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g634 ( .A1(n_197), .A2(n_235), .B1(n_484), .B2(n_487), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g915 ( .A(n_198), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_200), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_201), .A2(n_208), .B1(n_556), .B2(n_944), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_202), .A2(n_304), .B1(n_453), .B2(n_531), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_204), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_206), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_207), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_210), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_213), .A2(n_296), .B1(n_434), .B2(n_496), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_216), .A2(n_301), .B1(n_583), .B2(n_847), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_217), .B(n_673), .Y(n_894) );
XNOR2x2_ASAP7_75t_L g744 ( .A(n_218), .B(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_220), .A2(n_336), .B1(n_489), .B2(n_977), .Y(n_1005) );
INVx2_ASAP7_75t_L g358 ( .A(n_221), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g955 ( .A1(n_223), .A2(n_234), .B1(n_583), .B2(n_924), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_224), .B(n_521), .Y(n_841) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_227), .A2(n_346), .B1(n_432), .B2(n_489), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_229), .Y(n_754) );
AOI22xp33_ASAP7_75t_SL g639 ( .A1(n_230), .A2(n_342), .B1(n_572), .B2(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_233), .A2(n_318), .B1(n_515), .B2(n_623), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_239), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_241), .A2(n_277), .B1(n_425), .B2(n_580), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_242), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_243), .A2(n_337), .B1(n_574), .B2(n_576), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_244), .B(n_701), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_245), .A2(n_646), .B1(n_681), .B2(n_682), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_245), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_247), .A2(n_343), .B1(n_442), .B2(n_446), .Y(n_951) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_248), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g1041 ( .A(n_249), .Y(n_1041) );
OA22x2_ASAP7_75t_L g989 ( .A1(n_253), .A2(n_990), .B1(n_991), .B2(n_1010), .Y(n_989) );
CKINVDCx20_ASAP7_75t_R g990 ( .A(n_253), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_254), .A2(n_276), .B1(n_798), .B2(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g376 ( .A(n_257), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_257), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_258), .A2(n_341), .B1(n_484), .B2(n_603), .Y(n_956) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_259), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_262), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g985 ( .A(n_265), .Y(n_985) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_269), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_270), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g930 ( .A(n_271), .Y(n_930) );
CKINVDCx20_ASAP7_75t_R g994 ( .A(n_272), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_278), .B(n_701), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_281), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g827 ( .A1(n_282), .A2(n_335), .B1(n_492), .B2(n_494), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_285), .A2(n_300), .B1(n_453), .B2(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_286), .A2(n_323), .B1(n_487), .B2(n_489), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_287), .A2(n_310), .B1(n_511), .B2(n_515), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_288), .Y(n_720) );
AND2x2_ASAP7_75t_L g357 ( .A(n_289), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g724 ( .A(n_290), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_292), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_293), .Y(n_904) );
INVx1_ASAP7_75t_L g354 ( .A(n_294), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_295), .Y(n_758) );
OA22x2_ASAP7_75t_L g616 ( .A1(n_298), .A2(n_617), .B1(n_618), .B2(n_642), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_298), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_299), .B(n_629), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_307), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_308), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g970 ( .A(n_312), .Y(n_970) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_315), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_316), .Y(n_864) );
INVx1_ASAP7_75t_L g957 ( .A(n_317), .Y(n_957) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_319), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_320), .B(n_509), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_322), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_324), .A2(n_330), .B1(n_535), .B2(n_824), .Y(n_1074) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_326), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_333), .Y(n_653) );
INVx1_ASAP7_75t_L g497 ( .A(n_334), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_338), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_340), .B(n_556), .Y(n_721) );
OA22x2_ASAP7_75t_SL g853 ( .A1(n_345), .A2(n_854), .B1(n_855), .B2(n_881), .Y(n_853) );
INVx1_ASAP7_75t_L g881 ( .A(n_345), .Y(n_881) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_347), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_348), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_349), .Y(n_719) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_354), .Y(n_1026) );
OAI21xp5_ASAP7_75t_L g1062 ( .A1(n_355), .A2(n_1025), .B(n_1063), .Y(n_1062) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_685), .B1(n_1020), .B2(n_1021), .C(n_1022), .Y(n_359) );
INVx1_ASAP7_75t_L g1020 ( .A(n_360), .Y(n_1020) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_540), .B1(n_683), .B2(n_684), .Y(n_360) );
INVx1_ASAP7_75t_L g683 ( .A(n_361), .Y(n_683) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_460), .B2(n_539), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_422), .Y(n_367) );
NOR3xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_393), .C(n_411), .Y(n_368) );
OAI22xp5_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_386), .B1(n_387), .B2(n_392), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_370), .A2(n_387), .B1(n_549), .B2(n_550), .Y(n_548) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g859 ( .A(n_371), .Y(n_859) );
INVx1_ASAP7_75t_SL g938 ( .A(n_371), .Y(n_938) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx3_ASAP7_75t_L g467 ( .A(n_372), .Y(n_467) );
OAI221xp5_ASAP7_75t_L g605 ( .A1(n_372), .A2(n_389), .B1(n_606), .B2(n_607), .C(n_608), .Y(n_605) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_372), .Y(n_781) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_381), .Y(n_372) );
INVx2_ASAP7_75t_L g454 ( .A(n_373), .Y(n_454) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_379), .Y(n_373) );
AND2x2_ASAP7_75t_L g391 ( .A(n_374), .B(n_379), .Y(n_391) );
AND2x2_ASAP7_75t_L g433 ( .A(n_374), .B(n_417), .Y(n_433) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g398 ( .A(n_375), .B(n_379), .Y(n_398) );
AND2x2_ASAP7_75t_L g406 ( .A(n_375), .B(n_385), .Y(n_406) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_378), .Y(n_380) );
INVx2_ASAP7_75t_L g417 ( .A(n_379), .Y(n_417) );
INVx1_ASAP7_75t_L g437 ( .A(n_379), .Y(n_437) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_382), .B(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g432 ( .A(n_382), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g520 ( .A(n_382), .B(n_454), .Y(n_520) );
AND2x6_ASAP7_75t_L g522 ( .A(n_382), .B(n_391), .Y(n_522) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g400 ( .A(n_383), .Y(n_400) );
INVx1_ASAP7_75t_L g405 ( .A(n_383), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_383), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_383), .B(n_385), .Y(n_438) );
AND2x2_ASAP7_75t_L g399 ( .A(n_384), .B(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g429 ( .A(n_385), .B(n_410), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_387), .A2(n_467), .B1(n_715), .B2(n_716), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_387), .A2(n_858), .B1(n_859), .B2(n_860), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_387), .A2(n_779), .B1(n_915), .B2(n_916), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_387), .A2(n_937), .B1(n_938), .B2(n_939), .Y(n_936) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx3_ASAP7_75t_L g965 ( .A(n_389), .Y(n_965) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g470 ( .A(n_390), .Y(n_470) );
AND2x4_ASAP7_75t_L g425 ( .A(n_391), .B(n_399), .Y(n_425) );
AND2x2_ASAP7_75t_L g428 ( .A(n_391), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_391), .B(n_429), .Y(n_655) );
OAI21xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B(n_401), .Y(n_393) );
OAI21xp5_ASAP7_75t_SL g609 ( .A1(n_395), .A2(n_610), .B(n_611), .Y(n_609) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_395), .A2(n_621), .B(n_622), .Y(n_620) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx4_ASAP7_75t_L g472 ( .A(n_397), .Y(n_472) );
INVx2_ASAP7_75t_L g718 ( .A(n_397), .Y(n_718) );
INVx2_ASAP7_75t_L g762 ( .A(n_397), .Y(n_762) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_397), .Y(n_814) );
AND2x6_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
AND2x4_ASAP7_75t_L g408 ( .A(n_398), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g565 ( .A(n_398), .Y(n_565) );
AND2x2_ASAP7_75t_L g443 ( .A(n_399), .B(n_433), .Y(n_443) );
AND2x6_ASAP7_75t_L g453 ( .A(n_399), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g508 ( .A(n_402), .Y(n_508) );
BUFx4f_ASAP7_75t_SL g708 ( .A(n_402), .Y(n_708) );
BUFx12f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_403), .Y(n_556) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_403), .Y(n_766) );
AND2x4_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g416 ( .A(n_405), .B(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g415 ( .A(n_406), .B(n_416), .Y(n_415) );
NAND2x1p5_ASAP7_75t_L g420 ( .A(n_406), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g515 ( .A(n_406), .B(n_516), .Y(n_515) );
BUFx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_408), .Y(n_511) );
BUFx2_ASAP7_75t_SL g709 ( .A(n_408), .Y(n_709) );
INVx1_ASAP7_75t_L g566 ( .A(n_409), .Y(n_566) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B1(n_418), .B2(n_419), .Y(n_411) );
OAI221xp5_ASAP7_75t_SL g551 ( .A1(n_413), .A2(n_503), .B1(n_552), .B2(n_553), .C(n_554), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_415), .Y(n_479) );
BUFx4f_ASAP7_75t_SL g623 ( .A(n_415), .Y(n_623) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_415), .Y(n_680) );
BUFx2_ASAP7_75t_L g1053 ( .A(n_415), .Y(n_1053) );
INVx1_ASAP7_75t_L g421 ( .A(n_417), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_419), .A2(n_918), .B1(n_919), .B2(n_920), .Y(n_917) );
BUFx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_420), .A2(n_476), .B1(n_477), .B2(n_480), .Y(n_475) );
INVx4_ASAP7_75t_L g560 ( .A(n_420), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_420), .A2(n_564), .B1(n_675), .B2(n_676), .Y(n_674) );
AND2x2_ASAP7_75t_L g600 ( .A(n_421), .B(n_448), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_439), .C(n_449), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_430), .Y(n_423) );
INVx6_ASAP7_75t_L g493 ( .A(n_425), .Y(n_493) );
BUFx3_ASAP7_75t_L g579 ( .A(n_425), .Y(n_579) );
BUFx3_ASAP7_75t_L g603 ( .A(n_425), .Y(n_603) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g494 ( .A(n_427), .Y(n_494) );
BUFx3_ASAP7_75t_L g575 ( .A(n_427), .Y(n_575) );
INVx5_ASAP7_75t_L g599 ( .A(n_427), .Y(n_599) );
INVx4_ASAP7_75t_L g636 ( .A(n_427), .Y(n_636) );
INVx8_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_429), .B(n_433), .Y(n_459) );
AND2x2_ASAP7_75t_L g485 ( .A(n_429), .B(n_433), .Y(n_485) );
INVx1_ASAP7_75t_L g670 ( .A(n_431), .Y(n_670) );
BUFx2_ASAP7_75t_L g873 ( .A(n_431), .Y(n_873) );
BUFx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx3_ASAP7_75t_L g496 ( .A(n_432), .Y(n_496) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_432), .Y(n_585) );
INVx2_ASAP7_75t_L g830 ( .A(n_432), .Y(n_830) );
BUFx3_ASAP7_75t_L g929 ( .A(n_432), .Y(n_929) );
AND2x4_ASAP7_75t_L g447 ( .A(n_433), .B(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_L g576 ( .A(n_435), .Y(n_576) );
BUFx4f_ASAP7_75t_SL g731 ( .A(n_435), .Y(n_731) );
BUFx2_ASAP7_75t_L g752 ( .A(n_435), .Y(n_752) );
BUFx2_ASAP7_75t_L g798 ( .A(n_435), .Y(n_798) );
INVx6_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g637 ( .A(n_436), .Y(n_637) );
INVx1_ASAP7_75t_L g953 ( .A(n_436), .Y(n_953) );
INVx1_ASAP7_75t_SL g980 ( .A(n_436), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_436), .A2(n_564), .B1(n_1047), .B2(n_1048), .Y(n_1046) );
OR2x6_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g516 ( .A(n_437), .Y(n_516) );
INVx1_ASAP7_75t_L g448 ( .A(n_438), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_444), .B2(n_445), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g488 ( .A(n_443), .Y(n_488) );
BUFx2_ASAP7_75t_SL g531 ( .A(n_443), .Y(n_531) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_443), .Y(n_571) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
BUFx2_ASAP7_75t_L g489 ( .A(n_447), .Y(n_489) );
BUFx2_ASAP7_75t_SL g532 ( .A(n_447), .Y(n_532) );
BUFx3_ASAP7_75t_L g588 ( .A(n_447), .Y(n_588) );
BUFx3_ASAP7_75t_L g706 ( .A(n_447), .Y(n_706) );
BUFx3_ASAP7_75t_L g847 ( .A(n_447), .Y(n_847) );
BUFx3_ASAP7_75t_L g876 ( .A(n_447), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_455), .B1(n_456), .B2(n_457), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx5_ASAP7_75t_SL g668 ( .A(n_452), .Y(n_668) );
INVx4_ASAP7_75t_L g824 ( .A(n_452), .Y(n_824) );
INVx11_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx11_ASAP7_75t_L g527 ( .A(n_453), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_457), .A2(n_493), .B1(n_758), .B2(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g663 ( .A(n_458), .Y(n_663) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g539 ( .A(n_460), .Y(n_539) );
OA22x2_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B1(n_498), .B2(n_538), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
XOR2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_497), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_481), .Y(n_463) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_471), .C(n_475), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B1(n_468), .B2(n_469), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_467), .A2(n_699), .B1(n_1041), .B2(n_1042), .Y(n_1040) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_SL g699 ( .A(n_470), .Y(n_699) );
INVx2_ASAP7_75t_L g783 ( .A(n_470), .Y(n_783) );
OAI21xp5_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_473), .B(n_474), .Y(n_471) );
INVx4_ASAP7_75t_L g504 ( .A(n_472), .Y(n_504) );
BUFx2_ASAP7_75t_L g942 ( .A(n_472), .Y(n_942) );
OAI221xp5_ASAP7_75t_L g717 ( .A1(n_477), .A2(n_718), .B1(n_719), .B2(n_720), .C(n_721), .Y(n_717) );
INVx2_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_SL g971 ( .A(n_478), .Y(n_971) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g919 ( .A(n_479), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_490), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_486), .Y(n_482) );
INVx1_ASAP7_75t_L g735 ( .A(n_484), .Y(n_735) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx3_ASAP7_75t_L g529 ( .A(n_485), .Y(n_529) );
BUFx3_ASAP7_75t_L g581 ( .A(n_485), .Y(n_581) );
BUFx3_ASAP7_75t_L g794 ( .A(n_485), .Y(n_794) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g597 ( .A(n_488), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_495), .Y(n_490) );
INVxp67_ASAP7_75t_L g661 ( .A(n_492), .Y(n_661) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g535 ( .A(n_493), .Y(n_535) );
INVx3_ASAP7_75t_L g640 ( .A(n_493), .Y(n_640) );
INVx2_ASAP7_75t_L g899 ( .A(n_493), .Y(n_899) );
INVx1_ASAP7_75t_L g538 ( .A(n_498), .Y(n_538) );
INVx1_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_501), .B(n_523), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_512), .Y(n_501) );
OAI21xp5_ASAP7_75t_SL g502 ( .A1(n_503), .A2(n_505), .B(n_506), .Y(n_502) );
OAI21xp33_ASAP7_75t_SL g784 ( .A1(n_503), .A2(n_785), .B(n_786), .Y(n_784) );
OAI221xp5_ASAP7_75t_L g861 ( .A1(n_503), .A2(n_862), .B1(n_863), .B2(n_864), .C(n_865), .Y(n_861) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g973 ( .A(n_507), .Y(n_973) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_517), .Y(n_512) );
BUFx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx3_ASAP7_75t_L g631 ( .A(n_515), .Y(n_631) );
INVx1_ASAP7_75t_L g770 ( .A(n_515), .Y(n_770) );
BUFx2_ASAP7_75t_L g787 ( .A(n_515), .Y(n_787) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx5_ASAP7_75t_L g629 ( .A(n_519), .Y(n_629) );
INVx2_ASAP7_75t_L g701 ( .A(n_519), .Y(n_701) );
INVx2_ASAP7_75t_L g840 ( .A(n_519), .Y(n_840) );
INVx4_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_SL g627 ( .A(n_522), .Y(n_627) );
BUFx2_ASAP7_75t_L g673 ( .A(n_522), .Y(n_673) );
BUFx4f_ASAP7_75t_L g819 ( .A(n_522), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_533), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_530), .Y(n_524) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx4_ASAP7_75t_L g572 ( .A(n_527), .Y(n_572) );
INVx4_ASAP7_75t_L g875 ( .A(n_527), .Y(n_875) );
INVx2_ASAP7_75t_SL g924 ( .A(n_527), .Y(n_924) );
OAI21xp33_ASAP7_75t_SL g1043 ( .A1(n_527), .A2(n_1044), .B(n_1045), .Y(n_1043) );
BUFx4f_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g1073 ( .A(n_529), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
INVx1_ASAP7_75t_L g684 ( .A(n_540), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B1(n_612), .B2(n_613), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OAI22xp5_ASAP7_75t_SL g543 ( .A1(n_544), .A2(n_545), .B1(n_591), .B2(n_592), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g590 ( .A(n_546), .Y(n_590) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_567), .Y(n_546) );
NOR3xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .C(n_557), .Y(n_547) );
BUFx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g789 ( .A(n_556), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_561), .B2(n_562), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_559), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_559), .A2(n_946), .B1(n_947), .B2(n_948), .Y(n_945) );
INVx3_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g868 ( .A(n_560), .Y(n_868) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g948 ( .A(n_563), .Y(n_948) );
CKINVDCx16_ASAP7_75t_R g563 ( .A(n_564), .Y(n_563) );
BUFx2_ASAP7_75t_L g725 ( .A(n_564), .Y(n_725) );
OR2x6_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_577), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_573), .Y(n_568) );
BUFx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx3_ASAP7_75t_L g729 ( .A(n_571), .Y(n_729) );
BUFx6f_ASAP7_75t_L g749 ( .A(n_571), .Y(n_749) );
INVx3_ASAP7_75t_L g978 ( .A(n_571), .Y(n_978) );
INVx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVxp67_ASAP7_75t_L g657 ( .A(n_576), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_582), .Y(n_577) );
BUFx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx4_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_584), .A2(n_754), .B1(n_755), .B2(n_756), .Y(n_753) );
INVx4_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_587), .A2(n_649), .B1(n_650), .B2(n_651), .Y(n_648) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_588), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_591), .A2(n_592), .B1(n_616), .B2(n_643), .Y(n_615) );
INVx2_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
XNOR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
NOR4xp75_ASAP7_75t_L g594 ( .A(n_595), .B(n_601), .C(n_605), .D(n_609), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVxp67_ASAP7_75t_L g650 ( .A(n_597), .Y(n_650) );
BUFx6f_ASAP7_75t_L g880 ( .A(n_599), .Y(n_880) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI22xp5_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_615), .B1(n_644), .B2(n_645), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g643 ( .A(n_616), .Y(n_643) );
INVx1_ASAP7_75t_L g642 ( .A(n_618), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_632), .Y(n_618) );
NOR2xp67_ASAP7_75t_L g619 ( .A(n_620), .B(n_624), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_628), .C(n_630), .Y(n_624) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g1002 ( .A(n_627), .Y(n_1002) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_629), .Y(n_672) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_633), .B(n_638), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_636), .Y(n_751) );
INVx2_ASAP7_75t_L g797 ( .A(n_636), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g682 ( .A(n_646), .Y(n_682) );
AND4x1_ASAP7_75t_L g646 ( .A(n_647), .B(n_658), .C(n_671), .D(n_677), .Y(n_646) );
NOR2xp33_ASAP7_75t_SL g647 ( .A(n_648), .B(n_652), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B1(n_656), .B2(n_657), .Y(n_652) );
BUFx2_ASAP7_75t_R g654 ( .A(n_655), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_664), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_661), .A2(n_663), .B1(n_982), .B2(n_983), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_669), .B2(n_670), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g755 ( .A(n_668), .Y(n_755) );
INVx3_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx4_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g863 ( .A(n_680), .Y(n_863) );
BUFx2_ASAP7_75t_L g944 ( .A(n_680), .Y(n_944) );
INVx1_ASAP7_75t_L g1021 ( .A(n_685), .Y(n_1021) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_804), .B1(n_1018), .B2(n_1019), .Y(n_685) );
INVx1_ASAP7_75t_L g1018 ( .A(n_686), .Y(n_1018) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_741), .B1(n_742), .B2(n_803), .Y(n_686) );
INVx1_ASAP7_75t_SL g803 ( .A(n_687), .Y(n_803) );
BUFx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI22xp5_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_690), .B1(n_711), .B2(n_740), .Y(n_688) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
XNOR2xp5_ASAP7_75t_L g772 ( .A(n_691), .B(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
XOR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_710), .Y(n_692) );
NAND4xp75_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .C(n_703), .D(n_707), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
OA211x2_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B(n_700), .C(n_702), .Y(n_697) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g740 ( .A(n_711), .Y(n_740) );
INVx2_ASAP7_75t_L g739 ( .A(n_712), .Y(n_739) );
AND2x2_ASAP7_75t_SL g712 ( .A(n_713), .B(n_726), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_717), .C(n_722), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g890 ( .A1(n_718), .A2(n_891), .B(n_892), .Y(n_890) );
OAI22xp5_ASAP7_75t_SL g788 ( .A1(n_725), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_725), .A2(n_867), .B1(n_868), .B2(n_869), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_732), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_736), .Y(n_732) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_772), .B1(n_801), .B2(n_802), .Y(n_743) );
INVx2_ASAP7_75t_L g801 ( .A(n_744), .Y(n_801) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_746), .B(n_760), .Y(n_745) );
NOR3xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_753), .C(n_757), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_750), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_767), .Y(n_760) );
OAI21xp5_ASAP7_75t_SL g761 ( .A1(n_762), .A2(n_763), .B(n_764), .Y(n_761) );
OAI21xp5_ASAP7_75t_SL g835 ( .A1(n_762), .A2(n_836), .B(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g997 ( .A(n_765), .Y(n_997) );
BUFx4f_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g911 ( .A(n_766), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g802 ( .A(n_772), .Y(n_802) );
XNOR2x1_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
AND2x2_ASAP7_75t_L g775 ( .A(n_776), .B(n_792), .Y(n_775) );
NOR3xp33_ASAP7_75t_L g776 ( .A(n_777), .B(n_784), .C(n_788), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_782), .B2(n_783), .Y(n_777) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
AND4x1_ASAP7_75t_L g792 ( .A(n_793), .B(n_795), .C(n_799), .D(n_800), .Y(n_792) );
INVx3_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g1019 ( .A(n_804), .Y(n_1019) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_882), .B1(n_1016), .B2(n_1017), .Y(n_804) );
INVx2_ASAP7_75t_SL g1016 ( .A(n_805), .Y(n_1016) );
XNOR2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_853), .Y(n_805) );
OAI22x1_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .B1(n_832), .B2(n_852), .Y(n_806) );
INVx3_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
XOR2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_831), .Y(n_808) );
NAND2xp5_ASAP7_75t_SL g809 ( .A(n_810), .B(n_821), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_816), .Y(n_810) );
OAI21xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_813), .B(n_815), .Y(n_811) );
OAI221xp5_ASAP7_75t_L g909 ( .A1(n_813), .A2(n_910), .B1(n_911), .B2(n_912), .C(n_913), .Y(n_909) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_SL g995 ( .A(n_814), .Y(n_995) );
NAND3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .C(n_820), .Y(n_816) );
NOR2x1_ASAP7_75t_L g821 ( .A(n_822), .B(n_826), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_825), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_830), .A2(n_985), .B1(n_986), .B2(n_987), .Y(n_984) );
INVx3_ASAP7_75t_L g852 ( .A(n_832), .Y(n_852) );
XOR2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_851), .Y(n_832) );
NAND2x1_ASAP7_75t_SL g833 ( .A(n_834), .B(n_843), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_835), .B(n_838), .Y(n_834) );
NAND3xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_841), .C(n_842), .Y(n_838) );
BUFx2_ASAP7_75t_L g967 ( .A(n_840), .Y(n_967) );
NOR2x1_ASAP7_75t_L g843 ( .A(n_844), .B(n_848), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
BUFx2_ASAP7_75t_L g988 ( .A(n_847), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
INVx2_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
AND2x2_ASAP7_75t_SL g855 ( .A(n_856), .B(n_870), .Y(n_855) );
NOR3xp33_ASAP7_75t_L g856 ( .A(n_857), .B(n_861), .C(n_866), .Y(n_856) );
OAI222xp33_ASAP7_75t_L g993 ( .A1(n_863), .A2(n_994), .B1(n_995), .B2(n_996), .C1(n_997), .C2(n_998), .Y(n_993) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_877), .Y(n_870) );
NAND2xp5_ASAP7_75t_SL g871 ( .A(n_872), .B(n_874), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_878), .B(n_879), .Y(n_877) );
INVx1_ASAP7_75t_L g1017 ( .A(n_882), .Y(n_1017) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_883), .A2(n_884), .B1(n_932), .B2(n_1015), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
OAI22xp5_ASAP7_75t_SL g884 ( .A1(n_885), .A2(n_886), .B1(n_905), .B2(n_931), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
XOR2x2_ASAP7_75t_L g887 ( .A(n_888), .B(n_904), .Y(n_887) );
NAND3x1_ASAP7_75t_L g888 ( .A(n_889), .B(n_897), .C(n_901), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_890), .B(n_893), .Y(n_889) );
NAND3xp33_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .C(n_896), .Y(n_893) );
AND2x2_ASAP7_75t_L g897 ( .A(n_898), .B(n_900), .Y(n_897) );
AND2x2_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
INVx1_ASAP7_75t_L g931 ( .A(n_905), .Y(n_931) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
XOR2x2_ASAP7_75t_L g906 ( .A(n_907), .B(n_930), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_908), .B(n_921), .Y(n_907) );
NOR3xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_914), .C(n_917), .Y(n_908) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_926), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_923), .B(n_925), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_927), .B(n_928), .Y(n_926) );
INVx1_ASAP7_75t_L g1015 ( .A(n_932), .Y(n_1015) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_958), .B1(n_1013), .B2(n_1014), .Y(n_932) );
INVx1_ASAP7_75t_L g1013 ( .A(n_933), .Y(n_1013) );
XOR2x2_ASAP7_75t_L g933 ( .A(n_934), .B(n_957), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_935), .B(n_949), .Y(n_934) );
NOR3xp33_ASAP7_75t_L g935 ( .A(n_936), .B(n_940), .C(n_945), .Y(n_935) );
OAI21xp33_ASAP7_75t_L g940 ( .A1(n_941), .A2(n_942), .B(n_943), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g949 ( .A(n_950), .B(n_954), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_951), .B(n_952), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_955), .B(n_956), .Y(n_954) );
INVx1_ASAP7_75t_L g1014 ( .A(n_958), .Y(n_1014) );
AOI22xp5_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_989), .B1(n_1011), .B2(n_1012), .Y(n_958) );
INVx2_ASAP7_75t_L g1012 ( .A(n_959), .Y(n_1012) );
XNOR2x1_ASAP7_75t_L g959 ( .A(n_960), .B(n_961), .Y(n_959) );
AND2x2_ASAP7_75t_L g961 ( .A(n_962), .B(n_974), .Y(n_961) );
OAI211xp5_ASAP7_75t_L g963 ( .A1(n_964), .A2(n_965), .B(n_966), .C(n_968), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_970), .A2(n_971), .B1(n_972), .B2(n_973), .Y(n_969) );
NOR3xp33_ASAP7_75t_L g974 ( .A(n_975), .B(n_981), .C(n_984), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_979), .Y(n_975) );
INVx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g1011 ( .A(n_989), .Y(n_1011) );
INVx1_ASAP7_75t_SL g1010 ( .A(n_991), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_992), .B(n_1003), .Y(n_991) );
NOR2x1_ASAP7_75t_L g992 ( .A(n_993), .B(n_999), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1001), .Y(n_999) );
NOR2xp33_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1007), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1006), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1009), .Y(n_1007) );
INVx1_ASAP7_75t_SL g1022 ( .A(n_1023), .Y(n_1022) );
NOR2x1_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1028), .Y(n_1023) );
OR2x2_ASAP7_75t_SL g1081 ( .A(n_1024), .B(n_1029), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1027), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
HB1xp67_ASAP7_75t_L g1057 ( .A(n_1026), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1026), .B(n_1060), .Y(n_1063) );
CKINVDCx16_ASAP7_75t_R g1060 ( .A(n_1027), .Y(n_1060) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_1029), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1031), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1034), .Y(n_1032) );
OAI322xp33_ASAP7_75t_L g1035 ( .A1(n_1036), .A2(n_1057), .A3(n_1058), .B1(n_1061), .B2(n_1064), .C1(n_1065), .C2(n_1079), .Y(n_1035) );
INVx2_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1049), .Y(n_1038) );
NOR3xp33_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1043), .C(n_1046), .Y(n_1039) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1054), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1052), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1056), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
CKINVDCx16_ASAP7_75t_R g1061 ( .A(n_1062), .Y(n_1061) );
NAND4xp75_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1070), .C(n_1075), .D(n_1078), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1069), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1074), .Y(n_1070) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
AND2x2_ASAP7_75t_SL g1075 ( .A(n_1076), .B(n_1077), .Y(n_1075) );
CKINVDCx20_ASAP7_75t_R g1079 ( .A(n_1080), .Y(n_1079) );
CKINVDCx20_ASAP7_75t_R g1080 ( .A(n_1081), .Y(n_1080) );
endmodule