module fake_netlist_1_6477_n_704 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_704);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_704;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_72), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_4), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_28), .Y(n_84) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_64), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_54), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_65), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_0), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_30), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_13), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_62), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_77), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_6), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_32), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_29), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_36), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_0), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_26), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_22), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_76), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_15), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_4), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_73), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_61), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_39), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_37), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_57), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_27), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_60), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_23), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_17), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_50), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_24), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_21), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_31), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_21), .Y(n_116) );
INVxp33_ASAP7_75t_SL g117 ( .A(n_22), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_75), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_1), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_45), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_79), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_15), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_59), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_53), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_7), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_33), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_41), .Y(n_127) );
INVxp67_ASAP7_75t_SL g128 ( .A(n_78), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_46), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_42), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_82), .Y(n_131) );
XNOR2xp5_ASAP7_75t_L g132 ( .A(n_117), .B(n_1), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_84), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_129), .B(n_2), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_95), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_84), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_87), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_83), .B(n_2), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_95), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_95), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_90), .B(n_3), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_92), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_90), .B(n_3), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_85), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_92), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_101), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_96), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_96), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_101), .B(n_5), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_98), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_83), .B(n_5), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_98), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_93), .B(n_6), .Y(n_155) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_103), .A2(n_44), .B(n_80), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_96), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_103), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_119), .B(n_7), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_104), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_93), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_130), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_104), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_97), .B(n_99), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_105), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_97), .B(n_8), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_105), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_108), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_99), .B(n_8), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_108), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_156), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_146), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_141), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_164), .B(n_122), .Y(n_175) );
INVx2_ASAP7_75t_SL g176 ( .A(n_161), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
OR2x2_ASAP7_75t_L g178 ( .A(n_148), .B(n_114), .Y(n_178) );
OR2x2_ASAP7_75t_SL g179 ( .A(n_161), .B(n_116), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_156), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_162), .B(n_125), .Y(n_182) );
INVx1_ASAP7_75t_SL g183 ( .A(n_148), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_142), .Y(n_184) );
AO22x2_ASAP7_75t_L g185 ( .A1(n_145), .A2(n_109), .B1(n_110), .B2(n_126), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_164), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_162), .B(n_113), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_164), .B(n_102), .Y(n_188) );
INVxp67_ASAP7_75t_L g189 ( .A(n_145), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_136), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_131), .B(n_133), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_142), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_136), .Y(n_193) );
NOR2x1p5_ASAP7_75t_L g194 ( .A(n_145), .B(n_111), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_162), .B(n_91), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_136), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_142), .Y(n_197) );
NAND2xp33_ASAP7_75t_L g198 ( .A(n_131), .B(n_118), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_151), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_149), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_133), .B(n_134), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_162), .B(n_86), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_134), .B(n_102), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_136), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_137), .B(n_112), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_136), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_136), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_151), .B(n_116), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_149), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_149), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_137), .B(n_107), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_150), .Y(n_213) );
BUFx8_ASAP7_75t_SL g214 ( .A(n_151), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_138), .B(n_122), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_150), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_157), .Y(n_217) );
OAI221xp5_ASAP7_75t_L g218 ( .A1(n_140), .A2(n_88), .B1(n_128), .B2(n_89), .C(n_94), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_157), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_156), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_138), .Y(n_222) );
INVx1_ASAP7_75t_SL g223 ( .A(n_143), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_143), .B(n_115), .Y(n_224) );
BUFx2_ASAP7_75t_L g225 ( .A(n_153), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_139), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_156), .Y(n_227) );
INVx5_ASAP7_75t_L g228 ( .A(n_153), .Y(n_228) );
INVx1_ASAP7_75t_SL g229 ( .A(n_153), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_139), .B(n_109), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_144), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_144), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_147), .B(n_110), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_156), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_192), .Y(n_235) );
INVxp67_ASAP7_75t_SL g236 ( .A(n_186), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_222), .Y(n_237) );
BUFx4f_ASAP7_75t_L g238 ( .A(n_191), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_222), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_176), .B(n_170), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_183), .Y(n_241) );
AND3x2_ASAP7_75t_SL g242 ( .A(n_185), .B(n_106), .C(n_120), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_176), .B(n_135), .Y(n_243) );
AOI211xp5_ASAP7_75t_L g244 ( .A1(n_218), .A2(n_132), .B(n_159), .C(n_140), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_186), .Y(n_245) );
NOR2xp33_ASAP7_75t_R g246 ( .A(n_172), .B(n_100), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_227), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_222), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_227), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_182), .B(n_170), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_222), .Y(n_251) );
BUFx3_ASAP7_75t_L g252 ( .A(n_186), .Y(n_252) );
INVx6_ASAP7_75t_L g253 ( .A(n_228), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_228), .B(n_152), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_231), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_231), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_192), .Y(n_257) );
BUFx4f_ASAP7_75t_L g258 ( .A(n_191), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_231), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_192), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_227), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_185), .A2(n_152), .B1(n_168), .B2(n_167), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_231), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_226), .A2(n_147), .B(n_168), .C(n_167), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_228), .B(n_165), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_185), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_191), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_212), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_223), .B(n_132), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_212), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_214), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_228), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_229), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_212), .Y(n_274) );
CKINVDCx11_ASAP7_75t_R g275 ( .A(n_175), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_228), .B(n_154), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_177), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_191), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_225), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_227), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_178), .B(n_154), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_201), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_177), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_201), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_201), .B(n_228), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_201), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_173), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_225), .B(n_158), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_175), .B(n_169), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_173), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_174), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_174), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_224), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_189), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_177), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_180), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_190), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_180), .Y(n_298) );
NAND2x1_ASAP7_75t_L g299 ( .A(n_226), .B(n_158), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_175), .B(n_169), .Y(n_300) );
O2A1O1Ixp5_ASAP7_75t_L g301 ( .A1(n_171), .A2(n_165), .B(n_163), .C(n_160), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_175), .B(n_163), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_197), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_241), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_267), .Y(n_305) );
BUFx12f_ASAP7_75t_L g306 ( .A(n_271), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_262), .A2(n_185), .B1(n_179), .B2(n_233), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_266), .A2(n_185), .B1(n_238), .B2(n_258), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_266), .A2(n_245), .B1(n_252), .B2(n_194), .Y(n_309) );
AOI22xp33_ASAP7_75t_SL g310 ( .A1(n_293), .A2(n_224), .B1(n_208), .B2(n_188), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_241), .B(n_178), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_273), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_244), .A2(n_199), .B1(n_194), .B2(n_208), .Y(n_313) );
AND3x1_ASAP7_75t_SL g314 ( .A(n_246), .B(n_179), .C(n_124), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_238), .A2(n_233), .B1(n_203), .B2(n_215), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_267), .Y(n_316) );
INVx4_ASAP7_75t_L g317 ( .A(n_238), .Y(n_317) );
OR2x6_ASAP7_75t_SL g318 ( .A(n_271), .B(n_155), .Y(n_318) );
BUFx12f_ASAP7_75t_L g319 ( .A(n_275), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_288), .B(n_188), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_SL g321 ( .A1(n_264), .A2(n_234), .B(n_221), .C(n_232), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_245), .A2(n_215), .B1(n_203), .B2(n_233), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_299), .A2(n_221), .B(n_234), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_235), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_245), .A2(n_215), .B1(n_203), .B2(n_233), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_278), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_258), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_244), .A2(n_198), .B1(n_202), .B2(n_203), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_278), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_235), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_258), .A2(n_215), .B1(n_232), .B2(n_230), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_282), .Y(n_332) );
INVx4_ASAP7_75t_L g333 ( .A(n_252), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_282), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_288), .B(n_205), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_269), .B(n_155), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_281), .B(n_211), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_279), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_SL g339 ( .A1(n_299), .A2(n_234), .B(n_221), .C(n_210), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_284), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_294), .B(n_187), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_269), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_236), .B(n_197), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_284), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_286), .Y(n_345) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_242), .Y(n_346) );
NOR2xp67_ASAP7_75t_L g347 ( .A(n_243), .B(n_184), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_240), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_289), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_286), .B(n_166), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_302), .B(n_166), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_250), .B(n_210), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_254), .Y(n_353) );
NAND2xp33_ASAP7_75t_L g354 ( .A(n_247), .B(n_227), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_247), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_287), .A2(n_160), .B1(n_220), .B2(n_219), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_308), .A2(n_300), .B1(n_303), .B2(n_298), .Y(n_357) );
OAI222xp33_ASAP7_75t_L g358 ( .A1(n_308), .A2(n_242), .B1(n_298), .B2(n_296), .C1(n_292), .C2(n_291), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_304), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_307), .A2(n_303), .B1(n_296), .B2(n_292), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_348), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_310), .A2(n_195), .B1(n_290), .B2(n_291), .C(n_287), .Y(n_362) );
OAI21x1_ASAP7_75t_L g363 ( .A1(n_323), .A2(n_301), .B(n_237), .Y(n_363) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_346), .A2(n_242), .B1(n_253), .B2(n_290), .Y(n_364) );
NAND2x1_ASAP7_75t_L g365 ( .A(n_317), .B(n_235), .Y(n_365) );
O2A1O1Ixp33_ASAP7_75t_SL g366 ( .A1(n_356), .A2(n_123), .B(n_121), .C(n_124), .Y(n_366) );
O2A1O1Ixp33_ASAP7_75t_SL g367 ( .A1(n_356), .A2(n_121), .B(n_123), .C(n_126), .Y(n_367) );
CKINVDCx6p67_ASAP7_75t_R g368 ( .A(n_319), .Y(n_368) );
AND2x4_ASAP7_75t_SL g369 ( .A(n_317), .B(n_320), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_305), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_333), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_320), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_315), .A2(n_260), .B1(n_235), .B2(n_257), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_336), .B(n_313), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_310), .B(n_265), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_342), .A2(n_285), .B1(n_276), .B2(n_200), .C(n_220), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_337), .B(n_257), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_L g378 ( .A1(n_337), .A2(n_200), .B(n_209), .C(n_213), .Y(n_378) );
AO31x2_ASAP7_75t_L g379 ( .A1(n_323), .A2(n_171), .A3(n_181), .B(n_216), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_324), .A2(n_251), .B(n_237), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g381 ( .A1(n_328), .A2(n_263), .B(n_239), .Y(n_381) );
OR2x6_ASAP7_75t_L g382 ( .A(n_315), .B(n_272), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_311), .B(n_272), .Y(n_383) );
BUFx8_ASAP7_75t_L g384 ( .A(n_306), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_339), .A2(n_247), .B(n_261), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_335), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_307), .A2(n_251), .B1(n_239), .B2(n_255), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g388 ( .A1(n_312), .A2(n_253), .B1(n_257), .B2(n_260), .Y(n_388) );
OAI211xp5_ASAP7_75t_L g389 ( .A1(n_374), .A2(n_309), .B(n_312), .C(n_341), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_357), .A2(n_331), .B1(n_322), .B2(n_325), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_357), .A2(n_331), .B1(n_352), .B2(n_350), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_374), .A2(n_335), .B1(n_338), .B2(n_350), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_360), .A2(n_352), .B1(n_350), .B2(n_351), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_382), .Y(n_394) );
AOI21xp33_ASAP7_75t_L g395 ( .A1(n_362), .A2(n_333), .B(n_327), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_361), .B(n_372), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_364), .A2(n_349), .B1(n_353), .B2(n_347), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_370), .Y(n_398) );
OAI211xp5_ASAP7_75t_SL g399 ( .A1(n_386), .A2(n_314), .B(n_318), .C(n_115), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_375), .A2(n_326), .B1(n_329), .B2(n_345), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_377), .Y(n_401) );
OAI21xp5_ASAP7_75t_L g402 ( .A1(n_378), .A2(n_343), .B(n_321), .Y(n_402) );
OR2x6_ASAP7_75t_L g403 ( .A(n_382), .B(n_373), .Y(n_403) );
AOI222xp33_ASAP7_75t_L g404 ( .A1(n_358), .A2(n_360), .B1(n_369), .B2(n_384), .C1(n_387), .C2(n_359), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_383), .Y(n_405) );
OAI211xp5_ASAP7_75t_L g406 ( .A1(n_366), .A2(n_316), .B(n_344), .C(n_340), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_379), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_387), .A2(n_334), .B1(n_332), .B2(n_219), .Y(n_408) );
AOI21x1_ASAP7_75t_L g409 ( .A1(n_385), .A2(n_190), .B(n_193), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_384), .Y(n_410) );
AOI211x1_ASAP7_75t_L g411 ( .A1(n_381), .A2(n_209), .B(n_213), .C(n_216), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_382), .A2(n_253), .B1(n_256), .B2(n_255), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_379), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_378), .A2(n_257), .B1(n_260), .B2(n_268), .Y(n_414) );
BUFx2_ASAP7_75t_R g415 ( .A(n_368), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_379), .Y(n_416) );
AOI222xp33_ASAP7_75t_L g417 ( .A1(n_393), .A2(n_369), .B1(n_376), .B2(n_217), .C1(n_371), .C2(n_171), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_398), .B(n_379), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_405), .B(n_371), .Y(n_419) );
AOI33xp33_ASAP7_75t_L g420 ( .A1(n_392), .A2(n_367), .A3(n_366), .B1(n_106), .B2(n_120), .B3(n_127), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_407), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g422 ( .A1(n_391), .A2(n_403), .B1(n_390), .B2(n_394), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_398), .B(n_217), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_404), .B(n_184), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_404), .A2(n_388), .B1(n_184), .B2(n_330), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_396), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_401), .B(n_184), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_401), .B(n_363), .Y(n_428) );
INVxp67_ASAP7_75t_L g429 ( .A(n_407), .Y(n_429) );
OAI211xp5_ASAP7_75t_L g430 ( .A1(n_399), .A2(n_367), .B(n_106), .C(n_127), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_394), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g432 ( .A1(n_403), .A2(n_365), .B1(n_171), .B2(n_181), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_403), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_413), .Y(n_434) );
OAI22xp33_ASAP7_75t_L g435 ( .A1(n_403), .A2(n_181), .B1(n_253), .B2(n_270), .Y(n_435) );
BUFx2_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_389), .A2(n_127), .B1(n_120), .B2(n_256), .C(n_263), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_411), .B(n_181), .C(n_227), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_407), .Y(n_439) );
OR2x2_ASAP7_75t_SL g440 ( .A(n_416), .B(n_9), .Y(n_440) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_397), .B(n_9), .C(n_10), .D(n_11), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_400), .A2(n_259), .B1(n_248), .B2(n_268), .C(n_260), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_395), .A2(n_268), .B1(n_270), .B2(n_380), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_416), .A2(n_268), .B1(n_270), .B2(n_274), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_406), .A2(n_270), .B1(n_274), .B2(n_259), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_416), .B(n_10), .Y(n_446) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_413), .A2(n_190), .B(n_206), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_411), .B(n_248), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_409), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
OAI22xp33_ASAP7_75t_L g451 ( .A1(n_408), .A2(n_355), .B1(n_280), .B2(n_261), .Y(n_451) );
AOI221xp5_ASAP7_75t_SL g452 ( .A1(n_402), .A2(n_354), .B1(n_193), .B2(n_196), .C(n_204), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_408), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_418), .B(n_412), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_434), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_421), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_418), .B(n_11), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_453), .B(n_414), .Y(n_458) );
OAI31xp33_ASAP7_75t_L g459 ( .A1(n_441), .A2(n_415), .A3(n_13), .B(n_14), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_453), .B(n_280), .Y(n_460) );
OAI22xp33_ASAP7_75t_L g461 ( .A1(n_441), .A2(n_410), .B1(n_355), .B2(n_280), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_421), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_429), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_446), .B(n_12), .Y(n_464) );
OR2x2_ASAP7_75t_SL g465 ( .A(n_439), .B(n_410), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_428), .B(n_247), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_434), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_439), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_434), .Y(n_469) );
AOI31xp33_ASAP7_75t_L g470 ( .A1(n_433), .A2(n_12), .A3(n_14), .B(n_16), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_440), .A2(n_355), .B1(n_280), .B2(n_261), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_428), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_449), .Y(n_473) );
INVx4_ASAP7_75t_L g474 ( .A(n_436), .Y(n_474) );
OAI31xp33_ASAP7_75t_L g475 ( .A1(n_430), .A2(n_16), .A3(n_17), .B(n_18), .Y(n_475) );
OAI33xp33_ASAP7_75t_L g476 ( .A1(n_422), .A2(n_18), .A3(n_19), .B1(n_20), .B2(n_207), .B3(n_206), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_449), .Y(n_477) );
INVx4_ASAP7_75t_L g478 ( .A(n_436), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_426), .B(n_19), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_429), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_447), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_446), .Y(n_482) );
BUFx3_ASAP7_75t_L g483 ( .A(n_431), .Y(n_483) );
OAI221xp5_ASAP7_75t_SL g484 ( .A1(n_420), .A2(n_20), .B1(n_207), .B2(n_206), .C(n_204), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_424), .A2(n_193), .B1(n_196), .B2(n_204), .C(n_207), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_433), .B(n_196), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_419), .Y(n_487) );
AOI33xp33_ASAP7_75t_L g488 ( .A1(n_424), .A2(n_297), .A3(n_295), .B1(n_283), .B2(n_277), .B3(n_40), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_433), .B(n_25), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_449), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_450), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_450), .B(n_34), .Y(n_492) );
AOI221xp5_ASAP7_75t_L g493 ( .A1(n_437), .A2(n_247), .B1(n_249), .B2(n_261), .C(n_280), .Y(n_493) );
OAI33xp33_ASAP7_75t_L g494 ( .A1(n_419), .A2(n_35), .A3(n_38), .B1(n_43), .B2(n_47), .B3(n_48), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_431), .Y(n_495) );
AND2x4_ASAP7_75t_SL g496 ( .A(n_423), .B(n_261), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_431), .B(n_249), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_450), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_423), .B(n_49), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_448), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_427), .B(n_51), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_448), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_427), .B(n_52), .Y(n_503) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_432), .A2(n_297), .B(n_295), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_437), .B(n_249), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_417), .A2(n_249), .B1(n_277), .B2(n_283), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_447), .B(n_55), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_461), .B(n_452), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_483), .Y(n_509) );
NAND4xp75_ASAP7_75t_L g510 ( .A(n_459), .B(n_452), .C(n_440), .D(n_442), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_457), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_457), .B(n_417), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_483), .Y(n_513) );
NAND2xp33_ASAP7_75t_L g514 ( .A(n_471), .B(n_425), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_487), .B(n_447), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_472), .B(n_438), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_463), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_457), .B(n_430), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_456), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_454), .B(n_438), .Y(n_520) );
NAND4xp75_ASAP7_75t_L g521 ( .A(n_459), .B(n_442), .C(n_445), .D(n_435), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_463), .B(n_443), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_454), .B(n_444), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_456), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_454), .B(n_445), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_462), .B(n_56), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_487), .B(n_451), .Y(n_527) );
NOR3xp33_ASAP7_75t_L g528 ( .A(n_470), .B(n_58), .C(n_63), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_474), .B(n_66), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_462), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_468), .Y(n_531) );
INVx3_ASAP7_75t_L g532 ( .A(n_481), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_468), .B(n_67), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_480), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_482), .B(n_68), .Y(n_535) );
OAI221xp5_ASAP7_75t_L g536 ( .A1(n_479), .A2(n_249), .B1(n_70), .B2(n_71), .C(n_74), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_480), .B(n_69), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_482), .B(n_81), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_500), .B(n_502), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_455), .B(n_469), .Y(n_540) );
OR2x6_ASAP7_75t_L g541 ( .A(n_471), .B(n_478), .Y(n_541) );
INVxp67_ASAP7_75t_SL g542 ( .A(n_481), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_464), .B(n_500), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_464), .B(n_495), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_455), .B(n_469), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_465), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_467), .B(n_469), .Y(n_547) );
OAI211xp5_ASAP7_75t_SL g548 ( .A1(n_475), .A2(n_488), .B(n_485), .C(n_506), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_467), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_467), .B(n_502), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_465), .Y(n_551) );
NOR2xp67_ASAP7_75t_L g552 ( .A(n_481), .B(n_478), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_458), .B(n_499), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_498), .Y(n_554) );
INVxp67_ASAP7_75t_SL g555 ( .A(n_481), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_498), .B(n_491), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_458), .B(n_499), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_495), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_474), .B(n_478), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_473), .B(n_490), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_473), .B(n_490), .Y(n_561) );
NOR2xp67_ASAP7_75t_SL g562 ( .A(n_507), .B(n_489), .Y(n_562) );
OAI21xp33_ASAP7_75t_L g563 ( .A1(n_470), .A2(n_507), .B(n_484), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_476), .A2(n_484), .B1(n_475), .B2(n_494), .C(n_485), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_473), .B(n_491), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_474), .B(n_478), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_534), .B(n_491), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_544), .B(n_511), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_519), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_524), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_546), .B(n_474), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_517), .B(n_490), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_552), .B(n_496), .Y(n_573) );
INVxp67_ASAP7_75t_SL g574 ( .A(n_542), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_539), .B(n_477), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_563), .B(n_507), .Y(n_576) );
OAI21xp5_ASAP7_75t_L g577 ( .A1(n_564), .A2(n_493), .B(n_489), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_560), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_508), .A2(n_493), .B(n_494), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_509), .Y(n_580) );
BUFx2_ASAP7_75t_L g581 ( .A(n_509), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_561), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_520), .B(n_496), .Y(n_583) );
AND2x4_ASAP7_75t_L g584 ( .A(n_541), .B(n_477), .Y(n_584) );
NOR2xp67_ASAP7_75t_SL g585 ( .A(n_537), .B(n_503), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_530), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_510), .A2(n_505), .B(n_492), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_531), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_558), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_554), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_539), .B(n_477), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_543), .B(n_466), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_550), .B(n_460), .Y(n_593) );
NOR2x1_ASAP7_75t_L g594 ( .A(n_529), .B(n_503), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_559), .B(n_466), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_541), .B(n_486), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_558), .Y(n_597) );
NOR2x1_ASAP7_75t_L g598 ( .A(n_529), .B(n_501), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_559), .B(n_460), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_550), .Y(n_600) );
BUFx5_ASAP7_75t_L g601 ( .A(n_529), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_513), .B(n_486), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_556), .B(n_504), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_566), .B(n_497), .Y(n_604) );
OAI31xp33_ASAP7_75t_SL g605 ( .A1(n_551), .A2(n_501), .A3(n_476), .B(n_504), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_514), .A2(n_504), .B1(n_505), .B2(n_497), .Y(n_606) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_528), .B(n_504), .C(n_514), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_515), .B(n_557), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_523), .B(n_525), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_540), .B(n_547), .Y(n_610) );
AND2x4_ASAP7_75t_L g611 ( .A(n_541), .B(n_532), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_540), .B(n_547), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_545), .B(n_565), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_523), .B(n_525), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_569), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_570), .Y(n_616) );
XOR2x2_ASAP7_75t_L g617 ( .A(n_594), .B(n_512), .Y(n_617) );
AND2x4_ASAP7_75t_SL g618 ( .A(n_573), .B(n_541), .Y(n_618) );
INVx3_ASAP7_75t_L g619 ( .A(n_573), .Y(n_619) );
INVxp67_ASAP7_75t_L g620 ( .A(n_597), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_598), .A2(n_518), .B1(n_537), .B2(n_555), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_586), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_588), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_605), .A2(n_508), .B(n_548), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_590), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_609), .B(n_516), .Y(n_626) );
XNOR2x1_ASAP7_75t_L g627 ( .A(n_614), .B(n_521), .Y(n_627) );
A2O1A1Ixp33_ASAP7_75t_SL g628 ( .A1(n_577), .A2(n_536), .B(n_562), .C(n_532), .Y(n_628) );
NOR2xp33_ASAP7_75t_R g629 ( .A(n_580), .B(n_553), .Y(n_629) );
AOI21xp33_ASAP7_75t_SL g630 ( .A1(n_576), .A2(n_522), .B(n_532), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_607), .B(n_522), .C(n_516), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_568), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_600), .B(n_516), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_610), .Y(n_634) );
NOR2x1_ASAP7_75t_L g635 ( .A(n_581), .B(n_526), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_613), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_604), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_608), .B(n_549), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_613), .Y(n_639) );
AND2x2_ASAP7_75t_SL g640 ( .A(n_611), .B(n_526), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_610), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_612), .B(n_527), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_592), .B(n_582), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_578), .B(n_538), .Y(n_644) );
XOR2x2_ASAP7_75t_L g645 ( .A(n_587), .B(n_533), .Y(n_645) );
XNOR2xp5_ASAP7_75t_L g646 ( .A(n_612), .B(n_535), .Y(n_646) );
XOR2xp5_ASAP7_75t_L g647 ( .A(n_595), .B(n_538), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_575), .Y(n_648) );
AOI21xp33_ASAP7_75t_L g649 ( .A1(n_571), .A2(n_535), .B(n_533), .Y(n_649) );
NOR4xp25_ASAP7_75t_L g650 ( .A(n_587), .B(n_577), .C(n_589), .D(n_572), .Y(n_650) );
AOI221x1_ASAP7_75t_L g651 ( .A1(n_579), .A2(n_611), .B1(n_572), .B2(n_596), .C(n_591), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_589), .B(n_591), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_593), .B(n_599), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_585), .B(n_596), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_593), .B(n_603), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_567), .Y(n_656) );
AOI31xp33_ASAP7_75t_L g657 ( .A1(n_579), .A2(n_574), .A3(n_606), .B(n_584), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_567), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_603), .A2(n_584), .B(n_602), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_601), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_583), .B(n_601), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_601), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_601), .A2(n_576), .B1(n_563), .B2(n_594), .Y(n_663) );
INVxp67_ASAP7_75t_L g664 ( .A(n_601), .Y(n_664) );
NAND3xp33_ASAP7_75t_L g665 ( .A(n_605), .B(n_607), .C(n_589), .Y(n_665) );
OAI21xp33_ASAP7_75t_L g666 ( .A1(n_605), .A2(n_607), .B(n_576), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_569), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_581), .Y(n_668) );
AOI211xp5_ASAP7_75t_L g669 ( .A1(n_624), .A2(n_650), .B(n_666), .C(n_665), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_627), .A2(n_617), .B1(n_663), .B2(n_621), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_619), .B(n_637), .Y(n_671) );
AOI321xp33_ASAP7_75t_L g672 ( .A1(n_621), .A2(n_630), .A3(n_654), .B1(n_659), .B2(n_635), .C(n_652), .Y(n_672) );
XNOR2x2_ASAP7_75t_L g673 ( .A(n_645), .B(n_631), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_668), .B(n_620), .Y(n_674) );
OAI21xp5_ASAP7_75t_L g675 ( .A1(n_651), .A2(n_657), .B(n_628), .Y(n_675) );
XOR2x2_ASAP7_75t_L g676 ( .A(n_646), .B(n_647), .Y(n_676) );
OAI211xp5_ASAP7_75t_L g677 ( .A1(n_629), .A2(n_654), .B(n_619), .C(n_661), .Y(n_677) );
NAND2x1_ASAP7_75t_L g678 ( .A(n_661), .B(n_652), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_656), .Y(n_679) );
XNOR2xp5_ASAP7_75t_L g680 ( .A(n_640), .B(n_618), .Y(n_680) );
AO22x2_ASAP7_75t_L g681 ( .A1(n_632), .A2(n_664), .B1(n_667), .B2(n_622), .Y(n_681) );
AOI211xp5_ASAP7_75t_SL g682 ( .A1(n_669), .A2(n_649), .B(n_662), .C(n_626), .Y(n_682) );
OAI211xp5_ASAP7_75t_SL g683 ( .A1(n_669), .A2(n_655), .B(n_642), .C(n_633), .Y(n_683) );
OAI221xp5_ASAP7_75t_R g684 ( .A1(n_670), .A2(n_653), .B1(n_636), .B2(n_639), .C(n_641), .Y(n_684) );
OAI221xp5_ASAP7_75t_SL g685 ( .A1(n_670), .A2(n_633), .B1(n_634), .B2(n_644), .C(n_660), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_681), .B(n_648), .Y(n_686) );
AOI211xp5_ASAP7_75t_L g687 ( .A1(n_675), .A2(n_660), .B(n_616), .C(n_623), .Y(n_687) );
OAI211xp5_ASAP7_75t_L g688 ( .A1(n_672), .A2(n_615), .B(n_625), .C(n_638), .Y(n_688) );
NOR4xp25_ASAP7_75t_L g689 ( .A(n_673), .B(n_643), .C(n_658), .D(n_638), .Y(n_689) );
NOR2x1p5_ASAP7_75t_L g690 ( .A(n_686), .B(n_678), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_686), .Y(n_691) );
AO22x2_ASAP7_75t_L g692 ( .A1(n_688), .A2(n_677), .B1(n_671), .B2(n_679), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_684), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_683), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_691), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_691), .Y(n_696) );
NAND5xp2_ASAP7_75t_L g697 ( .A(n_694), .B(n_682), .C(n_687), .D(n_685), .E(n_689), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_696), .Y(n_698) );
XNOR2xp5_ASAP7_75t_L g699 ( .A(n_695), .B(n_676), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_698), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_699), .A2(n_693), .B1(n_695), .B2(n_680), .C(n_692), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_700), .Y(n_702) );
OAI22xp33_ASAP7_75t_L g703 ( .A1(n_702), .A2(n_701), .B1(n_692), .B2(n_697), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_703), .A2(n_690), .B1(n_674), .B2(n_681), .Y(n_704) );
endmodule