module real_jpeg_24201_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_216;
wire n_179;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_73),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_1),
.A2(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

INVx8_ASAP7_75t_SL g34 ( 
.A(n_4),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_5),
.A2(n_60),
.B1(n_69),
.B2(n_70),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_60),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_6),
.A2(n_24),
.B1(n_39),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_45),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_6),
.A2(n_45),
.B1(n_54),
.B2(n_55),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_6),
.A2(n_45),
.B1(n_69),
.B2(n_70),
.Y(n_167)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_7),
.B(n_42),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_7),
.B(n_65),
.C(n_69),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_7),
.A2(n_28),
.B1(n_54),
.B2(n_55),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_7),
.B(n_58),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_7),
.A2(n_85),
.B1(n_89),
.B2(n_167),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_10),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_69),
.B1(n_70),
.B2(n_76),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_11),
.A2(n_69),
.B1(n_70),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_13),
.A2(n_27),
.B1(n_40),
.B2(n_50),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_13),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_13),
.A2(n_50),
.B1(n_69),
.B2(n_70),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_14),
.A2(n_69),
.B1(n_70),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_14),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_84),
.Y(n_112)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_15),
.Y(n_86)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_15),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_104),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_91),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_21),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_46),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_22),
.B(n_48),
.C(n_61),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_28),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_28),
.B(n_68),
.Y(n_174)
);

HAxp5_ASAP7_75t_SL g185 ( 
.A(n_28),
.B(n_36),
.CON(n_185),
.SN(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_29),
.A2(n_33),
.B(n_36),
.C(n_80),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_30),
.B(n_34),
.C(n_35),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_31),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_32),
.A2(n_44),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_38)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_36),
.B1(n_53),
.B2(n_56),
.Y(n_57)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_36),
.B(n_54),
.C(n_56),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_61),
.B2(n_62),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_58),
.B2(n_59),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_49),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_51),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_51),
.A2(n_58),
.B1(n_94),
.B2(n_185),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_53),
.A2(n_55),
.B(n_185),
.C(n_186),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_55),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_55),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_58),
.B(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_59),
.Y(n_125)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_71),
.B(n_74),
.Y(n_62)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_63),
.A2(n_68),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_63),
.A2(n_68),
.B1(n_143),
.B2(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_63),
.A2(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_68),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_70),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_72),
.B(n_77),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_77),
.A2(n_114),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_78),
.B(n_91),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_81),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_87),
.B2(n_89),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_87),
.B(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_85),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_85),
.A2(n_160),
.B1(n_167),
.B2(n_176),
.Y(n_175)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_86),
.Y(n_101)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_86),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_103),
.Y(n_110)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_90),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.C(n_99),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_92),
.B(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_202)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_101),
.A2(n_158),
.B1(n_159),
.B2(n_161),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_117),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_115),
.B2(n_116),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_110),
.A2(n_154),
.B(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_128),
.B2(n_129),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_128),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_212),
.B(n_216),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_197),
.B(n_211),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_181),
.B(n_196),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_155),
.B(n_180),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_144),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_144),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_140),
.B1(n_141),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_151),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_164),
.B(n_179),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_162),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_162),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_173),
.B(n_178),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_174),
.B(n_175),
.Y(n_178)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_195),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_195),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_191),
.C(n_194),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_193),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_199),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_206),
.C(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_215),
.Y(n_216)
);


endmodule