module fake_jpeg_11155_n_570 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_570);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_570;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_58),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_60),
.B(n_69),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_61),
.B(n_72),
.Y(n_135)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_62),
.Y(n_139)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_25),
.B(n_0),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_64),
.B(n_91),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_65),
.B(n_73),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_71),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_27),
.B(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_27),
.B(n_17),
.Y(n_73)
);

NAND2x1_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_0),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_74),
.B(n_2),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_75),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_76),
.B(n_85),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_79),
.Y(n_198)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_82),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_29),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_87),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_42),
.B(n_1),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_92),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_93),
.Y(n_200)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_94),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_96),
.B(n_97),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_31),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_29),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_98),
.B(n_101),
.Y(n_149)
);

AND2x4_ASAP7_75t_L g99 ( 
.A(n_26),
.B(n_54),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_99),
.B(n_123),
.Y(n_187)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_29),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_107),
.Y(n_213)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_109),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_113),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_33),
.B(n_48),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_126),
.Y(n_142)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_39),
.Y(n_116)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_117),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_33),
.B(n_16),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_119),
.B(n_124),
.Y(n_212)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_32),
.Y(n_120)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

BUFx12_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_122),
.Y(n_185)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_38),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_35),
.B(n_16),
.Y(n_124)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_38),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_125),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_35),
.B(n_15),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_58),
.A2(n_115),
.B1(n_66),
.B2(n_67),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_130),
.A2(n_144),
.B1(n_147),
.B2(n_151),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_56),
.B1(n_41),
.B2(n_54),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_136),
.A2(n_138),
.B1(n_150),
.B2(n_190),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_56),
.B1(n_41),
.B2(n_54),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_140),
.B(n_82),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_111),
.A2(n_56),
.B1(n_28),
.B2(n_50),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_102),
.A2(n_50),
.B1(n_28),
.B2(n_55),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_64),
.A2(n_47),
.B1(n_57),
.B2(n_19),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_90),
.A2(n_50),
.B1(n_28),
.B2(n_55),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_64),
.B(n_47),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_153),
.B(n_164),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_59),
.A2(n_57),
.B1(n_19),
.B2(n_21),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_158),
.A2(n_167),
.B1(n_176),
.B2(n_181),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_91),
.B(n_51),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_53),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_165),
.B(n_192),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_83),
.A2(n_53),
.B1(n_51),
.B2(n_46),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_91),
.B(n_45),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_168),
.B(n_170),
.Y(n_221)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_74),
.A2(n_46),
.B(n_45),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_86),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_174),
.B(n_182),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_99),
.A2(n_30),
.B1(n_23),
.B2(n_21),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_70),
.A2(n_30),
.B1(n_23),
.B2(n_5),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_125),
.A2(n_14),
.B(n_13),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_87),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_184),
.A2(n_196),
.B1(n_201),
.B2(n_207),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_88),
.A2(n_95),
.B1(n_89),
.B2(n_93),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_117),
.B(n_14),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_99),
.B(n_13),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_194),
.B(n_206),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_77),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_L g197 ( 
.A1(n_118),
.A2(n_38),
.B1(n_4),
.B2(n_7),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_197),
.A2(n_210),
.B1(n_128),
.B2(n_146),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_106),
.A2(n_3),
.B1(n_8),
.B2(n_10),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_68),
.A2(n_38),
.B1(n_10),
.B2(n_11),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_202),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_121),
.B(n_8),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_103),
.A2(n_8),
.B1(n_80),
.B2(n_107),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_79),
.A2(n_92),
.B1(n_75),
.B2(n_112),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_92),
.B1(n_122),
.B2(n_203),
.Y(n_231)
);

AO22x2_ASAP7_75t_L g210 ( 
.A1(n_123),
.A2(n_82),
.B1(n_86),
.B2(n_62),
.Y(n_210)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_216),
.Y(n_343)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_141),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_218),
.B(n_226),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_220),
.B(n_261),
.Y(n_335)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_149),
.B(n_62),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_225),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_158),
.A2(n_167),
.B1(n_188),
.B2(n_138),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_227),
.A2(n_250),
.B1(n_263),
.B2(n_130),
.Y(n_297)
);

BUFx12f_ASAP7_75t_L g228 ( 
.A(n_154),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_228),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_166),
.B(n_75),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_229),
.B(n_235),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_231),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_205),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_232),
.B(n_233),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_135),
.B(n_122),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_166),
.B(n_140),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_236),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_142),
.B(n_212),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_237),
.B(n_239),
.Y(n_315)
);

AOI21xp33_ASAP7_75t_L g239 ( 
.A1(n_129),
.A2(n_187),
.B(n_192),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_127),
.B(n_172),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_240),
.B(n_245),
.Y(n_340)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_162),
.Y(n_241)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_241),
.Y(n_304)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_195),
.Y(n_242)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_242),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_187),
.B(n_189),
.C(n_214),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_243),
.B(n_282),
.C(n_284),
.Y(n_328)
);

BUFx12_ASAP7_75t_L g244 ( 
.A(n_139),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_244),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_165),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_246),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_186),
.B(n_199),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_248),
.B(n_249),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_185),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_136),
.A2(n_200),
.B1(n_159),
.B2(n_178),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_175),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_251),
.Y(n_337)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_155),
.Y(n_252)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_252),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_137),
.Y(n_253)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_253),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_131),
.B(n_145),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_254),
.Y(n_290)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_134),
.Y(n_255)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_255),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_133),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_256),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_162),
.Y(n_258)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_258),
.Y(n_331)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_210),
.B(n_152),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_270),
.Y(n_296)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_179),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_204),
.Y(n_262)
);

INVx11_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_147),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_264),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_128),
.A2(n_132),
.B1(n_145),
.B2(n_146),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_265),
.A2(n_267),
.B1(n_272),
.B2(n_274),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_177),
.B(n_163),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_266),
.Y(n_325)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_161),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_133),
.B(n_198),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_180),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_143),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_271),
.B(n_286),
.Y(n_342)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_201),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_213),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_178),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_285),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_198),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_144),
.B(n_151),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_279),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_210),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_156),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_132),
.B(n_209),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_280),
.B(n_281),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_210),
.B(n_159),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_200),
.B(n_156),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_215),
.B(n_183),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_283),
.A2(n_287),
.B(n_288),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_169),
.B(n_171),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_169),
.Y(n_285)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_137),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_215),
.B(n_183),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_171),
.B(n_157),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_157),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_289),
.A2(n_258),
.B1(n_217),
.B2(n_236),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_297),
.A2(n_298),
.B1(n_310),
.B2(n_313),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_273),
.A2(n_207),
.B1(n_181),
.B2(n_184),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_235),
.A2(n_196),
.B(n_208),
.C(n_221),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_299),
.B(n_302),
.Y(n_359)
);

A2O1A1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_220),
.A2(n_219),
.B(n_229),
.C(n_260),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_247),
.A2(n_278),
.B1(n_263),
.B2(n_245),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_234),
.A2(n_222),
.B1(n_269),
.B2(n_281),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_311),
.A2(n_320),
.B1(n_322),
.B2(n_332),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_247),
.A2(n_277),
.B1(n_257),
.B2(n_224),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_230),
.B1(n_243),
.B2(n_238),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_317),
.A2(n_319),
.B1(n_339),
.B2(n_297),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_279),
.A2(n_289),
.B1(n_285),
.B2(n_223),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_220),
.A2(n_242),
.B1(n_282),
.B2(n_271),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_282),
.A2(n_246),
.B(n_270),
.C(n_256),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_321),
.A2(n_296),
.B(n_300),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_262),
.A2(n_275),
.B1(n_255),
.B2(n_251),
.Y(n_322)
);

AOI32xp33_ASAP7_75t_L g326 ( 
.A1(n_226),
.A2(n_218),
.A3(n_262),
.B1(n_276),
.B2(n_228),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_326),
.A2(n_228),
.B(n_296),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_329),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_216),
.A2(n_267),
.B1(n_261),
.B2(n_252),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_241),
.B(n_259),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_335),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_286),
.A2(n_274),
.B1(n_253),
.B2(n_244),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_272),
.B(n_244),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_345),
.A2(n_351),
.B(n_368),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_301),
.B(n_325),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_357),
.Y(n_401)
);

INVx5_ASAP7_75t_SL g347 ( 
.A(n_327),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_347),
.Y(n_393)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_295),
.Y(n_348)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_338),
.B(n_228),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_372),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_352),
.A2(n_356),
.B(n_361),
.Y(n_415)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_353),
.Y(n_400)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_307),
.Y(n_355)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_355),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_314),
.A2(n_296),
.B(n_338),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_294),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_307),
.Y(n_358)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_358),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_327),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_360),
.B(n_363),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_313),
.A2(n_300),
.B(n_344),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_364),
.B(n_374),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_340),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_366),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_319),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_301),
.B(n_325),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_367),
.B(n_369),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_299),
.A2(n_344),
.B(n_341),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_318),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_290),
.B(n_315),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_370),
.B(n_373),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_311),
.A2(n_298),
.B(n_302),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_371),
.A2(n_374),
.B(n_381),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_328),
.B(n_317),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_343),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_292),
.A2(n_336),
.B(n_320),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_376),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_332),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_321),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_379),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_290),
.B(n_309),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_378),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_292),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_312),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_380),
.A2(n_305),
.B1(n_295),
.B2(n_304),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_326),
.A2(n_316),
.B(n_342),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_383),
.A2(n_385),
.B(n_386),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_316),
.A2(n_335),
.B1(n_291),
.B2(n_333),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_384),
.A2(n_306),
.B1(n_334),
.B2(n_323),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_342),
.A2(n_335),
.B(n_308),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_342),
.A2(n_329),
.B(n_306),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_291),
.A2(n_333),
.B(n_312),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_387),
.A2(n_359),
.B(n_352),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_390),
.A2(n_409),
.B1(n_410),
.B2(n_366),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_354),
.A2(n_324),
.B1(n_303),
.B2(n_334),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_394),
.A2(n_395),
.B1(n_376),
.B2(n_349),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_354),
.A2(n_324),
.B1(n_303),
.B2(n_337),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_379),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_406),
.Y(n_429)
);

XOR2x2_ASAP7_75t_L g398 ( 
.A(n_356),
.B(n_323),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_398),
.A2(n_405),
.B(n_407),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_330),
.C(n_304),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_403),
.B(n_422),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_347),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_351),
.A2(n_305),
.B(n_331),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g408 ( 
.A(n_359),
.B(n_330),
.CI(n_337),
.CON(n_408),
.SN(n_408)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_413),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_362),
.A2(n_331),
.B1(n_343),
.B2(n_371),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_362),
.A2(n_383),
.B1(n_377),
.B2(n_381),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_347),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_416),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_361),
.A2(n_368),
.B(n_345),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_421),
.A2(n_391),
.B(n_412),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_423),
.A2(n_437),
.B1(n_450),
.B2(n_452),
.Y(n_475)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_411),
.Y(n_424)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_424),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_425),
.A2(n_427),
.B1(n_453),
.B2(n_408),
.Y(n_479)
);

OAI22x1_ASAP7_75t_SL g427 ( 
.A1(n_392),
.A2(n_384),
.B1(n_387),
.B2(n_386),
.Y(n_427)
);

NAND3xp33_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_378),
.C(n_370),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_428),
.B(n_436),
.Y(n_462)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_411),
.Y(n_432)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_432),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_414),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_439),
.Y(n_454)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_399),
.Y(n_435)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_435),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_414),
.Y(n_436)
);

AOI32xp33_ASAP7_75t_L g437 ( 
.A1(n_421),
.A2(n_350),
.A3(n_385),
.B1(n_382),
.B2(n_357),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_438),
.A2(n_391),
.B(n_407),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_401),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_401),
.B(n_363),
.Y(n_440)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_440),
.Y(n_481)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_399),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_441),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_419),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_443),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_353),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_397),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_445),
.Y(n_460)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_400),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_389),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_446),
.Y(n_478)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g455 ( 
.A1(n_447),
.A2(n_449),
.B1(n_451),
.B2(n_406),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_420),
.B(n_369),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_448),
.B(n_420),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_389),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_409),
.A2(n_382),
.B1(n_355),
.B2(n_358),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_402),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_410),
.A2(n_360),
.B1(n_373),
.B2(n_375),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_412),
.A2(n_348),
.B1(n_416),
.B2(n_388),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_455),
.B(n_458),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_422),
.C(n_396),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_465),
.C(n_466),
.Y(n_485)
);

INVx3_ASAP7_75t_SL g458 ( 
.A(n_436),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_459),
.A2(n_463),
.B(n_468),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_438),
.A2(n_392),
.B(n_404),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_434),
.B(n_396),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_427),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_403),
.C(n_415),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_415),
.C(n_388),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_426),
.A2(n_404),
.B(n_408),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_423),
.A2(n_394),
.B1(n_397),
.B2(n_395),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_470),
.B(n_425),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_398),
.C(n_390),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_477),
.C(n_480),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g472 ( 
.A(n_442),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_472),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_474),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_433),
.A2(n_405),
.B1(n_413),
.B2(n_393),
.Y(n_476)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_476),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_431),
.B(n_398),
.C(n_402),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_479),
.A2(n_430),
.B1(n_444),
.B2(n_450),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_453),
.B(n_417),
.C(n_408),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_482),
.B(n_498),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_464),
.B(n_426),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_500),
.Y(n_506)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_454),
.Y(n_488)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_488),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_457),
.B(n_439),
.C(n_424),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_489),
.B(n_502),
.C(n_467),
.Y(n_510)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_460),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_493),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_460),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_495),
.A2(n_481),
.B1(n_480),
.B2(n_456),
.Y(n_511)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_461),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_SL g517 ( 
.A1(n_496),
.A2(n_497),
.B1(n_499),
.B2(n_503),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_465),
.B(n_437),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_454),
.Y(n_499)
);

NAND2xp67_ASAP7_75t_SL g500 ( 
.A(n_462),
.B(n_448),
.Y(n_500)
);

FAx1_ASAP7_75t_SL g501 ( 
.A(n_468),
.B(n_430),
.CI(n_440),
.CON(n_501),
.SN(n_501)
);

OAI322xp33_ASAP7_75t_L g505 ( 
.A1(n_501),
.A2(n_456),
.A3(n_481),
.B1(n_477),
.B2(n_471),
.C1(n_474),
.C2(n_467),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_466),
.B(n_432),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_461),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_483),
.A2(n_459),
.B(n_479),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_504),
.A2(n_518),
.B(n_494),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_505),
.A2(n_491),
.B1(n_501),
.B2(n_502),
.Y(n_523)
);

OA21x2_ASAP7_75t_L g507 ( 
.A1(n_497),
.A2(n_470),
.B(n_463),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_507),
.A2(n_511),
.B1(n_482),
.B2(n_492),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_496),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_508),
.B(n_514),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_510),
.B(n_515),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_484),
.Y(n_512)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_512),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_458),
.C(n_475),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_458),
.C(n_449),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_489),
.B(n_478),
.C(n_469),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_516),
.B(n_520),
.C(n_486),
.Y(n_522)
);

BUFx12f_ASAP7_75t_SL g518 ( 
.A(n_500),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_486),
.B(n_478),
.C(n_469),
.Y(n_520)
);

AO21x1_ASAP7_75t_L g542 ( 
.A1(n_521),
.A2(n_517),
.B(n_509),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_522),
.B(n_529),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_523),
.B(n_506),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_504),
.A2(n_483),
.B(n_494),
.Y(n_524)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_524),
.Y(n_536)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_519),
.Y(n_527)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_527),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_507),
.A2(n_495),
.B1(n_498),
.B2(n_491),
.Y(n_528)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_528),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_487),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_530),
.B(n_507),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_520),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g543 ( 
.A(n_531),
.Y(n_543)
);

NAND4xp25_ASAP7_75t_SL g532 ( 
.A(n_518),
.B(n_443),
.C(n_501),
.D(n_393),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_532),
.B(n_516),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_515),
.B(n_503),
.C(n_452),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_533),
.B(n_510),
.C(n_514),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_535),
.B(n_539),
.Y(n_552)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_537),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_541),
.B(n_532),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_542),
.B(n_545),
.C(n_524),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_SL g545 ( 
.A1(n_525),
.A2(n_512),
.B1(n_511),
.B2(n_473),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_540),
.B(n_526),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_546),
.B(n_548),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_547),
.B(n_541),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_543),
.A2(n_534),
.B(n_522),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_549),
.A2(n_550),
.B(n_551),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_538),
.B(n_533),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_540),
.B(n_528),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_545),
.B(n_473),
.Y(n_553)
);

AO21x1_ASAP7_75t_L g558 ( 
.A1(n_553),
.A2(n_536),
.B(n_521),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_555),
.B(n_556),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_552),
.B(n_539),
.C(n_544),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_550),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_557),
.A2(n_558),
.B1(n_554),
.B2(n_542),
.Y(n_561)
);

OAI32xp33_ASAP7_75t_L g565 ( 
.A1(n_561),
.A2(n_562),
.A3(n_563),
.B1(n_558),
.B2(n_529),
.Y(n_565)
);

AOI21x1_ASAP7_75t_L g562 ( 
.A1(n_560),
.A2(n_553),
.B(n_523),
.Y(n_562)
);

AOI21x1_ASAP7_75t_L g563 ( 
.A1(n_559),
.A2(n_506),
.B(n_513),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_565),
.A2(n_566),
.B(n_435),
.Y(n_567)
);

BUFx24_ASAP7_75t_SL g566 ( 
.A(n_564),
.Y(n_566)
);

AO21x1_ASAP7_75t_L g568 ( 
.A1(n_567),
.A2(n_417),
.B(n_441),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_568),
.A2(n_445),
.B(n_447),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_451),
.B(n_490),
.Y(n_570)
);


endmodule