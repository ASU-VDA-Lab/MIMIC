module fake_netlist_1_594_n_681 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_681);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_681;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_30), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_53), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_59), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_66), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_47), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_15), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_37), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_18), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_1), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_58), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_44), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_4), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_68), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_24), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_3), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_33), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_69), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_7), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_17), .Y(n_96) );
HB1xp67_ASAP7_75t_L g97 ( .A(n_74), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_56), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_7), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_35), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_61), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_26), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_6), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_36), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_9), .Y(n_105) );
NOR2xp67_ASAP7_75t_L g106 ( .A(n_6), .B(n_60), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_2), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_21), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_54), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_46), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_67), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_1), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_32), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_16), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_57), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_40), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_50), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_2), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_5), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_49), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_28), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_52), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_78), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_97), .B(n_0), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_112), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_78), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_85), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_119), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_103), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_83), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_119), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_86), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_80), .Y(n_135) );
NOR2xp33_ASAP7_75t_R g136 ( .A(n_81), .B(n_34), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_80), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_79), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_89), .B(n_8), .Y(n_139) );
INVxp67_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
AND3x1_ASAP7_75t_L g141 ( .A(n_96), .B(n_8), .C(n_9), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_82), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_93), .Y(n_143) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_87), .B(n_77), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_87), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_109), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_79), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_88), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_122), .B(n_10), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_88), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_107), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_122), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_104), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_84), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_90), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_85), .B(n_10), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_90), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_96), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_99), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_91), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_91), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_99), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_123), .Y(n_163) );
OAI21x1_ASAP7_75t_L g164 ( .A1(n_123), .A2(n_38), .B(n_75), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_105), .Y(n_165) );
NOR2xp33_ASAP7_75t_R g166 ( .A(n_94), .B(n_31), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_140), .B(n_124), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_156), .B(n_105), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_153), .B(n_124), .Y(n_169) );
NAND2x1p5_ASAP7_75t_L g170 ( .A(n_156), .B(n_121), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_125), .B(n_110), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_156), .B(n_121), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_156), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_130), .Y(n_174) );
INVx4_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_163), .Y(n_176) );
AO22x2_ASAP7_75t_L g177 ( .A1(n_144), .A2(n_120), .B1(n_108), .B2(n_113), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_157), .B(n_120), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_142), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_160), .B(n_108), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_125), .B(n_118), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_127), .Y(n_182) );
AND2x6_ASAP7_75t_L g183 ( .A(n_128), .B(n_118), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_163), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_132), .B(n_92), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_128), .A2(n_116), .B1(n_113), .B2(n_95), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_135), .Y(n_188) );
INVx8_ASAP7_75t_L g189 ( .A(n_143), .Y(n_189) );
BUFx2_ASAP7_75t_L g190 ( .A(n_133), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_163), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_144), .A2(n_116), .B1(n_92), .B2(n_95), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_163), .Y(n_193) );
CKINVDCx8_ASAP7_75t_R g194 ( .A(n_134), .Y(n_194) );
AO22x2_ASAP7_75t_L g195 ( .A1(n_135), .A2(n_102), .B1(n_115), .B2(n_114), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_163), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_154), .B(n_117), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_138), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_137), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_165), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_138), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_137), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_145), .B(n_117), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_161), .B(n_115), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_145), .Y(n_205) );
NAND2x1p5_ASAP7_75t_L g206 ( .A(n_126), .B(n_114), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_146), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_148), .B(n_111), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_148), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_150), .B(n_111), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_150), .B(n_110), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_138), .Y(n_212) );
NOR2xp33_ASAP7_75t_SL g213 ( .A(n_131), .B(n_102), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_155), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_155), .B(n_101), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_147), .A2(n_101), .B(n_100), .C(n_98), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_158), .B(n_100), .Y(n_217) );
INVxp33_ASAP7_75t_L g218 ( .A(n_139), .Y(n_218) );
NAND3xp33_ASAP7_75t_L g219 ( .A(n_149), .B(n_98), .C(n_94), .Y(n_219) );
AND2x6_ASAP7_75t_L g220 ( .A(n_147), .B(n_106), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_129), .B(n_11), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_147), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_152), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_152), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_221), .Y(n_225) );
NAND3xp33_ASAP7_75t_SL g226 ( .A(n_174), .B(n_159), .C(n_151), .Y(n_226) );
OR2x6_ASAP7_75t_L g227 ( .A(n_175), .B(n_131), .Y(n_227) );
INVx4_ASAP7_75t_L g228 ( .A(n_170), .Y(n_228) );
INVx3_ASAP7_75t_SL g229 ( .A(n_189), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_173), .A2(n_152), .B(n_164), .C(n_129), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_221), .Y(n_231) );
INVx4_ASAP7_75t_L g232 ( .A(n_170), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_176), .Y(n_233) );
NAND3xp33_ASAP7_75t_SL g234 ( .A(n_174), .B(n_162), .C(n_166), .Y(n_234) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_200), .Y(n_235) );
BUFx2_ASAP7_75t_L g236 ( .A(n_207), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_200), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_183), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_189), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_176), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_221), .Y(n_241) );
NOR3xp33_ASAP7_75t_SL g242 ( .A(n_192), .B(n_141), .C(n_162), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_208), .B(n_164), .Y(n_243) );
BUFx5_ASAP7_75t_L g244 ( .A(n_183), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_208), .B(n_129), .Y(n_245) );
INVx2_ASAP7_75t_SL g246 ( .A(n_195), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_183), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_195), .B(n_129), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_168), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_168), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_168), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_183), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_172), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_183), .Y(n_254) );
INVxp67_ASAP7_75t_L g255 ( .A(n_190), .Y(n_255) );
NAND2xp33_ASAP7_75t_L g256 ( .A(n_177), .B(n_136), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_172), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_195), .B(n_12), .Y(n_258) );
INVx6_ASAP7_75t_L g259 ( .A(n_172), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_198), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_208), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_218), .B(n_41), .Y(n_262) );
NAND2x1p5_ASAP7_75t_L g263 ( .A(n_179), .B(n_13), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_194), .Y(n_264) );
AND2x6_ASAP7_75t_L g265 ( .A(n_210), .B(n_42), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_210), .Y(n_266) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_179), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_188), .A2(n_39), .B(n_72), .Y(n_268) );
INVx4_ASAP7_75t_L g269 ( .A(n_210), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_211), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_189), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_182), .Y(n_272) );
INVx2_ASAP7_75t_SL g273 ( .A(n_211), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_211), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_215), .Y(n_275) );
INVx2_ASAP7_75t_SL g276 ( .A(n_215), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_215), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_177), .A2(n_175), .B1(n_180), .B2(n_178), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_204), .B(n_14), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_199), .B(n_29), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_184), .Y(n_281) );
INVxp67_ASAP7_75t_SL g282 ( .A(n_202), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_177), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_222), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_186), .B(n_14), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_178), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_228), .B(n_178), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_228), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_229), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_228), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_266), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_243), .A2(n_214), .B(n_209), .Y(n_292) );
INVxp67_ASAP7_75t_L g293 ( .A(n_236), .Y(n_293) );
INVx2_ASAP7_75t_SL g294 ( .A(n_266), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_238), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_238), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_284), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_238), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_246), .A2(n_175), .B1(n_204), .B2(n_180), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_266), .B(n_204), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_269), .B(n_180), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_238), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_260), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_259), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_232), .B(n_217), .Y(n_305) );
BUFx4_ASAP7_75t_SL g306 ( .A(n_264), .Y(n_306) );
OR2x6_ASAP7_75t_L g307 ( .A(n_232), .B(n_206), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_232), .B(n_169), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_247), .B(n_206), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_269), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_269), .B(n_167), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_278), .A2(n_218), .B1(n_194), .B2(n_187), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_235), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_246), .A2(n_197), .B1(n_219), .B2(n_213), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_261), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_237), .B(n_197), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_229), .B(n_205), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_254), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_259), .Y(n_319) );
BUFx4f_ASAP7_75t_L g320 ( .A(n_247), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_270), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_247), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_279), .B(n_171), .Y(n_323) );
BUFx12f_ASAP7_75t_L g324 ( .A(n_239), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_255), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_279), .B(n_203), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_279), .B(n_203), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_272), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_225), .A2(n_216), .B(n_181), .C(n_224), .Y(n_329) );
BUFx12f_ASAP7_75t_L g330 ( .A(n_239), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_243), .A2(n_181), .B(n_216), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_274), .Y(n_332) );
CKINVDCx11_ASAP7_75t_R g333 ( .A(n_264), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_273), .A2(n_220), .B1(n_187), .B2(n_223), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_267), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_275), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_288), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_297), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_295), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_288), .Y(n_340) );
NAND3xp33_ASAP7_75t_L g341 ( .A(n_331), .B(n_256), .C(n_230), .Y(n_341) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_299), .B(n_256), .C(n_230), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_323), .B(n_285), .Y(n_343) );
OAI21x1_ASAP7_75t_L g344 ( .A1(n_292), .A2(n_280), .B(n_268), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_302), .Y(n_345) );
INVx3_ASAP7_75t_SL g346 ( .A(n_289), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_323), .B(n_285), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_297), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_290), .B(n_270), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_293), .B(n_286), .Y(n_350) );
NAND2xp33_ASAP7_75t_R g351 ( .A(n_317), .B(n_271), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_312), .A2(n_227), .B1(n_283), .B2(n_234), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_295), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_315), .Y(n_354) );
AOI22xp33_ASAP7_75t_SL g355 ( .A1(n_323), .A2(n_258), .B1(n_227), .B2(n_263), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_315), .B(n_282), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_325), .B(n_226), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_308), .B(n_276), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_316), .A2(n_227), .B1(n_271), .B2(n_273), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_326), .A2(n_227), .B1(n_258), .B2(n_231), .Y(n_360) );
INVx4_ASAP7_75t_L g361 ( .A(n_295), .Y(n_361) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_324), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_332), .B(n_277), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_332), .Y(n_364) );
NOR2xp33_ASAP7_75t_SL g365 ( .A(n_320), .B(n_254), .Y(n_365) );
AOI21xp33_ASAP7_75t_L g366 ( .A1(n_326), .A2(n_262), .B(n_248), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_309), .A2(n_280), .B(n_263), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_295), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_337), .B(n_290), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_338), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g371 ( .A1(n_337), .A2(n_305), .B1(n_324), .B2(n_330), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_355), .A2(n_305), .B1(n_326), .B2(n_327), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_355), .A2(n_305), .B1(n_327), .B2(n_333), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_352), .A2(n_327), .B1(n_333), .B2(n_287), .Y(n_374) );
NOR2x1_ASAP7_75t_SL g375 ( .A(n_361), .B(n_295), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_337), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_338), .B(n_248), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g378 ( .A1(n_360), .A2(n_242), .B1(n_314), .B2(n_301), .C(n_300), .Y(n_378) );
OAI221xp5_ASAP7_75t_SL g379 ( .A1(n_360), .A2(n_335), .B1(n_317), .B2(n_328), .C(n_313), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_348), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_348), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_354), .Y(n_382) );
OAI221xp5_ASAP7_75t_SL g383 ( .A1(n_359), .A2(n_334), .B1(n_307), .B2(n_336), .C(n_245), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_357), .A2(n_308), .B1(n_265), .B2(n_276), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_354), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_364), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_343), .A2(n_308), .B1(n_265), .B2(n_321), .Y(n_387) );
AO21x2_ASAP7_75t_L g388 ( .A1(n_341), .A2(n_329), .B(n_241), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_368), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_364), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_363), .Y(n_391) );
OAI21xp33_ASAP7_75t_L g392 ( .A1(n_341), .A2(n_336), .B(n_311), .Y(n_392) );
AOI222xp33_ASAP7_75t_L g393 ( .A1(n_343), .A2(n_330), .B1(n_257), .B2(n_253), .C1(n_251), .C2(n_250), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_340), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_342), .B(n_184), .C(n_191), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_347), .A2(n_220), .B1(n_265), .B2(n_321), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_378), .A2(n_347), .B1(n_342), .B2(n_366), .C(n_350), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_370), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_370), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_393), .A2(n_366), .B1(n_358), .B2(n_265), .Y(n_401) );
AOI33xp33_ASAP7_75t_L g402 ( .A1(n_371), .A2(n_358), .A3(n_304), .B1(n_319), .B2(n_340), .B3(n_198), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_373), .A2(n_350), .B(n_290), .C(n_356), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_379), .A2(n_356), .B1(n_346), .B2(n_363), .Y(n_404) );
AO21x1_ASAP7_75t_SL g405 ( .A1(n_376), .A2(n_391), .B(n_372), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_394), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_371), .B(n_346), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_395), .A2(n_353), .B(n_339), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_385), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_385), .B(n_346), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_385), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_380), .Y(n_412) );
BUFx5_ASAP7_75t_L g413 ( .A(n_391), .Y(n_413) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_379), .B(n_351), .C(n_306), .D(n_249), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_394), .Y(n_415) );
OAI211xp5_ASAP7_75t_SL g416 ( .A1(n_393), .A2(n_201), .B(n_212), .C(n_310), .Y(n_416) );
AND2x6_ASAP7_75t_L g417 ( .A(n_389), .B(n_368), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_378), .A2(n_265), .B1(n_220), .B2(n_349), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_380), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_376), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_381), .B(n_367), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_382), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_382), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_386), .B(n_349), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_369), .Y(n_426) );
OAI22xp5_ASAP7_75t_SL g427 ( .A1(n_374), .A2(n_362), .B1(n_307), .B2(n_349), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_369), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_383), .A2(n_259), .B1(n_361), .B2(n_349), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_386), .Y(n_430) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_402), .B(n_383), .C(n_384), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_399), .B(n_390), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_399), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_422), .B(n_388), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_412), .B(n_390), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_412), .Y(n_436) );
INVxp67_ASAP7_75t_L g437 ( .A(n_406), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_422), .B(n_388), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_419), .B(n_377), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_397), .Y(n_440) );
INVx4_ASAP7_75t_L g441 ( .A(n_413), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_401), .A2(n_387), .B1(n_396), .B2(n_369), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_408), .A2(n_395), .B(n_392), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_400), .B(n_388), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_417), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_419), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_400), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_397), .B(n_409), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_413), .Y(n_449) );
OAI21xp5_ASAP7_75t_L g450 ( .A1(n_404), .A2(n_392), .B(n_367), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_409), .B(n_388), .Y(n_451) );
NAND5xp2_ASAP7_75t_SL g452 ( .A(n_403), .B(n_396), .C(n_362), .D(n_17), .E(n_18), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_424), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_411), .B(n_389), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_413), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_414), .B(n_307), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_411), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_421), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_424), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_430), .B(n_389), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_430), .B(n_389), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_421), .Y(n_462) );
BUFx8_ASAP7_75t_L g463 ( .A(n_413), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_423), .Y(n_464) );
AOI33xp33_ASAP7_75t_L g465 ( .A1(n_418), .A2(n_377), .A3(n_212), .B1(n_201), .B2(n_369), .B3(n_196), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_423), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_413), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_413), .B(n_389), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_413), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_413), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_405), .B(n_389), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_417), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_415), .Y(n_473) );
INVx3_ASAP7_75t_L g474 ( .A(n_417), .Y(n_474) );
INVx4_ASAP7_75t_L g475 ( .A(n_417), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_425), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_417), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_405), .B(n_426), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_463), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_448), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_436), .Y(n_481) );
NOR2xp33_ASAP7_75t_SL g482 ( .A(n_463), .B(n_414), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_473), .Y(n_483) );
INVx3_ASAP7_75t_SL g484 ( .A(n_441), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_436), .Y(n_485) );
NOR4xp25_ASAP7_75t_SL g486 ( .A(n_449), .B(n_407), .C(n_398), .D(n_427), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_433), .B(n_410), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_434), .B(n_428), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_433), .B(n_410), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_434), .B(n_420), .Y(n_490) );
AND2x2_ASAP7_75t_SL g491 ( .A(n_441), .B(n_449), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_448), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_463), .Y(n_493) );
AND2x4_ASAP7_75t_L g494 ( .A(n_474), .B(n_417), .Y(n_494) );
NOR2x1_ASAP7_75t_L g495 ( .A(n_441), .B(n_429), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_456), .B(n_427), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_434), .B(n_389), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_437), .B(n_15), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_447), .B(n_429), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_476), .B(n_377), .Y(n_500) );
BUFx2_ASAP7_75t_L g501 ( .A(n_463), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_476), .B(n_220), .Y(n_502) );
AND3x2_ASAP7_75t_L g503 ( .A(n_455), .B(n_365), .C(n_19), .Y(n_503) );
OAI21xp5_ASAP7_75t_SL g504 ( .A1(n_431), .A2(n_416), .B(n_345), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_439), .B(n_220), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_465), .A2(n_367), .B(n_345), .C(n_365), .Y(n_506) );
NOR4xp25_ASAP7_75t_SL g507 ( .A(n_455), .B(n_375), .C(n_19), .D(n_20), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_473), .Y(n_508) );
AND4x1_ASAP7_75t_L g509 ( .A(n_431), .B(n_16), .C(n_20), .D(n_21), .Y(n_509) );
NOR2x1_ASAP7_75t_L g510 ( .A(n_441), .B(n_361), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_458), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_438), .B(n_375), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_437), .B(n_22), .Y(n_513) );
NAND2x1_ASAP7_75t_SL g514 ( .A(n_474), .B(n_361), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_458), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_439), .B(n_417), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_446), .B(n_22), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_448), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_452), .A2(n_265), .B1(n_345), .B2(n_344), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_467), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_447), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_446), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_467), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_453), .B(n_345), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_435), .B(n_307), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_453), .B(n_353), .Y(n_526) );
NOR2xp33_ASAP7_75t_R g527 ( .A(n_463), .B(n_368), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_459), .B(n_339), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_460), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_459), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_460), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_438), .B(n_344), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_435), .B(n_339), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_432), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_432), .Y(n_535) );
AOI322xp5_ASAP7_75t_L g536 ( .A1(n_496), .A2(n_438), .A3(n_478), .B1(n_462), .B2(n_464), .C1(n_466), .C2(n_452), .Y(n_536) );
AOI21xp33_ASAP7_75t_L g537 ( .A1(n_498), .A2(n_432), .B(n_444), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_479), .A2(n_469), .B1(n_470), .B2(n_442), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g539 ( .A1(n_513), .A2(n_442), .B1(n_450), .B2(n_462), .C(n_464), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_506), .A2(n_450), .B(n_470), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_534), .B(n_451), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_482), .A2(n_478), .B1(n_469), .B2(n_451), .Y(n_542) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_479), .B(n_501), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_535), .B(n_451), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_525), .A2(n_478), .B1(n_471), .B2(n_474), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_483), .B(n_466), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_487), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_508), .B(n_474), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_487), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_501), .A2(n_471), .B1(n_445), .B2(n_475), .Y(n_550) );
NOR2x1_ASAP7_75t_L g551 ( .A(n_510), .B(n_475), .Y(n_551) );
OAI211xp5_ASAP7_75t_L g552 ( .A1(n_486), .A2(n_527), .B(n_504), .C(n_493), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_480), .B(n_458), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_481), .Y(n_554) );
AOI211xp5_ASAP7_75t_SL g555 ( .A1(n_506), .A2(n_471), .B(n_468), .C(n_477), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_492), .B(n_440), .Y(n_556) );
INVx2_ASAP7_75t_SL g557 ( .A(n_493), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_485), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_522), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_491), .A2(n_475), .B1(n_445), .B2(n_440), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_509), .B(n_475), .Y(n_561) );
OAI22xp33_ASAP7_75t_L g562 ( .A1(n_484), .A2(n_445), .B1(n_472), .B2(n_477), .Y(n_562) );
OAI211xp5_ASAP7_75t_L g563 ( .A1(n_527), .A2(n_477), .B(n_472), .C(n_444), .Y(n_563) );
OAI21xp33_ASAP7_75t_L g564 ( .A1(n_491), .A2(n_512), .B(n_490), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g565 ( .A1(n_512), .A2(n_461), .B(n_460), .Y(n_565) );
OAI21xp33_ASAP7_75t_SL g566 ( .A1(n_495), .A2(n_468), .B(n_472), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_530), .Y(n_567) );
OAI32xp33_ASAP7_75t_L g568 ( .A1(n_489), .A2(n_457), .A3(n_440), .B1(n_468), .B2(n_461), .Y(n_568) );
OAI22x1_ASAP7_75t_L g569 ( .A1(n_484), .A2(n_457), .B1(n_461), .B2(n_454), .Y(n_569) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_517), .A2(n_443), .B1(n_457), .B2(n_454), .C(n_185), .Y(n_570) );
NAND2xp33_ASAP7_75t_L g571 ( .A(n_489), .B(n_521), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_490), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_520), .A2(n_443), .B(n_454), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_488), .B(n_23), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_518), .B(n_344), .Y(n_575) );
OAI22xp33_ASAP7_75t_L g576 ( .A1(n_499), .A2(n_353), .B1(n_320), .B2(n_291), .Y(n_576) );
OAI32xp33_ASAP7_75t_L g577 ( .A1(n_523), .A2(n_196), .A3(n_193), .B1(n_185), .B2(n_302), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_488), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_529), .B(n_193), .Y(n_579) );
AOI31xp33_ASAP7_75t_L g580 ( .A1(n_499), .A2(n_291), .A3(n_294), .B(n_303), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_500), .B(n_25), .Y(n_581) );
AOI22xp33_ASAP7_75t_SL g582 ( .A1(n_494), .A2(n_516), .B1(n_531), .B2(n_532), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_532), .A2(n_303), .B1(n_310), .B2(n_294), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_497), .B(n_191), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_505), .A2(n_310), .B1(n_259), .B2(n_184), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_497), .B(n_184), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_503), .A2(n_191), .B1(n_318), .B2(n_260), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_537), .B(n_524), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_556), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_554), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_558), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_557), .Y(n_592) );
CKINVDCx16_ASAP7_75t_R g593 ( .A(n_574), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_539), .A2(n_502), .B1(n_519), .B2(n_533), .C(n_494), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_572), .B(n_494), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_547), .B(n_515), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_559), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_561), .Y(n_598) );
NOR3xp33_ASAP7_75t_SL g599 ( .A(n_552), .B(n_528), .C(n_526), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_543), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_567), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_549), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_578), .B(n_515), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_546), .B(n_511), .Y(n_604) );
NOR3xp33_ASAP7_75t_SL g605 ( .A(n_564), .B(n_507), .C(n_514), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_582), .B(n_511), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_571), .B(n_514), .Y(n_607) );
NOR3xp33_ASAP7_75t_SL g608 ( .A(n_566), .B(n_27), .C(n_43), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_541), .B(n_191), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_544), .B(n_45), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_548), .B(n_48), .Y(n_611) );
XNOR2xp5_ASAP7_75t_L g612 ( .A(n_543), .B(n_51), .Y(n_612) );
NAND2xp33_ASAP7_75t_R g613 ( .A(n_573), .B(n_55), .Y(n_613) );
NOR3xp33_ASAP7_75t_SL g614 ( .A(n_538), .B(n_62), .C(n_63), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_569), .B(n_320), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_551), .B(n_322), .Y(n_616) );
AOI211xp5_ASAP7_75t_L g617 ( .A1(n_560), .A2(n_247), .B(n_252), .C(n_322), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_553), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_575), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_580), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_584), .Y(n_621) );
XOR2x2_ASAP7_75t_L g622 ( .A(n_560), .B(n_64), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_536), .B(n_65), .Y(n_623) );
NAND2xp33_ASAP7_75t_R g624 ( .A(n_540), .B(n_70), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_590), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_591), .Y(n_626) );
AOI21xp33_ASAP7_75t_L g627 ( .A1(n_620), .A2(n_580), .B(n_581), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_588), .B(n_565), .Y(n_628) );
AOI21xp33_ASAP7_75t_SL g629 ( .A1(n_593), .A2(n_562), .B(n_550), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_597), .Y(n_630) );
AO22x2_ASAP7_75t_L g631 ( .A1(n_601), .A2(n_563), .B1(n_555), .B2(n_568), .Y(n_631) );
XNOR2x1_ASAP7_75t_L g632 ( .A(n_622), .B(n_545), .Y(n_632) );
OAI211xp5_ASAP7_75t_SL g633 ( .A1(n_599), .A2(n_555), .B(n_587), .C(n_570), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_600), .B(n_542), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_602), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_622), .A2(n_576), .B(n_577), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_588), .B(n_586), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_604), .Y(n_638) );
OAI32xp33_ASAP7_75t_L g639 ( .A1(n_613), .A2(n_579), .A3(n_583), .B1(n_585), .B2(n_318), .Y(n_639) );
INVxp67_ASAP7_75t_SL g640 ( .A(n_613), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_606), .A2(n_260), .B1(n_318), .B2(n_322), .C(n_298), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_618), .B(n_71), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_603), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_592), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_621), .B(n_76), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_600), .B(n_322), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_598), .B(n_322), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_638), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_643), .B(n_619), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_632), .A2(n_594), .B1(n_623), .B2(n_607), .Y(n_650) );
INVx6_ASAP7_75t_L g651 ( .A(n_644), .Y(n_651) );
AOI322xp5_ASAP7_75t_L g652 ( .A1(n_640), .A2(n_607), .A3(n_595), .B1(n_615), .B2(n_589), .C1(n_605), .C2(n_608), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_625), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_628), .B(n_619), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g655 ( .A1(n_640), .A2(n_615), .B1(n_589), .B2(n_621), .C1(n_612), .C2(n_610), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_629), .B(n_596), .Y(n_656) );
XNOR2xp5_ASAP7_75t_L g657 ( .A(n_637), .B(n_614), .Y(n_657) );
AND2x4_ASAP7_75t_L g658 ( .A(n_634), .B(n_616), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_631), .A2(n_611), .B1(n_616), .B2(n_609), .C(n_617), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_626), .Y(n_660) );
NAND4xp75_ASAP7_75t_L g661 ( .A(n_636), .B(n_624), .C(n_298), .D(n_296), .Y(n_661) );
OAI222xp33_ASAP7_75t_L g662 ( .A1(n_630), .A2(n_624), .B1(n_240), .B2(n_233), .C1(n_296), .C2(n_298), .Y(n_662) );
OAI321xp33_ASAP7_75t_L g663 ( .A1(n_633), .A2(n_296), .A3(n_298), .B1(n_252), .B2(n_281), .C(n_233), .Y(n_663) );
OAI322xp33_ASAP7_75t_L g664 ( .A1(n_635), .A2(n_296), .A3(n_298), .B1(n_252), .B2(n_240), .C1(n_281), .C2(n_244), .Y(n_664) );
OAI211xp5_ASAP7_75t_SL g665 ( .A1(n_627), .A2(n_244), .B(n_252), .C(n_296), .Y(n_665) );
AOI211xp5_ASAP7_75t_SL g666 ( .A1(n_633), .A2(n_244), .B(n_281), .C(n_647), .Y(n_666) );
NAND4xp25_ASAP7_75t_L g667 ( .A(n_639), .B(n_244), .C(n_281), .D(n_641), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_631), .Y(n_668) );
A2O1A1Ixp33_ASAP7_75t_L g669 ( .A1(n_646), .A2(n_244), .B(n_642), .C(n_631), .Y(n_669) );
AND2x4_ASAP7_75t_L g670 ( .A(n_658), .B(n_648), .Y(n_670) );
NOR4xp25_ASAP7_75t_L g671 ( .A(n_668), .B(n_650), .C(n_669), .D(n_656), .Y(n_671) );
INVx1_ASAP7_75t_SL g672 ( .A(n_651), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_657), .A2(n_667), .B(n_659), .C(n_663), .Y(n_673) );
OAI322xp33_ASAP7_75t_L g674 ( .A1(n_672), .A2(n_654), .A3(n_660), .B1(n_653), .B2(n_649), .C1(n_655), .C2(n_651), .Y(n_674) );
NOR4xp25_ASAP7_75t_L g675 ( .A(n_671), .B(n_662), .C(n_665), .D(n_645), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_670), .B(n_658), .Y(n_676) );
INVx8_ASAP7_75t_L g677 ( .A(n_676), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_674), .A2(n_673), .B(n_670), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_677), .A2(n_675), .B1(n_661), .B2(n_652), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_679), .A2(n_678), .B1(n_666), .B2(n_664), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_680), .A2(n_244), .B(n_678), .Y(n_681) );
endmodule