module fake_jpeg_29812_n_325 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_12),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_12),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_12),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_25),
.Y(n_82)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_56),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_59),
.B(n_60),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_19),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_82),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_63),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_80),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_28),
.B1(n_15),
.B2(n_29),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_73),
.A2(n_79),
.B1(n_84),
.B2(n_13),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_35),
.B1(n_33),
.B2(n_29),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_23),
.C(n_26),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_40),
.A2(n_45),
.B1(n_44),
.B2(n_39),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_21),
.B1(n_31),
.B2(n_17),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_87),
.A2(n_88),
.B1(n_92),
.B2(n_126),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_21),
.B1(n_31),
.B2(n_17),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_89),
.B(n_95),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_91),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_21),
.B1(n_31),
.B2(n_17),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_62),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_97),
.B(n_103),
.Y(n_152)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_34),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_105),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_68),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_104),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_34),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_34),
.B(n_22),
.C(n_26),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_13),
.B(n_77),
.C(n_20),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_67),
.A2(n_26),
.B1(n_22),
.B2(n_33),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_25),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_110),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_109),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_68),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_114),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_22),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_31),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_67),
.A2(n_13),
.B1(n_31),
.B2(n_21),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_13),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_84),
.A2(n_13),
.B1(n_31),
.B2(n_21),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_68),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_0),
.Y(n_129)
);

BUFx8_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_81),
.A2(n_21),
.B1(n_13),
.B2(n_20),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_129),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_102),
.C(n_121),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_131),
.B(n_6),
.C(n_7),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_118),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_95),
.B(n_0),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_139),
.B(n_141),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_99),
.A2(n_101),
.B1(n_127),
.B2(n_116),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g194 ( 
.A(n_143),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_86),
.A2(n_113),
.B1(n_77),
.B2(n_105),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_123),
.B1(n_112),
.B2(n_98),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_86),
.A2(n_66),
.B1(n_61),
.B2(n_32),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_155),
.B(n_158),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_66),
.B1(n_61),
.B2(n_32),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_160),
.B1(n_101),
.B2(n_97),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_103),
.A2(n_32),
.B(n_20),
.C(n_2),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_99),
.A2(n_0),
.B(n_1),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_106),
.A2(n_32),
.B1(n_20),
.B2(n_3),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_165),
.A2(n_175),
.B1(n_149),
.B2(n_133),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_166),
.B(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_171),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_144),
.B1(n_140),
.B2(n_131),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_170),
.B1(n_183),
.B2(n_190),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_128),
.B1(n_111),
.B2(n_100),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_91),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_96),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_180),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_139),
.B(n_93),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_177),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_117),
.B1(n_115),
.B2(n_104),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_118),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_146),
.B(n_89),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_125),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_125),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_189),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_147),
.A2(n_109),
.B1(n_90),
.B2(n_32),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_20),
.Y(n_184)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_136),
.Y(n_186)
);

AOI22x1_ASAP7_75t_L g187 ( 
.A1(n_141),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_151),
.B(n_148),
.Y(n_221)
);

NOR2x1_ASAP7_75t_L g188 ( 
.A(n_129),
.B(n_3),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_8),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_4),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_138),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_152),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_9),
.B1(n_11),
.B2(n_148),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_6),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_195),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_151),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_7),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_163),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_205),
.B1(n_170),
.B2(n_194),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_158),
.B(n_155),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_188),
.B(n_182),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_194),
.A2(n_133),
.B1(n_150),
.B2(n_132),
.Y(n_205)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_157),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_215),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_149),
.B(n_157),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_211),
.A2(n_212),
.B(n_224),
.Y(n_241)
);

AND2x6_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_149),
.Y(n_212)
);

AO22x1_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_132),
.B1(n_162),
.B2(n_130),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_164),
.B(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_189),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_130),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_218),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_145),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_219),
.B(n_190),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_183),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_165),
.B1(n_194),
.B2(n_175),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_176),
.A2(n_136),
.B(n_137),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_204),
.B1(n_214),
.B2(n_199),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_180),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_242),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_218),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_233),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_245),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_211),
.A2(n_187),
.B(n_181),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_237),
.B(n_244),
.Y(n_259)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_239),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_240),
.A2(n_246),
.B1(n_214),
.B2(n_199),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_193),
.C(n_196),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_197),
.A2(n_187),
.B1(n_179),
.B2(n_191),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_186),
.B(n_145),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_248),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_200),
.A2(n_153),
.B(n_137),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_210),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_228),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_257),
.A2(n_265),
.B1(n_267),
.B2(n_233),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_215),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_264),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_234),
.A2(n_204),
.B1(n_200),
.B2(n_216),
.Y(n_263)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_263),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_219),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_248),
.B(n_213),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_203),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_225),
.A2(n_212),
.B1(n_202),
.B2(n_217),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_268),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_247),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_269),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_270),
.A2(n_259),
.B1(n_267),
.B2(n_265),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_249),
.A2(n_246),
.B1(n_235),
.B2(n_240),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_283),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_241),
.C(n_227),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_277),
.Y(n_284)
);

OAI31xp33_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_241),
.A3(n_236),
.B(n_237),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_275),
.A2(n_282),
.B(n_251),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_281),
.Y(n_286)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_203),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_279),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_250),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_253),
.B(n_206),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_280),
.A2(n_258),
.B1(n_244),
.B2(n_239),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_228),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_206),
.B(n_227),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_260),
.A2(n_231),
.B1(n_236),
.B2(n_209),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_290),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_274),
.A2(n_252),
.B1(n_256),
.B2(n_255),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_287),
.A2(n_288),
.B1(n_220),
.B2(n_222),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_269),
.A2(n_275),
.B1(n_270),
.B2(n_251),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_292),
.B(n_276),
.Y(n_298)
);

AOI21xp33_ASAP7_75t_L g292 ( 
.A1(n_273),
.A2(n_243),
.B(n_238),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_269),
.A2(n_229),
.B1(n_221),
.B2(n_232),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_229),
.B1(n_221),
.B2(n_281),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_272),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_302),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_299),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_221),
.B(n_207),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_303),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_272),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_153),
.Y(n_304)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_304),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_11),
.B1(n_220),
.B2(n_296),
.Y(n_305)
);

NOR2x1_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_287),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_311),
.Y(n_313)
);

AOI21xp33_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_284),
.B(n_294),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_297),
.B(n_291),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_302),
.C(n_289),
.Y(n_314)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_314),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_288),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_315),
.B(n_316),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_294),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_299),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_306),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_293),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_310),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_319),
.C(n_313),
.Y(n_323)
);

AOI321xp33_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_313),
.A3(n_318),
.B1(n_320),
.B2(n_309),
.C(n_305),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_301),
.Y(n_325)
);


endmodule