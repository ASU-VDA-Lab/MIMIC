module fake_netlist_6_4827_n_1693 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1693);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1693;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_16),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_112),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_109),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_1),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_40),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_58),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_114),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_121),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_88),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_31),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_65),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_21),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_35),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_116),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_4),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_17),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_30),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_69),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_115),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_47),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_24),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_124),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_17),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_126),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_22),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_76),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_81),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_63),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_125),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_24),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_73),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_64),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_4),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_83),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_90),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_66),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_26),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_67),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_46),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_26),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_47),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_3),
.Y(n_207)
);

BUFx8_ASAP7_75t_SL g208 ( 
.A(n_51),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_100),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_136),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_70),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_147),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_144),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_12),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_133),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_30),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_27),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_34),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_127),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_57),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_16),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_55),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_72),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_71),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_45),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_9),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_40),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_7),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_28),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_11),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_10),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_19),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_99),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_41),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_148),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_151),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_89),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_53),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_51),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_108),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_60),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_94),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_6),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_130),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_104),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_68),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_84),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_102),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_119),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_111),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_138),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_10),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_12),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_92),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_59),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_43),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_43),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_139),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_62),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_145),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_3),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_78),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_152),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_101),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_132),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_113),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_28),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_1),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_39),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_87),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_41),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_56),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_36),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_106),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_153),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_46),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_5),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_13),
.Y(n_279)
);

BUFx2_ASAP7_75t_SL g280 ( 
.A(n_44),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_38),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_20),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_22),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_128),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_18),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_48),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_155),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_39),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_48),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_54),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_7),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_82),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_5),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_21),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_154),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_91),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_129),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_98),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_74),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_140),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_52),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_14),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_117),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_105),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_75),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_107),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_80),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_86),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_20),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_31),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_208),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_158),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_228),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_201),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_228),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_228),
.Y(n_317)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_201),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_159),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_184),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_199),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_160),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_182),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_228),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_228),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_285),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_0),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_182),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_163),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_165),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_2),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_197),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_225),
.B(n_2),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_269),
.B(n_6),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_166),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_157),
.Y(n_338)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_162),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_168),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_183),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_188),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_278),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_171),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_278),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_167),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_278),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_278),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_161),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_176),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_177),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_180),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_190),
.B(n_8),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_181),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_190),
.B(n_8),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_276),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_186),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_187),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_189),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_269),
.B(n_9),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_200),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_183),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_191),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_203),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_210),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_211),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_212),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_169),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_213),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_219),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_161),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_234),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_236),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_254),
.B(n_11),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_254),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_257),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_239),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_170),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_175),
.B(n_310),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_257),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_195),
.B(n_13),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_242),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_248),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_250),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_320),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_312),
.Y(n_387)
);

AND3x2_ASAP7_75t_L g388 ( 
.A(n_353),
.B(n_277),
.C(n_243),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_321),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_313),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_319),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_322),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_316),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_317),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_379),
.B(n_306),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_340),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_342),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_356),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_324),
.B(n_325),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_330),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_325),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_332),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_337),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_331),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_331),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_314),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_343),
.B(n_255),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_350),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_379),
.B(n_175),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_345),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_347),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_347),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_356),
.B(n_274),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_351),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_352),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_348),
.B(n_238),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_348),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_314),
.B(n_263),
.Y(n_424)
);

XOR2x2_ASAP7_75t_L g425 ( 
.A(n_318),
.B(n_216),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_342),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_349),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_344),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_371),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_359),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_375),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_354),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_376),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_357),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_358),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_314),
.B(n_310),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_336),
.B(n_276),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_376),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_365),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_380),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_366),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_361),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_327),
.B(n_188),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_380),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_364),
.Y(n_447)
);

AND2x6_ASAP7_75t_L g448 ( 
.A(n_327),
.B(n_188),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_333),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_333),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g451 ( 
.A(n_355),
.B(n_205),
.C(n_191),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_449),
.B(n_369),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_414),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_411),
.Y(n_457)
);

INVx6_ASAP7_75t_L g458 ( 
.A(n_411),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_450),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_411),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_449),
.B(n_238),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_338),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_396),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_195),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_426),
.B(n_243),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_397),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_387),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_399),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_438),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_424),
.B(n_346),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_424),
.B(n_339),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_398),
.B(n_196),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_426),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_412),
.B(n_368),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_426),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_385),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_398),
.B(n_196),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_414),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_419),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_439),
.A2(n_335),
.B1(n_384),
.B2(n_315),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_398),
.B(n_198),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_390),
.Y(n_484)
);

AND2x6_ASAP7_75t_L g485 ( 
.A(n_438),
.B(n_198),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_397),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_412),
.B(n_370),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_426),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_390),
.Y(n_489)
);

OR2x6_ASAP7_75t_L g490 ( 
.A(n_452),
.B(n_326),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_390),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_438),
.B(n_378),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_395),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_439),
.A2(n_315),
.B1(n_334),
.B2(n_360),
.Y(n_494)
);

BUFx10_ASAP7_75t_L g495 ( 
.A(n_393),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_414),
.B(n_372),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_395),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_444),
.B(n_373),
.Y(n_498)
);

INVxp33_ASAP7_75t_SL g499 ( 
.A(n_419),
.Y(n_499)
);

INVx5_ASAP7_75t_L g500 ( 
.A(n_445),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_391),
.B(n_377),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_392),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_451),
.A2(n_381),
.B1(n_341),
.B2(n_362),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_395),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_394),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_426),
.B(n_246),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_416),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_452),
.B(n_382),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_452),
.B(n_383),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_408),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_391),
.B(n_164),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_444),
.B(n_326),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_391),
.B(n_400),
.Y(n_514)
);

AND2x6_ASAP7_75t_L g515 ( 
.A(n_426),
.B(n_215),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_416),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_444),
.B(n_328),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_392),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_408),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_444),
.B(n_341),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_392),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_409),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_409),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_416),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_404),
.B(n_406),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_391),
.B(n_400),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_410),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_386),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_410),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_392),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_400),
.B(n_402),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_400),
.B(n_192),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_445),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_425),
.B(n_360),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_451),
.B(n_362),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_402),
.B(n_193),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_402),
.B(n_246),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_407),
.B(n_363),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_415),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_402),
.B(n_245),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_392),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_413),
.B(n_420),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_415),
.Y(n_543)
);

NOR2x1_ASAP7_75t_L g544 ( 
.A(n_403),
.B(n_336),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_389),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_421),
.B(n_284),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_422),
.B(n_215),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_423),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_445),
.B(n_448),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_433),
.B(n_284),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_418),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_436),
.B(n_363),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_423),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_417),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_417),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_418),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_437),
.B(n_222),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_422),
.B(n_220),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_445),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_429),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_417),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_447),
.B(n_188),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_422),
.B(n_220),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_448),
.A2(n_291),
.B1(n_205),
.B2(n_206),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_423),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_422),
.B(n_188),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_445),
.A2(n_206),
.B1(n_233),
.B2(n_240),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_403),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_425),
.B(n_311),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_430),
.B(n_280),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_445),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_388),
.B(n_374),
.Y(n_572)
);

AND2x6_ASAP7_75t_L g573 ( 
.A(n_430),
.B(n_223),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_388),
.B(n_172),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_427),
.B(n_173),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_423),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_423),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_435),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_445),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_423),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_435),
.B(n_209),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_445),
.A2(n_233),
.B1(n_302),
.B2(n_291),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_401),
.B(n_323),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_435),
.Y(n_584)
);

NAND3x1_ASAP7_75t_L g585 ( 
.A(n_425),
.B(n_289),
.C(n_283),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_435),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_448),
.A2(n_262),
.B1(n_240),
.B2(n_253),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_427),
.B(n_174),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_435),
.Y(n_589)
);

BUFx4f_ASAP7_75t_L g590 ( 
.A(n_448),
.Y(n_590)
);

AND3x2_ASAP7_75t_L g591 ( 
.A(n_432),
.B(n_262),
.C(n_253),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_432),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_448),
.Y(n_593)
);

AND2x6_ASAP7_75t_L g594 ( 
.A(n_434),
.B(n_223),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_448),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_434),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_448),
.A2(n_329),
.B1(n_268),
.B2(n_229),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_448),
.B(n_264),
.Y(n_598)
);

INVx5_ASAP7_75t_L g599 ( 
.A(n_435),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_568),
.B(n_427),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_471),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_477),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_454),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_476),
.A2(n_401),
.B1(n_275),
.B2(n_265),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_469),
.B(n_431),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_454),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_477),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_590),
.B(n_209),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_538),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_453),
.B(n_178),
.Y(n_610)
);

AOI221xp5_ASAP7_75t_L g611 ( 
.A1(n_535),
.A2(n_226),
.B1(n_270),
.B2(n_221),
.C(n_294),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_457),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_492),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_487),
.B(n_427),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_590),
.B(n_209),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_487),
.B(n_224),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_455),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_463),
.B(n_179),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_463),
.B(n_185),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_500),
.B(n_533),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_520),
.B(n_472),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_457),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_471),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_456),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_476),
.A2(n_287),
.B1(n_266),
.B2(n_271),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_538),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_459),
.B(n_224),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_500),
.B(n_533),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_520),
.B(n_237),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_473),
.B(n_194),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_L g631 ( 
.A1(n_534),
.A2(n_374),
.B1(n_281),
.B2(n_283),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_549),
.A2(n_237),
.B(n_241),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_552),
.B(n_480),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_473),
.B(n_241),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_575),
.B(n_247),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_575),
.B(n_588),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_588),
.B(n_247),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_R g638 ( 
.A(n_495),
.B(n_441),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_478),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_552),
.B(n_443),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_535),
.B(n_202),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_592),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_544),
.B(n_249),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_512),
.B(n_249),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_517),
.B(n_204),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_502),
.A2(n_297),
.B1(n_251),
.B2(n_308),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_596),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_532),
.A2(n_297),
.B1(n_251),
.B2(n_308),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_513),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_478),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_494),
.B(n_280),
.Y(n_651)
);

O2A1O1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_462),
.A2(n_281),
.B(n_289),
.C(n_302),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_496),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_464),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_536),
.B(n_252),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_540),
.B(n_252),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_477),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_513),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_517),
.B(n_207),
.Y(n_659)
);

A2O1A1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_504),
.A2(n_290),
.B(n_259),
.C(n_260),
.Y(n_660)
);

NAND2x1p5_ASAP7_75t_L g661 ( 
.A(n_593),
.B(n_256),
.Y(n_661)
);

BUFx12f_ASAP7_75t_L g662 ( 
.A(n_495),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_467),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_465),
.B(n_256),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_509),
.B(n_274),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_458),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_470),
.Y(n_667)
);

INVxp33_ASAP7_75t_L g668 ( 
.A(n_583),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_465),
.B(n_259),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_510),
.B(n_274),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_465),
.B(n_260),
.Y(n_671)
);

INVxp33_ASAP7_75t_L g672 ( 
.A(n_542),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_465),
.B(n_261),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_465),
.B(n_261),
.Y(n_674)
);

OAI221xp5_ASAP7_75t_L g675 ( 
.A1(n_504),
.A2(n_307),
.B1(n_290),
.B2(n_267),
.C(n_446),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_484),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_468),
.B(n_267),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_484),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_486),
.B(n_307),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_546),
.B(n_214),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_597),
.A2(n_296),
.B1(n_273),
.B2(n_292),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_533),
.B(n_295),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_501),
.B(n_428),
.Y(n_683)
);

A2O1A1Ixp33_ASAP7_75t_L g684 ( 
.A1(n_564),
.A2(n_446),
.B(n_442),
.C(n_440),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_474),
.A2(n_305),
.B1(n_298),
.B2(n_303),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_511),
.B(n_442),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_461),
.B(n_440),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_519),
.B(n_428),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_525),
.B(n_309),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_522),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_528),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_474),
.A2(n_304),
.B1(n_300),
.B2(n_276),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_523),
.B(n_301),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_527),
.B(n_293),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_529),
.B(n_288),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_539),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_543),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_489),
.Y(n_698)
);

NOR3xp33_ASAP7_75t_L g699 ( 
.A(n_482),
.B(n_286),
.C(n_282),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_557),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_551),
.B(n_279),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_572),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_489),
.Y(n_703)
);

NOR2x1p5_ASAP7_75t_L g704 ( 
.A(n_569),
.B(n_272),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_475),
.A2(n_526),
.B(n_531),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_556),
.B(n_258),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_458),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_546),
.B(n_550),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_491),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_559),
.B(n_244),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_564),
.A2(n_235),
.B1(n_232),
.B2(n_231),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_490),
.B(n_230),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_477),
.B(n_227),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_572),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_550),
.B(n_557),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_559),
.B(n_218),
.Y(n_716)
);

O2A1O1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_462),
.A2(n_217),
.B(n_15),
.C(n_18),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_498),
.B(n_156),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_498),
.B(n_150),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_545),
.B(n_14),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_481),
.B(n_19),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_491),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_458),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_490),
.B(n_23),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_474),
.B(n_142),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_493),
.Y(n_726)
);

NOR2xp67_ASAP7_75t_L g727 ( 
.A(n_542),
.B(n_135),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_493),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_497),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_497),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_574),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_505),
.Y(n_732)
);

CKINVDCx8_ASAP7_75t_R g733 ( 
.A(n_560),
.Y(n_733)
);

INVx8_ASAP7_75t_L g734 ( 
.A(n_490),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_506),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_562),
.B(n_23),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_505),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_508),
.Y(n_738)
);

NOR3xp33_ASAP7_75t_L g739 ( 
.A(n_574),
.B(n_25),
.C(n_27),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_499),
.A2(n_25),
.B1(n_29),
.B2(n_32),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_474),
.B(n_61),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_508),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_516),
.Y(n_743)
);

AO221x1_ASAP7_75t_L g744 ( 
.A1(n_460),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.C(n_34),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_570),
.Y(n_745)
);

NOR2x1p5_ASAP7_75t_L g746 ( 
.A(n_506),
.B(n_585),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_474),
.B(n_79),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_516),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_479),
.B(n_77),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_593),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_570),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_524),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_524),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_567),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_479),
.B(n_93),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_570),
.B(n_37),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_479),
.B(n_96),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_571),
.B(n_85),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_562),
.B(n_37),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_479),
.A2(n_97),
.B1(n_131),
.B2(n_123),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_479),
.B(n_134),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_598),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_750),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_715),
.B(n_579),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_705),
.A2(n_514),
.B(n_595),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_634),
.A2(n_537),
.B(n_566),
.C(n_507),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_621),
.B(n_483),
.Y(n_767)
);

BUFx8_ASAP7_75t_L g768 ( 
.A(n_662),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_621),
.B(n_483),
.Y(n_769)
);

AOI21x1_ASAP7_75t_L g770 ( 
.A1(n_608),
.A2(n_537),
.B(n_466),
.Y(n_770)
);

CKINVDCx10_ASAP7_75t_R g771 ( 
.A(n_720),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_636),
.A2(n_571),
.B(n_595),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_616),
.B(n_483),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_754),
.A2(n_567),
.B1(n_587),
.B2(n_582),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_641),
.B(n_715),
.Y(n_775)
);

AO21x1_ASAP7_75t_L g776 ( 
.A1(n_635),
.A2(n_507),
.B(n_466),
.Y(n_776)
);

O2A1O1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_641),
.A2(n_566),
.B(n_581),
.C(n_582),
.Y(n_777)
);

AOI21x1_ASAP7_75t_L g778 ( 
.A1(n_608),
.A2(n_580),
.B(n_503),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_614),
.A2(n_579),
.B1(n_587),
.B2(n_581),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_602),
.A2(n_607),
.B(n_620),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_618),
.B(n_483),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_750),
.Y(n_782)
);

BUFx4f_ASAP7_75t_L g783 ( 
.A(n_734),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_601),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_617),
.Y(n_785)
);

A2O1A1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_630),
.A2(n_578),
.B(n_586),
.C(n_584),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_618),
.B(n_483),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_638),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_619),
.B(n_485),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_750),
.B(n_708),
.Y(n_790)
);

AND2x2_ASAP7_75t_SL g791 ( 
.A(n_754),
.B(n_578),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_750),
.B(n_586),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_602),
.A2(n_577),
.B(n_589),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_675),
.A2(n_594),
.B1(n_573),
.B2(n_485),
.Y(n_794)
);

O2A1O1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_660),
.A2(n_554),
.B(n_555),
.C(n_561),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_619),
.B(n_485),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_607),
.A2(n_589),
.B(n_553),
.Y(n_797)
);

AOI21x1_ASAP7_75t_L g798 ( 
.A1(n_615),
.A2(n_565),
.B(n_584),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_660),
.A2(n_554),
.B(n_561),
.C(n_555),
.Y(n_799)
);

AO21x2_ASAP7_75t_L g800 ( 
.A1(n_637),
.A2(n_485),
.B(n_515),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_702),
.B(n_591),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_620),
.A2(n_589),
.B(n_553),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_628),
.A2(n_589),
.B(n_553),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_630),
.A2(n_521),
.B(n_530),
.C(n_576),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_609),
.B(n_521),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_649),
.A2(n_518),
.B1(n_576),
.B2(n_530),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_610),
.B(n_485),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_610),
.B(n_573),
.Y(n_808)
);

OA21x2_ASAP7_75t_L g809 ( 
.A1(n_632),
.A2(n_515),
.B(n_594),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_628),
.A2(n_553),
.B(n_541),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_626),
.B(n_42),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_645),
.B(n_594),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_645),
.B(n_594),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_623),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_659),
.B(n_594),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_659),
.B(n_573),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_657),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_657),
.A2(n_541),
.B(n_599),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_633),
.B(n_573),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_658),
.B(n_573),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_700),
.B(n_547),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_672),
.B(n_460),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_600),
.A2(n_548),
.B(n_518),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_657),
.A2(n_541),
.B(n_599),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_613),
.B(n_591),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_708),
.B(n_563),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_731),
.B(n_653),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_710),
.A2(n_599),
.B(n_548),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_723),
.B(n_563),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_710),
.A2(n_515),
.B(n_558),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_615),
.A2(n_515),
.B(n_558),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_721),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_612),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_SL g834 ( 
.A(n_699),
.B(n_563),
.C(n_558),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_665),
.B(n_563),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_727),
.B(n_563),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_716),
.A2(n_515),
.B(n_558),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_716),
.A2(n_558),
.B(n_547),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_718),
.B(n_547),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_680),
.A2(n_547),
.B(n_44),
.C(n_45),
.Y(n_840)
);

OAI321xp33_ASAP7_75t_L g841 ( 
.A1(n_740),
.A2(n_42),
.A3(n_49),
.B1(n_50),
.B2(n_52),
.C(n_103),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_758),
.A2(n_110),
.B(n_118),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_667),
.B(n_49),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_629),
.B(n_50),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_668),
.B(n_624),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_719),
.B(n_612),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_642),
.B(n_647),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_721),
.B(n_651),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_680),
.A2(n_759),
.B(n_736),
.C(n_656),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_714),
.B(n_687),
.Y(n_850)
);

OAI321xp33_ASAP7_75t_L g851 ( 
.A1(n_740),
.A2(n_631),
.A3(n_736),
.B1(n_759),
.B2(n_611),
.C(n_646),
.Y(n_851)
);

BUFx12f_ASAP7_75t_L g852 ( 
.A(n_735),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_687),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_762),
.A2(n_612),
.B1(n_622),
.B2(n_663),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_713),
.A2(n_707),
.B(n_688),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_654),
.B(n_690),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_696),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_638),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_697),
.A2(n_689),
.B1(n_670),
.B2(n_655),
.Y(n_859)
);

AOI21x1_ASAP7_75t_L g860 ( 
.A1(n_683),
.A2(n_686),
.B(n_627),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_612),
.A2(n_622),
.B1(n_661),
.B2(n_723),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_622),
.Y(n_862)
);

AND2x2_ASAP7_75t_SL g863 ( 
.A(n_739),
.B(n_760),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_644),
.B(n_643),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_666),
.A2(n_761),
.B(n_757),
.Y(n_865)
);

NOR2x1_ASAP7_75t_L g866 ( 
.A(n_746),
.B(n_704),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_734),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_666),
.A2(n_725),
.B(n_755),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_648),
.A2(n_717),
.B(n_631),
.C(n_684),
.Y(n_869)
);

AOI21xp33_ASAP7_75t_L g870 ( 
.A1(n_604),
.A2(n_625),
.B(n_681),
.Y(n_870)
);

CKINVDCx11_ASAP7_75t_R g871 ( 
.A(n_733),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_741),
.A2(n_747),
.B(n_749),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_622),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_682),
.A2(n_603),
.B(n_703),
.Y(n_874)
);

NAND2x1_ASAP7_75t_L g875 ( 
.A(n_753),
.B(n_730),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_682),
.A2(n_698),
.B(n_606),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_650),
.A2(n_709),
.B(n_732),
.Y(n_877)
);

OAI21x1_ASAP7_75t_L g878 ( 
.A1(n_639),
.A2(n_748),
.B(n_730),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_745),
.A2(n_751),
.B(n_652),
.C(n_692),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_677),
.B(n_679),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_693),
.A2(n_694),
.B1(n_706),
.B2(n_701),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_722),
.A2(n_743),
.B(n_728),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_695),
.A2(n_726),
.B(n_737),
.C(n_738),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_676),
.A2(n_742),
.B(n_752),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_676),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_685),
.A2(n_756),
.B1(n_661),
.B2(n_712),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_678),
.A2(n_729),
.B(n_742),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_SL g888 ( 
.A1(n_684),
.A2(n_673),
.B(n_664),
.C(n_669),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_671),
.A2(n_674),
.B(n_711),
.C(n_724),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_711),
.A2(n_640),
.B(n_720),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_605),
.B(n_734),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_744),
.A2(n_720),
.B(n_691),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_621),
.B(n_633),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_636),
.A2(n_715),
.B1(n_621),
.B2(n_616),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_613),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_617),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_702),
.B(n_714),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_621),
.B(n_616),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_665),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_636),
.A2(n_715),
.B1(n_621),
.B2(n_616),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_705),
.A2(n_475),
.B(n_488),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_636),
.A2(n_614),
.B(n_641),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_609),
.B(n_534),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_621),
.B(n_616),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_705),
.A2(n_475),
.B(n_488),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_754),
.A2(n_641),
.B1(n_675),
.B2(n_535),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_617),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_715),
.B(n_636),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_641),
.A2(n_630),
.B(n_715),
.C(n_618),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_705),
.A2(n_475),
.B(n_488),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_609),
.B(n_534),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_621),
.B(n_616),
.Y(n_912)
);

BUFx12f_ASAP7_75t_L g913 ( 
.A(n_662),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_617),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_641),
.A2(n_630),
.B(n_715),
.C(n_618),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_621),
.B(n_616),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_641),
.A2(n_630),
.B(n_715),
.C(n_618),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_621),
.B(n_616),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_617),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_621),
.B(n_616),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_621),
.B(n_616),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_705),
.A2(n_475),
.B(n_488),
.Y(n_922)
);

O2A1O1Ixp5_ASAP7_75t_L g923 ( 
.A1(n_616),
.A2(n_632),
.B(n_636),
.C(n_635),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_705),
.A2(n_475),
.B(n_488),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_638),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_621),
.B(n_616),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_621),
.B(n_616),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_705),
.A2(n_475),
.B(n_488),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_636),
.A2(n_614),
.B(n_641),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_601),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_617),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_609),
.B(n_626),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_SL g933 ( 
.A1(n_660),
.A2(n_636),
.B(n_616),
.C(n_632),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_621),
.B(n_616),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_621),
.B(n_633),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_638),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_636),
.A2(n_614),
.B(n_641),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_705),
.A2(n_475),
.B(n_488),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_SL g939 ( 
.A(n_735),
.B(n_469),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_621),
.B(n_616),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_641),
.A2(n_630),
.B(n_715),
.C(n_618),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_636),
.A2(n_614),
.B(n_641),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_941),
.A2(n_929),
.B(n_902),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_775),
.B(n_908),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_774),
.A2(n_906),
.B1(n_894),
.B2(n_900),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_867),
.B(n_850),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_878),
.A2(n_765),
.B(n_798),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_846),
.A2(n_839),
.B(n_778),
.Y(n_948)
);

AO21x1_ASAP7_75t_L g949 ( 
.A1(n_937),
.A2(n_942),
.B(n_908),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_774),
.A2(n_906),
.B1(n_918),
.B2(n_920),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_898),
.A2(n_921),
.B1(n_916),
.B2(n_940),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_764),
.A2(n_772),
.B(n_933),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_904),
.B(n_912),
.Y(n_953)
);

OAI21x1_ASAP7_75t_L g954 ( 
.A1(n_874),
.A2(n_876),
.B(n_901),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_905),
.A2(n_922),
.B(n_910),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_871),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_924),
.A2(n_938),
.B(n_928),
.Y(n_957)
);

AOI21xp33_ASAP7_75t_L g958 ( 
.A1(n_851),
.A2(n_848),
.B(n_926),
.Y(n_958)
);

AO31x2_ASAP7_75t_L g959 ( 
.A1(n_776),
.A2(n_786),
.A3(n_804),
.B(n_849),
.Y(n_959)
);

O2A1O1Ixp5_ASAP7_75t_L g960 ( 
.A1(n_870),
.A2(n_923),
.B(n_927),
.C(n_934),
.Y(n_960)
);

BUFx10_ASAP7_75t_L g961 ( 
.A(n_891),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_893),
.B(n_935),
.Y(n_962)
);

AOI21xp33_ASAP7_75t_L g963 ( 
.A1(n_848),
.A2(n_863),
.B(n_844),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_862),
.Y(n_964)
);

AOI21x1_ASAP7_75t_L g965 ( 
.A1(n_846),
.A2(n_839),
.B(n_790),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_884),
.A2(n_887),
.B(n_868),
.Y(n_966)
);

AO21x1_ASAP7_75t_L g967 ( 
.A1(n_767),
.A2(n_769),
.B(n_790),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_864),
.B(n_881),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_850),
.B(n_853),
.Y(n_969)
);

AND3x4_ASAP7_75t_L g970 ( 
.A(n_866),
.B(n_801),
.C(n_897),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_862),
.Y(n_971)
);

BUFx4_ASAP7_75t_SL g972 ( 
.A(n_788),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_832),
.B(n_791),
.Y(n_973)
);

AOI21xp33_ASAP7_75t_L g974 ( 
.A1(n_863),
.A2(n_869),
.B(n_890),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_777),
.A2(n_923),
.B(n_859),
.C(n_889),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_852),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_865),
.A2(n_799),
.B(n_795),
.Y(n_977)
);

OAI22xp33_ASAP7_75t_L g978 ( 
.A1(n_903),
.A2(n_911),
.B1(n_899),
.B2(n_939),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_SL g979 ( 
.A1(n_764),
.A2(n_836),
.B(n_826),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_832),
.B(n_791),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_855),
.A2(n_828),
.B(n_770),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_779),
.A2(n_787),
.B(n_781),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_827),
.B(n_932),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_933),
.A2(n_773),
.B(n_872),
.Y(n_984)
);

INVx5_ASAP7_75t_L g985 ( 
.A(n_817),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_827),
.B(n_932),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_830),
.A2(n_837),
.B(n_802),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_886),
.A2(n_835),
.B1(n_854),
.B2(n_845),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_857),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_812),
.A2(n_816),
.B(n_813),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_807),
.A2(n_796),
.B(n_789),
.Y(n_991)
);

NAND2x1_ASAP7_75t_L g992 ( 
.A(n_763),
.B(n_782),
.Y(n_992)
);

INVxp67_ASAP7_75t_SL g993 ( 
.A(n_862),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_815),
.A2(n_808),
.B(n_766),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_803),
.A2(n_810),
.B(n_838),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_794),
.A2(n_811),
.B1(n_847),
.B2(n_856),
.Y(n_996)
);

OAI21x1_ASAP7_75t_SL g997 ( 
.A1(n_842),
.A2(n_819),
.B(n_831),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_880),
.B(n_805),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_883),
.A2(n_820),
.B(n_888),
.Y(n_999)
);

AOI21xp33_ASAP7_75t_L g1000 ( 
.A1(n_841),
.A2(n_821),
.B(n_822),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_853),
.B(n_895),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_823),
.A2(n_877),
.B(n_882),
.Y(n_1002)
);

NAND3xp33_ASAP7_75t_SL g1003 ( 
.A(n_858),
.B(n_925),
.C(n_936),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_862),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_896),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_805),
.B(n_822),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_907),
.Y(n_1007)
);

NAND3xp33_ASAP7_75t_L g1008 ( 
.A(n_845),
.B(n_895),
.C(n_892),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_780),
.A2(n_792),
.B(n_797),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_794),
.A2(n_840),
.B1(n_930),
.B2(n_814),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_809),
.A2(n_861),
.B(n_793),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_914),
.B(n_931),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_809),
.A2(n_792),
.B(n_800),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_919),
.B(n_885),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_784),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_897),
.B(n_801),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_825),
.Y(n_1017)
);

AO31x2_ASAP7_75t_L g1018 ( 
.A1(n_806),
.A2(n_879),
.A3(n_818),
.B(n_824),
.Y(n_1018)
);

AO21x1_ASAP7_75t_L g1019 ( 
.A1(n_860),
.A2(n_875),
.B(n_829),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_800),
.A2(n_834),
.B(n_763),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_834),
.A2(n_873),
.B(n_833),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_833),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_817),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_891),
.A2(n_783),
.B(n_843),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_913),
.A2(n_771),
.B(n_768),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_768),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_878),
.A2(n_765),
.B(n_798),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_895),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_775),
.A2(n_915),
.B1(n_917),
.B2(n_909),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_862),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_785),
.Y(n_1031)
);

CKINVDCx11_ASAP7_75t_R g1032 ( 
.A(n_871),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_857),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_878),
.A2(n_765),
.B(n_798),
.Y(n_1034)
);

AO31x2_ASAP7_75t_L g1035 ( 
.A1(n_776),
.A2(n_909),
.A3(n_917),
.B(n_915),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_775),
.B(n_908),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_893),
.B(n_935),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_893),
.B(n_935),
.Y(n_1038)
);

O2A1O1Ixp5_ASAP7_75t_L g1039 ( 
.A1(n_909),
.A2(n_917),
.B(n_941),
.C(n_915),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_775),
.B(n_609),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_878),
.A2(n_765),
.B(n_798),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_871),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_878),
.A2(n_765),
.B(n_798),
.Y(n_1043)
);

AO31x2_ASAP7_75t_L g1044 ( 
.A1(n_776),
.A2(n_909),
.A3(n_917),
.B(n_915),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_862),
.Y(n_1045)
);

O2A1O1Ixp5_ASAP7_75t_L g1046 ( 
.A1(n_909),
.A2(n_917),
.B(n_941),
.C(n_915),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_878),
.A2(n_765),
.B(n_798),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_867),
.B(n_850),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_775),
.B(n_609),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_775),
.B(n_908),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_775),
.B(n_908),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_775),
.B(n_908),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_775),
.B(n_908),
.Y(n_1053)
);

OAI33xp33_ASAP7_75t_L g1054 ( 
.A1(n_903),
.A2(n_631),
.A3(n_494),
.B1(n_534),
.B2(n_482),
.B3(n_315),
.Y(n_1054)
);

CKINVDCx6p67_ASAP7_75t_R g1055 ( 
.A(n_871),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_903),
.B(n_911),
.Y(n_1056)
);

NAND2x1_ASAP7_75t_L g1057 ( 
.A(n_763),
.B(n_657),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_862),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_909),
.A2(n_917),
.B(n_915),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_857),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_878),
.A2(n_765),
.B(n_798),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_775),
.B(n_908),
.Y(n_1062)
);

OR2x6_ASAP7_75t_L g1063 ( 
.A(n_852),
.B(n_734),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_785),
.Y(n_1064)
);

AND2x6_ASAP7_75t_L g1065 ( 
.A(n_835),
.B(n_750),
.Y(n_1065)
);

OA21x2_ASAP7_75t_L g1066 ( 
.A1(n_823),
.A2(n_786),
.B(n_878),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_909),
.A2(n_917),
.B(n_915),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_785),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_878),
.A2(n_765),
.B(n_798),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_857),
.Y(n_1070)
);

OAI21xp33_ASAP7_75t_SL g1071 ( 
.A1(n_774),
.A2(n_906),
.B(n_775),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_775),
.A2(n_906),
.B1(n_870),
.B2(n_863),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_909),
.A2(n_917),
.B(n_915),
.Y(n_1073)
);

BUFx10_ASAP7_75t_L g1074 ( 
.A(n_1042),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_962),
.B(n_1037),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_1016),
.B(n_969),
.Y(n_1076)
);

CKINVDCx11_ASAP7_75t_R g1077 ( 
.A(n_1032),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_964),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_1016),
.B(n_969),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_989),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_1055),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1033),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_1026),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_968),
.A2(n_943),
.B(n_1073),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1072),
.A2(n_953),
.B1(n_945),
.B2(n_1029),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_953),
.A2(n_945),
.B1(n_950),
.B2(n_951),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1040),
.A2(n_1038),
.B1(n_951),
.B2(n_950),
.Y(n_1087)
);

AO21x1_ASAP7_75t_L g1088 ( 
.A1(n_958),
.A2(n_974),
.B(n_1067),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_985),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_974),
.A2(n_963),
.B1(n_958),
.B2(n_1054),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_972),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_963),
.A2(n_1071),
.B1(n_986),
.B2(n_983),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_985),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1001),
.B(n_1017),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_1028),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1060),
.Y(n_1096)
);

OR2x6_ASAP7_75t_SL g1097 ( 
.A(n_1008),
.B(n_1056),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_956),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_1063),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_944),
.B(n_1036),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_944),
.B(n_1036),
.Y(n_1101)
);

BUFx2_ASAP7_75t_R g1102 ( 
.A(n_976),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_946),
.B(n_1048),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1070),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_998),
.A2(n_1059),
.B1(n_973),
.B2(n_980),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_1063),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_991),
.A2(n_982),
.B(n_994),
.Y(n_1107)
);

AO21x1_ASAP7_75t_L g1108 ( 
.A1(n_998),
.A2(n_1010),
.B(n_1006),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_961),
.B(n_1015),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_991),
.A2(n_984),
.B(n_990),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1039),
.A2(n_1046),
.B(n_975),
.C(n_978),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_946),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_SL g1113 ( 
.A1(n_1050),
.A2(n_1051),
.B(n_1062),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_1048),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_964),
.Y(n_1115)
);

NOR2x1_ASAP7_75t_R g1116 ( 
.A(n_973),
.B(n_980),
.Y(n_1116)
);

BUFx12f_ASAP7_75t_L g1117 ( 
.A(n_1063),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_961),
.Y(n_1118)
);

BUFx12f_ASAP7_75t_L g1119 ( 
.A(n_1004),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_970),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1004),
.Y(n_1121)
);

NAND2x1_ASAP7_75t_L g1122 ( 
.A(n_1065),
.B(n_971),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1050),
.B(n_1051),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1003),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1052),
.A2(n_1062),
.B1(n_1053),
.B2(n_988),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1052),
.A2(n_1053),
.B1(n_996),
.B2(n_1006),
.Y(n_1126)
);

NAND2xp33_ASAP7_75t_L g1127 ( 
.A(n_1065),
.B(n_985),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_1004),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_960),
.A2(n_1024),
.B(n_1000),
.C(n_996),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_L g1130 ( 
.A(n_1000),
.B(n_1010),
.C(n_999),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_1023),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_952),
.A2(n_979),
.B(n_1002),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_985),
.Y(n_1133)
);

NOR2x1_ASAP7_75t_SL g1134 ( 
.A(n_1022),
.B(n_1021),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1005),
.Y(n_1135)
);

AND2x2_ASAP7_75t_SL g1136 ( 
.A(n_1014),
.B(n_1007),
.Y(n_1136)
);

OA22x2_ASAP7_75t_L g1137 ( 
.A1(n_1025),
.A2(n_993),
.B1(n_1068),
.B2(n_1031),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_955),
.A2(n_957),
.B(n_1011),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1030),
.Y(n_1139)
);

HB1xp67_ASAP7_75t_L g1140 ( 
.A(n_1064),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_949),
.B(n_1044),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_1012),
.B(n_1035),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1011),
.A2(n_966),
.B(n_954),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_1030),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1045),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1035),
.B(n_1044),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1035),
.B(n_1044),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_967),
.A2(n_1065),
.B1(n_997),
.B2(n_1058),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_1045),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1058),
.Y(n_1150)
);

NOR4xp25_ASAP7_75t_L g1151 ( 
.A(n_959),
.B(n_965),
.C(n_1018),
.D(n_977),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1057),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1020),
.A2(n_987),
.B(n_1013),
.Y(n_1153)
);

AND2x2_ASAP7_75t_SL g1154 ( 
.A(n_1066),
.B(n_1065),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_981),
.A2(n_995),
.B(n_1009),
.Y(n_1155)
);

INVx5_ASAP7_75t_L g1156 ( 
.A(n_1065),
.Y(n_1156)
);

BUFx10_ASAP7_75t_L g1157 ( 
.A(n_992),
.Y(n_1157)
);

BUFx12f_ASAP7_75t_L g1158 ( 
.A(n_1019),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1018),
.B(n_948),
.Y(n_1159)
);

OR2x2_ASAP7_75t_L g1160 ( 
.A(n_959),
.B(n_1018),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1066),
.A2(n_947),
.B(n_1069),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_SL g1162 ( 
.A1(n_1034),
.A2(n_1041),
.B1(n_1043),
.B2(n_1047),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1061),
.B(n_962),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1032),
.Y(n_1165)
);

BUFx2_ASAP7_75t_SL g1166 ( 
.A(n_956),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_989),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1072),
.A2(n_775),
.B1(n_906),
.B2(n_909),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_953),
.B(n_951),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_1032),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_1028),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1072),
.A2(n_774),
.B1(n_906),
.B2(n_775),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1028),
.Y(n_1175)
);

OR2x2_ASAP7_75t_SL g1176 ( 
.A(n_1003),
.B(n_534),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_1032),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1056),
.B(n_903),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1016),
.B(n_969),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1040),
.B(n_609),
.Y(n_1182)
);

BUFx4_ASAP7_75t_SL g1183 ( 
.A(n_1026),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1072),
.A2(n_774),
.B1(n_906),
.B2(n_775),
.Y(n_1184)
);

NAND2xp33_ASAP7_75t_L g1185 ( 
.A(n_1072),
.B(n_774),
.Y(n_1185)
);

INVxp67_ASAP7_75t_L g1186 ( 
.A(n_1028),
.Y(n_1186)
);

OR2x6_ASAP7_75t_L g1187 ( 
.A(n_1063),
.B(n_1024),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1016),
.B(n_969),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_964),
.Y(n_1189)
);

INVx4_ASAP7_75t_L g1190 ( 
.A(n_985),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1056),
.B(n_903),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_985),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_962),
.B(n_1037),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1028),
.Y(n_1196)
);

NAND2xp33_ASAP7_75t_L g1197 ( 
.A(n_1072),
.B(n_774),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1016),
.B(n_969),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1056),
.B(n_903),
.Y(n_1199)
);

INVxp67_ASAP7_75t_SL g1200 ( 
.A(n_1140),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_1095),
.Y(n_1201)
);

OAI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1168),
.A2(n_1194),
.B1(n_1164),
.B2(n_1181),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1077),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1185),
.A2(n_1197),
.B1(n_1085),
.B2(n_1184),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1075),
.B(n_1193),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_SL g1206 ( 
.A1(n_1182),
.A2(n_1171),
.B1(n_1180),
.B2(n_1195),
.Y(n_1206)
);

INVx6_ASAP7_75t_L g1207 ( 
.A(n_1119),
.Y(n_1207)
);

BUFx12f_ASAP7_75t_L g1208 ( 
.A(n_1091),
.Y(n_1208)
);

INVx6_ASAP7_75t_L g1209 ( 
.A(n_1156),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1104),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1174),
.B(n_1178),
.Y(n_1211)
);

AO21x2_ASAP7_75t_L g1212 ( 
.A1(n_1138),
.A2(n_1155),
.B(n_1143),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1175),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1082),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1100),
.B(n_1101),
.Y(n_1215)
);

CKINVDCx11_ASAP7_75t_R g1216 ( 
.A(n_1170),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_SL g1217 ( 
.A1(n_1173),
.A2(n_1184),
.B1(n_1085),
.B2(n_1086),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1168),
.A2(n_1173),
.B1(n_1087),
.B2(n_1169),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1156),
.Y(n_1219)
);

BUFx2_ASAP7_75t_R g1220 ( 
.A(n_1081),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_SL g1221 ( 
.A1(n_1086),
.A2(n_1120),
.B1(n_1124),
.B2(n_1130),
.Y(n_1221)
);

INVxp33_ASAP7_75t_L g1222 ( 
.A(n_1191),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1096),
.Y(n_1223)
);

BUFx2_ASAP7_75t_R g1224 ( 
.A(n_1165),
.Y(n_1224)
);

INVx6_ASAP7_75t_L g1225 ( 
.A(n_1190),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1094),
.B(n_1076),
.Y(n_1226)
);

BUFx12f_ASAP7_75t_L g1227 ( 
.A(n_1074),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1167),
.Y(n_1228)
);

AO21x2_ASAP7_75t_L g1229 ( 
.A1(n_1132),
.A2(n_1153),
.B(n_1110),
.Y(n_1229)
);

CKINVDCx6p67_ASAP7_75t_R g1230 ( 
.A(n_1177),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1088),
.A2(n_1090),
.B1(n_1130),
.B2(n_1087),
.Y(n_1231)
);

INVx4_ASAP7_75t_SL g1232 ( 
.A(n_1187),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1108),
.A2(n_1169),
.B1(n_1092),
.B2(n_1105),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1187),
.B(n_1076),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1183),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1187),
.A2(n_1103),
.B1(n_1125),
.B2(n_1079),
.Y(n_1236)
);

CKINVDCx8_ASAP7_75t_R g1237 ( 
.A(n_1166),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1098),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1097),
.A2(n_1199),
.B1(n_1176),
.B2(n_1135),
.Y(n_1239)
);

BUFx8_ASAP7_75t_L g1240 ( 
.A(n_1083),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1103),
.A2(n_1125),
.B1(n_1198),
.B2(n_1079),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1172),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1196),
.Y(n_1243)
);

INVx6_ASAP7_75t_L g1244 ( 
.A(n_1192),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1131),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1106),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1142),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1179),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1179),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1105),
.A2(n_1107),
.B1(n_1126),
.B2(n_1084),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1078),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1145),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1123),
.B(n_1113),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1109),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1186),
.Y(n_1255)
);

BUFx8_ASAP7_75t_SL g1256 ( 
.A(n_1099),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1111),
.A2(n_1129),
.B(n_1126),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1123),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_SL g1259 ( 
.A1(n_1117),
.A2(n_1136),
.B1(n_1118),
.B2(n_1112),
.Y(n_1259)
);

AOI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1188),
.A2(n_1198),
.B1(n_1137),
.B2(n_1114),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1134),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1146),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1188),
.B(n_1116),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1116),
.B(n_1163),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1159),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1102),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1141),
.A2(n_1147),
.B(n_1160),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1089),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1149),
.B(n_1144),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1154),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1139),
.B(n_1144),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1139),
.B(n_1144),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1150),
.B(n_1128),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1150),
.B(n_1133),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1122),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1074),
.Y(n_1276)
);

OA21x2_ASAP7_75t_L g1277 ( 
.A1(n_1148),
.A2(n_1151),
.B(n_1162),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1150),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1133),
.A2(n_1158),
.B1(n_1093),
.B2(n_1152),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1157),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1127),
.A2(n_1152),
.B1(n_1115),
.B2(n_1121),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1115),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1157),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1152),
.A2(n_1121),
.B1(n_1189),
.B2(n_1151),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1121),
.A2(n_775),
.B1(n_1072),
.B2(n_1185),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1189),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1156),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1182),
.A2(n_640),
.B1(n_630),
.B2(n_429),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1080),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1161),
.A2(n_1027),
.B(n_947),
.Y(n_1290)
);

OAI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1168),
.A2(n_775),
.B1(n_851),
.B2(n_1174),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1173),
.A2(n_499),
.B1(n_419),
.B2(n_890),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1119),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1080),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1077),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1080),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1183),
.Y(n_1297)
);

INVx6_ASAP7_75t_L g1298 ( 
.A(n_1119),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1185),
.A2(n_775),
.B1(n_1072),
.B2(n_1197),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1183),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1080),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1080),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1080),
.Y(n_1303)
);

INVx6_ASAP7_75t_L g1304 ( 
.A(n_1119),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1080),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1080),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1095),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1185),
.A2(n_775),
.B1(n_1072),
.B2(n_1197),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1185),
.A2(n_775),
.B1(n_1072),
.B2(n_1197),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1267),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1262),
.B(n_1247),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1267),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1250),
.B(n_1257),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1290),
.A2(n_1250),
.B(n_1261),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1233),
.A2(n_1253),
.B(n_1277),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1270),
.B(n_1217),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1232),
.B(n_1265),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1270),
.B(n_1233),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1292),
.A2(n_1309),
.B1(n_1299),
.B2(n_1308),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1229),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1299),
.A2(n_1309),
.B(n_1308),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1277),
.B(n_1218),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1204),
.A2(n_1206),
.B1(n_1231),
.B2(n_1221),
.Y(n_1323)
);

AO21x2_ASAP7_75t_L g1324 ( 
.A1(n_1212),
.A2(n_1291),
.B(n_1264),
.Y(n_1324)
);

AO21x2_ASAP7_75t_L g1325 ( 
.A1(n_1212),
.A2(n_1291),
.B(n_1202),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1231),
.A2(n_1204),
.B(n_1284),
.Y(n_1326)
);

OR2x6_ASAP7_75t_L g1327 ( 
.A(n_1234),
.B(n_1232),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1209),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1214),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1223),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1277),
.B(n_1258),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1232),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1200),
.Y(n_1333)
);

NAND4xp25_ASAP7_75t_L g1334 ( 
.A(n_1211),
.B(n_1288),
.C(n_1239),
.D(n_1285),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1228),
.Y(n_1335)
);

INVx5_ASAP7_75t_L g1336 ( 
.A(n_1209),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1209),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1245),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1202),
.A2(n_1211),
.B1(n_1222),
.B2(n_1285),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1210),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1215),
.B(n_1236),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1289),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1294),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1296),
.B(n_1301),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1302),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1303),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1260),
.B(n_1275),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1305),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1306),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1254),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1216),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1252),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1222),
.B(n_1205),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1213),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1284),
.B(n_1241),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1219),
.A2(n_1287),
.B(n_1279),
.Y(n_1356)
);

AO21x2_ASAP7_75t_L g1357 ( 
.A1(n_1263),
.A2(n_1274),
.B(n_1280),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1226),
.B(n_1271),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1283),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1268),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1268),
.Y(n_1361)
);

NOR2x1p5_ASAP7_75t_L g1362 ( 
.A(n_1227),
.B(n_1230),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_1216),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1282),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1286),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1281),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1272),
.A2(n_1273),
.B(n_1269),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1225),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1278),
.A2(n_1271),
.B(n_1255),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1225),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1311),
.B(n_1243),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1331),
.B(n_1213),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1323),
.A2(n_1259),
.B1(n_1248),
.B2(n_1249),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1310),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1369),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1331),
.B(n_1271),
.Y(n_1376)
);

NOR2x1_ASAP7_75t_L g1377 ( 
.A(n_1360),
.B(n_1361),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1323),
.A2(n_1201),
.B1(n_1307),
.B2(n_1230),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1312),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1331),
.B(n_1251),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1322),
.B(n_1251),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1322),
.B(n_1315),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1369),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1369),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1322),
.B(n_1315),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1311),
.B(n_1242),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1369),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1327),
.B(n_1246),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1369),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1320),
.B(n_1276),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1321),
.A2(n_1319),
.B(n_1313),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1335),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1324),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1320),
.B(n_1266),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1327),
.B(n_1293),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1338),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1324),
.B(n_1293),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1324),
.B(n_1244),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1338),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1313),
.B(n_1237),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1324),
.B(n_1244),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1325),
.B(n_1237),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1327),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1378),
.A2(n_1319),
.B1(n_1339),
.B2(n_1321),
.Y(n_1404)
);

NAND3xp33_ASAP7_75t_L g1405 ( 
.A(n_1378),
.B(n_1334),
.C(n_1339),
.Y(n_1405)
);

OAI221xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1373),
.A2(n_1334),
.B1(n_1313),
.B2(n_1341),
.C(n_1355),
.Y(n_1406)
);

NAND2xp33_ASAP7_75t_L g1407 ( 
.A(n_1391),
.B(n_1362),
.Y(n_1407)
);

NOR3xp33_ASAP7_75t_L g1408 ( 
.A(n_1391),
.B(n_1366),
.C(n_1341),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1379),
.Y(n_1409)
);

OAI221xp5_ASAP7_75t_L g1410 ( 
.A1(n_1373),
.A2(n_1341),
.B1(n_1366),
.B2(n_1350),
.C(n_1351),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1371),
.B(n_1353),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_SL g1412 ( 
.A1(n_1402),
.A2(n_1355),
.B1(n_1326),
.B2(n_1316),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1395),
.A2(n_1355),
.B1(n_1326),
.B2(n_1347),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1400),
.A2(n_1326),
.B1(n_1350),
.B2(n_1332),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1400),
.B(n_1333),
.C(n_1326),
.Y(n_1415)
);

NAND3xp33_ASAP7_75t_L g1416 ( 
.A(n_1402),
.B(n_1333),
.C(n_1326),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1376),
.B(n_1318),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1402),
.A2(n_1316),
.B(n_1347),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1376),
.B(n_1318),
.Y(n_1419)
);

OAI221xp5_ASAP7_75t_SL g1420 ( 
.A1(n_1393),
.A2(n_1397),
.B1(n_1382),
.B2(n_1385),
.C(n_1316),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1403),
.B(n_1327),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1372),
.B(n_1352),
.Y(n_1422)
);

NAND4xp25_ASAP7_75t_L g1423 ( 
.A(n_1397),
.B(n_1344),
.C(n_1346),
.D(n_1345),
.Y(n_1423)
);

OAI221xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1393),
.A2(n_1327),
.B1(n_1318),
.B2(n_1359),
.C(n_1358),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1372),
.B(n_1357),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1372),
.B(n_1357),
.Y(n_1426)
);

NAND3xp33_ASAP7_75t_L g1427 ( 
.A(n_1393),
.B(n_1359),
.C(n_1340),
.Y(n_1427)
);

AOI221xp5_ASAP7_75t_L g1428 ( 
.A1(n_1397),
.A2(n_1340),
.B1(n_1342),
.B2(n_1343),
.C(n_1349),
.Y(n_1428)
);

NOR3xp33_ASAP7_75t_L g1429 ( 
.A(n_1398),
.B(n_1367),
.C(n_1368),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1376),
.B(n_1325),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1380),
.B(n_1325),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1386),
.B(n_1357),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1386),
.B(n_1357),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1394),
.B(n_1329),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_SL g1435 ( 
.A1(n_1395),
.A2(n_1347),
.B(n_1317),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1394),
.B(n_1396),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1380),
.B(n_1325),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1381),
.B(n_1314),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1394),
.B(n_1330),
.Y(n_1439)
);

NAND3xp33_ASAP7_75t_L g1440 ( 
.A(n_1390),
.B(n_1345),
.C(n_1348),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1392),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1398),
.A2(n_1356),
.B(n_1367),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1381),
.B(n_1382),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1396),
.B(n_1330),
.Y(n_1444)
);

OAI221xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1398),
.A2(n_1327),
.B1(n_1358),
.B2(n_1354),
.C(n_1343),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1395),
.B(n_1388),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1432),
.B(n_1399),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1409),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1421),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1409),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1443),
.B(n_1375),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1441),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1443),
.B(n_1375),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1441),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1433),
.B(n_1399),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1436),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1444),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1431),
.B(n_1383),
.Y(n_1458)
);

INVx4_ASAP7_75t_L g1459 ( 
.A(n_1421),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1405),
.B(n_1354),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1425),
.B(n_1384),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1437),
.B(n_1384),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1440),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1421),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1440),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1438),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1438),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1426),
.B(n_1374),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1437),
.B(n_1387),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1446),
.B(n_1401),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1430),
.B(n_1387),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1427),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1434),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1430),
.B(n_1389),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1405),
.A2(n_1363),
.B1(n_1395),
.B2(n_1347),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1416),
.B(n_1420),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1439),
.Y(n_1477)
);

OAI21xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1476),
.A2(n_1423),
.B(n_1428),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1452),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1450),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1452),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1452),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1463),
.B(n_1417),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1449),
.B(n_1419),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1476),
.B(n_1416),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1450),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1476),
.B(n_1415),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1459),
.B(n_1442),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_SL g1489 ( 
.A(n_1460),
.B(n_1406),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1470),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1463),
.B(n_1419),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1461),
.B(n_1463),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1454),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1449),
.B(n_1429),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1454),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1449),
.B(n_1435),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1460),
.B(n_1363),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1454),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1450),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1461),
.B(n_1415),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1448),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1465),
.B(n_1408),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1461),
.B(n_1423),
.Y(n_1503)
);

INVxp67_ASAP7_75t_SL g1504 ( 
.A(n_1470),
.Y(n_1504)
);

AOI21xp33_ASAP7_75t_L g1505 ( 
.A1(n_1472),
.A2(n_1407),
.B(n_1404),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1464),
.B(n_1435),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1464),
.B(n_1403),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1448),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1465),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1464),
.B(n_1403),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1450),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1464),
.B(n_1418),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1451),
.B(n_1401),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1451),
.B(n_1453),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1465),
.B(n_1411),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1447),
.B(n_1422),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1480),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1480),
.Y(n_1518)
);

OAI21xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1485),
.A2(n_1472),
.B(n_1459),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1506),
.B(n_1459),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1502),
.B(n_1456),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1502),
.B(n_1456),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1497),
.B(n_1363),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_SL g1524 ( 
.A(n_1505),
.B(n_1220),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1489),
.B(n_1473),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1485),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1480),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1489),
.B(n_1505),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1479),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1479),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1509),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1481),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1492),
.B(n_1447),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1481),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1478),
.B(n_1473),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1482),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1509),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1482),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1506),
.B(n_1459),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1493),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1515),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1492),
.B(n_1455),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1486),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1493),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1495),
.Y(n_1545)
);

NAND3xp33_ASAP7_75t_L g1546 ( 
.A(n_1487),
.B(n_1407),
.C(n_1475),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1478),
.A2(n_1414),
.B1(n_1412),
.B2(n_1475),
.Y(n_1547)
);

NAND2x1p5_ASAP7_75t_L g1548 ( 
.A(n_1487),
.B(n_1401),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1495),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1496),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1496),
.B(n_1459),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1515),
.B(n_1473),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1512),
.B(n_1459),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1498),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1486),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1512),
.B(n_1470),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1498),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1501),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1503),
.B(n_1455),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1526),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1529),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1528),
.A2(n_1546),
.B1(n_1547),
.B2(n_1525),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1537),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1529),
.Y(n_1564)
);

AND3x2_ASAP7_75t_L g1565 ( 
.A(n_1524),
.B(n_1490),
.C(n_1504),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1535),
.A2(n_1550),
.B1(n_1410),
.B2(n_1537),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1530),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1521),
.B(n_1503),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1522),
.A2(n_1413),
.B1(n_1500),
.B2(n_1494),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1559),
.B(n_1550),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1531),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1559),
.B(n_1483),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1523),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1541),
.B(n_1203),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1552),
.B(n_1483),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1556),
.A2(n_1500),
.B1(n_1494),
.B2(n_1490),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1530),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1553),
.B(n_1514),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1533),
.B(n_1491),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1532),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1533),
.B(n_1491),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1532),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1548),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_SL g1584 ( 
.A(n_1519),
.B(n_1224),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1542),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1534),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1553),
.B(n_1514),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1548),
.A2(n_1445),
.B1(n_1470),
.B2(n_1424),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1542),
.B(n_1484),
.Y(n_1589)
);

INVx4_ASAP7_75t_L g1590 ( 
.A(n_1517),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1520),
.B(n_1484),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1548),
.B(n_1516),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1520),
.B(n_1516),
.Y(n_1593)
);

AND2x2_ASAP7_75t_SL g1594 ( 
.A(n_1539),
.B(n_1395),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1534),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1560),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1571),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1561),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1590),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1562),
.A2(n_1539),
.B(n_1551),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1566),
.A2(n_1551),
.B1(n_1488),
.B2(n_1470),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1563),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1562),
.B(n_1477),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1563),
.B(n_1477),
.Y(n_1604)
);

INVxp67_ASAP7_75t_SL g1605 ( 
.A(n_1574),
.Y(n_1605)
);

OAI221xp5_ASAP7_75t_L g1606 ( 
.A1(n_1569),
.A2(n_1540),
.B1(n_1544),
.B2(n_1536),
.C(n_1554),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1590),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1584),
.A2(n_1488),
.B1(n_1395),
.B2(n_1510),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1564),
.Y(n_1609)
);

INVxp67_ASAP7_75t_SL g1610 ( 
.A(n_1574),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1588),
.A2(n_1488),
.B1(n_1507),
.B2(n_1510),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1569),
.A2(n_1488),
.B1(n_1467),
.B2(n_1466),
.Y(n_1612)
);

OAI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1576),
.A2(n_1538),
.B1(n_1557),
.B2(n_1545),
.C(n_1549),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1585),
.B(n_1477),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1567),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1573),
.B(n_1203),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1594),
.B(n_1507),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_SL g1618 ( 
.A1(n_1578),
.A2(n_1295),
.B1(n_1238),
.B2(n_1297),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1577),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1580),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1597),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1596),
.B(n_1295),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1619),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1605),
.B(n_1570),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1610),
.B(n_1568),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1602),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1602),
.B(n_1587),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1616),
.B(n_1587),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1616),
.B(n_1591),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1618),
.B(n_1591),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1619),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1599),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1603),
.B(n_1576),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1600),
.B(n_1578),
.Y(n_1634)
);

INVx1_ASAP7_75t_SL g1635 ( 
.A(n_1599),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1607),
.B(n_1578),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1607),
.B(n_1568),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1620),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1617),
.B(n_1594),
.Y(n_1639)
);

AOI221xp5_ASAP7_75t_L g1640 ( 
.A1(n_1633),
.A2(n_1606),
.B1(n_1613),
.B2(n_1612),
.C(n_1601),
.Y(n_1640)
);

AND4x2_ASAP7_75t_L g1641 ( 
.A(n_1626),
.B(n_1565),
.C(n_1611),
.D(n_1590),
.Y(n_1641)
);

OAI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1630),
.A2(n_1608),
.B1(n_1614),
.B2(n_1604),
.C(n_1609),
.Y(n_1642)
);

AOI211xp5_ASAP7_75t_L g1643 ( 
.A1(n_1625),
.A2(n_1598),
.B(n_1615),
.C(n_1617),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1621),
.A2(n_1595),
.B1(n_1586),
.B2(n_1582),
.C(n_1583),
.Y(n_1644)
);

OAI21xp33_ASAP7_75t_L g1645 ( 
.A1(n_1634),
.A2(n_1593),
.B(n_1589),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1635),
.B(n_1575),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1622),
.B(n_1581),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_SL g1648 ( 
.A(n_1624),
.B(n_1592),
.C(n_1238),
.Y(n_1648)
);

AOI222xp33_ASAP7_75t_L g1649 ( 
.A1(n_1637),
.A2(n_1583),
.B1(n_1538),
.B2(n_1545),
.C1(n_1549),
.C2(n_1557),
.Y(n_1649)
);

OAI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1627),
.A2(n_1572),
.B1(n_1579),
.B2(n_1558),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1646),
.Y(n_1651)
);

NOR2x1_ASAP7_75t_L g1652 ( 
.A(n_1648),
.B(n_1622),
.Y(n_1652)
);

NAND4xp75_ASAP7_75t_L g1653 ( 
.A(n_1640),
.B(n_1639),
.C(n_1636),
.D(n_1623),
.Y(n_1653)
);

AOI211x1_ASAP7_75t_L g1654 ( 
.A1(n_1642),
.A2(n_1629),
.B(n_1628),
.C(n_1639),
.Y(n_1654)
);

AND4x1_ASAP7_75t_L g1655 ( 
.A(n_1643),
.B(n_1638),
.C(n_1631),
.D(n_1240),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1647),
.Y(n_1656)
);

NOR3xp33_ASAP7_75t_L g1657 ( 
.A(n_1645),
.B(n_1632),
.C(n_1300),
.Y(n_1657)
);

NOR3x1_ASAP7_75t_L g1658 ( 
.A(n_1641),
.B(n_1235),
.C(n_1632),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1650),
.A2(n_1558),
.B(n_1518),
.Y(n_1659)
);

AOI211x1_ASAP7_75t_L g1660 ( 
.A1(n_1649),
.A2(n_1644),
.B(n_1508),
.C(n_1501),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1648),
.B(n_1208),
.Y(n_1661)
);

AND4x1_ASAP7_75t_L g1662 ( 
.A(n_1658),
.B(n_1240),
.C(n_1256),
.D(n_1227),
.Y(n_1662)
);

NAND5xp2_ASAP7_75t_L g1663 ( 
.A(n_1656),
.B(n_1362),
.C(n_1240),
.D(n_1256),
.E(n_1208),
.Y(n_1663)
);

AND4x2_ASAP7_75t_L g1664 ( 
.A(n_1652),
.B(n_1377),
.C(n_1543),
.D(n_1527),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1661),
.A2(n_1518),
.B(n_1517),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1653),
.A2(n_1555),
.B1(n_1543),
.B2(n_1527),
.Y(n_1666)
);

AND2x2_ASAP7_75t_SL g1667 ( 
.A(n_1657),
.B(n_1207),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1667),
.A2(n_1651),
.B1(n_1659),
.B2(n_1654),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1666),
.A2(n_1655),
.B1(n_1555),
.B2(n_1660),
.Y(n_1669)
);

NOR2x1_ASAP7_75t_L g1670 ( 
.A(n_1663),
.B(n_1486),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1664),
.Y(n_1671)
);

BUFx3_ASAP7_75t_L g1672 ( 
.A(n_1662),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1665),
.A2(n_1207),
.B1(n_1298),
.B2(n_1304),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1668),
.B(n_1457),
.Y(n_1674)
);

NAND4xp25_ASAP7_75t_L g1675 ( 
.A(n_1672),
.B(n_1354),
.C(n_1298),
.D(n_1304),
.Y(n_1675)
);

OAI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1669),
.A2(n_1207),
.B1(n_1298),
.B2(n_1304),
.Y(n_1676)
);

OAI211xp5_ASAP7_75t_L g1677 ( 
.A1(n_1671),
.A2(n_1336),
.B(n_1457),
.C(n_1499),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1673),
.A2(n_1328),
.B1(n_1337),
.B2(n_1513),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1674),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1678),
.B(n_1670),
.Y(n_1680)
);

NOR3xp33_ASAP7_75t_L g1681 ( 
.A(n_1676),
.B(n_1367),
.C(n_1368),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1680),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1679),
.B1(n_1677),
.B2(n_1681),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1683),
.A2(n_1675),
.B1(n_1511),
.B2(n_1499),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1683),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1685),
.B(n_1513),
.Y(n_1686)
);

OA22x2_ASAP7_75t_L g1687 ( 
.A1(n_1684),
.A2(n_1511),
.B1(n_1499),
.B2(n_1508),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1686),
.A2(n_1511),
.B(n_1468),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_SL g1689 ( 
.A(n_1687),
.B(n_1457),
.Y(n_1689)
);

OAI21xp33_ASAP7_75t_L g1690 ( 
.A1(n_1689),
.A2(n_1469),
.B(n_1462),
.Y(n_1690)
);

AOI322xp5_ASAP7_75t_L g1691 ( 
.A1(n_1690),
.A2(n_1688),
.A3(n_1469),
.B1(n_1462),
.B2(n_1474),
.C1(n_1471),
.C2(n_1458),
.Y(n_1691)
);

AOI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1691),
.A2(n_1462),
.B1(n_1469),
.B2(n_1365),
.C(n_1364),
.Y(n_1692)
);

AOI211xp5_ASAP7_75t_L g1693 ( 
.A1(n_1692),
.A2(n_1328),
.B(n_1337),
.C(n_1370),
.Y(n_1693)
);


endmodule