module real_aes_17211_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g105 ( .A(n_0), .B(n_106), .Y(n_105) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_1), .A2(n_32), .B1(n_141), .B2(n_153), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_2), .A2(n_9), .B1(n_520), .B2(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g106 ( .A(n_3), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_4), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_5), .A2(n_10), .B1(n_530), .B2(n_531), .Y(n_529) );
OR2x2_ASAP7_75t_L g113 ( .A(n_6), .B(n_28), .Y(n_113) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_7), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_8), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_11), .B(n_192), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_12), .A2(n_96), .B1(n_189), .B2(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_13), .A2(n_29), .B1(n_543), .B2(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_14), .B(n_192), .Y(n_585) );
OAI21x1_ASAP7_75t_L g136 ( .A1(n_15), .A2(n_43), .B(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_16), .B(n_281), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_17), .Y(n_525) );
INVx1_ASAP7_75t_L g827 ( .A(n_18), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_18), .B(n_828), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_19), .A2(n_36), .B1(n_179), .B2(n_197), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_20), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_21), .A2(n_41), .B1(n_179), .B2(n_520), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_22), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_23), .B(n_543), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_24), .B(n_144), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_25), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_26), .B(n_202), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_27), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_30), .A2(n_80), .B1(n_141), .B2(n_573), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_31), .A2(n_35), .B1(n_141), .B2(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_33), .A2(n_46), .B1(n_520), .B2(n_522), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_34), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_37), .B(n_192), .Y(n_242) );
INVx2_ASAP7_75t_L g832 ( .A(n_38), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_39), .B(n_193), .Y(n_276) );
INVx1_ASAP7_75t_L g111 ( .A(n_40), .Y(n_111) );
BUFx3_ASAP7_75t_L g835 ( .A(n_40), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_42), .B(n_161), .Y(n_283) );
AND2x2_ASAP7_75t_L g181 ( .A(n_44), .B(n_161), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_45), .B(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_47), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_48), .B(n_197), .Y(n_196) );
XNOR2x1_ASAP7_75t_L g122 ( .A(n_49), .B(n_123), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_49), .A2(n_75), .B1(n_845), .B2(n_846), .Y(n_844) );
INVx1_ASAP7_75t_SL g845 ( .A(n_49), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_50), .A2(n_67), .B1(n_197), .B2(n_522), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_51), .A2(n_70), .B1(n_141), .B2(n_533), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_52), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_53), .A2(n_146), .B(n_171), .C(n_172), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_54), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_55), .A2(n_93), .B1(n_520), .B2(n_531), .Y(n_594) );
INVx1_ASAP7_75t_L g137 ( .A(n_56), .Y(n_137) );
AND2x4_ASAP7_75t_L g158 ( .A(n_57), .B(n_159), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_58), .A2(n_59), .B1(n_179), .B2(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_60), .B(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_61), .B(n_161), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_62), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_63), .B(n_179), .Y(n_245) );
INVx1_ASAP7_75t_L g159 ( .A(n_64), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_65), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_66), .B(n_202), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_68), .B(n_141), .Y(n_140) );
NAND3xp33_ASAP7_75t_L g277 ( .A(n_69), .B(n_153), .C(n_193), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_71), .B(n_141), .Y(n_223) );
INVx2_ASAP7_75t_L g148 ( .A(n_72), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_73), .B(n_192), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_74), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g846 ( .A(n_75), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_75), .B(n_875), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_76), .B(n_199), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_77), .A2(n_92), .B1(n_171), .B2(n_179), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_78), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_79), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_81), .A2(n_87), .B1(n_144), .B2(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_82), .B(n_192), .Y(n_191) );
NAND2xp33_ASAP7_75t_SL g215 ( .A(n_83), .B(n_198), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_84), .B(n_190), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g855 ( .A(n_85), .Y(n_855) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_86), .B(n_202), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_88), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_89), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g121 ( .A(n_89), .Y(n_121) );
NAND2xp33_ASAP7_75t_L g588 ( .A(n_90), .B(n_192), .Y(n_588) );
NAND2xp33_ASAP7_75t_L g224 ( .A(n_91), .B(n_198), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_94), .B(n_161), .Y(n_160) );
NAND3xp33_ASAP7_75t_L g211 ( .A(n_95), .B(n_198), .C(n_210), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_97), .B(n_141), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_98), .B(n_144), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_114), .B(n_862), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx2_ASAP7_75t_SL g871 ( .A(n_105), .Y(n_871) );
INVx5_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx4_ASAP7_75t_L g850 ( .A(n_108), .Y(n_850) );
INVx3_ASAP7_75t_L g872 ( .A(n_108), .Y(n_872) );
AND2x6_ASAP7_75t_SL g108 ( .A(n_109), .B(n_112), .Y(n_108) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_112), .B(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NOR2x1_ASAP7_75t_L g861 ( .A(n_113), .B(n_835), .Y(n_861) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g115 ( .A(n_116), .B(n_839), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_826), .B1(n_836), .B2(n_837), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B(n_504), .Y(n_117) );
AOI21x1_ASAP7_75t_L g838 ( .A1(n_118), .A2(n_122), .B(n_504), .Y(n_838) );
INVx3_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx8_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g860 ( .A(n_120), .B(n_861), .Y(n_860) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g508 ( .A(n_121), .Y(n_508) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g847 ( .A(n_124), .Y(n_847) );
NAND2x1p5_ASAP7_75t_L g124 ( .A(n_125), .B(n_399), .Y(n_124) );
NOR2x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_334), .Y(n_125) );
NAND3xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_257), .C(n_307), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_182), .B(n_217), .C(n_234), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OR2x2_ASAP7_75t_L g473 ( .A(n_129), .B(n_392), .Y(n_473) );
OR2x2_ASAP7_75t_L g484 ( .A(n_129), .B(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_130), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g375 ( .A(n_130), .B(n_264), .Y(n_375) );
AND2x2_ASAP7_75t_L g496 ( .A(n_130), .B(n_306), .Y(n_496) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_162), .Y(n_130) );
INVx2_ASAP7_75t_L g326 ( .A(n_131), .Y(n_326) );
AND2x2_ASAP7_75t_L g341 ( .A(n_131), .B(n_293), .Y(n_341) );
AND2x2_ASAP7_75t_L g350 ( .A(n_131), .B(n_219), .Y(n_350) );
AND2x2_ASAP7_75t_L g419 ( .A(n_131), .B(n_305), .Y(n_419) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g232 ( .A(n_132), .Y(n_232) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_138), .B(n_160), .Y(n_132) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_133), .A2(n_186), .B(n_201), .Y(n_185) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_133), .A2(n_186), .B(n_201), .Y(n_300) );
OAI21xp33_ASAP7_75t_SL g391 ( .A1(n_133), .A2(n_138), .B(n_160), .Y(n_391) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g161 ( .A(n_134), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_134), .B(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_134), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
INVx2_ASAP7_75t_L g256 ( .A(n_135), .Y(n_256) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_136), .Y(n_203) );
OAI21x1_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_149), .B(n_157), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_143), .B(n_146), .Y(n_139) );
OAI22xp33_ASAP7_75t_L g177 ( .A1(n_141), .A2(n_178), .B1(n_179), .B2(n_180), .Y(n_177) );
INVx1_ASAP7_75t_L g522 ( .A(n_141), .Y(n_522) );
INVx1_ASAP7_75t_L g531 ( .A(n_141), .Y(n_531) );
INVx4_ASAP7_75t_L g533 ( .A(n_141), .Y(n_533) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g145 ( .A(n_142), .Y(n_145) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
INVx1_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
INVx2_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_142), .Y(n_179) );
INVx1_ASAP7_75t_L g190 ( .A(n_142), .Y(n_190) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_142), .Y(n_192) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_142), .Y(n_198) );
INVx1_ASAP7_75t_L g214 ( .A(n_142), .Y(n_214) );
INVx1_ASAP7_75t_L g253 ( .A(n_142), .Y(n_253) );
INVx1_ASAP7_75t_L g530 ( .A(n_144), .Y(n_530) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_146), .A2(n_213), .B(n_215), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_146), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_146), .A2(n_241), .B(n_242), .Y(n_240) );
BUFx4f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
BUFx8_ASAP7_75t_L g193 ( .A(n_148), .Y(n_193) );
INVx1_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_154), .Y(n_149) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g200 ( .A(n_156), .Y(n_200) );
OAI21x1_ASAP7_75t_L g186 ( .A1(n_157), .A2(n_187), .B(n_194), .Y(n_186) );
OAI21x1_ASAP7_75t_L g207 ( .A1(n_157), .A2(n_208), .B(n_212), .Y(n_207) );
AND2x4_ASAP7_75t_SL g229 ( .A(n_157), .B(n_203), .Y(n_229) );
OAI21x1_ASAP7_75t_L g239 ( .A1(n_157), .A2(n_240), .B(n_243), .Y(n_239) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_157), .A2(n_275), .B(n_278), .Y(n_274) );
BUFx10_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx10_ASAP7_75t_L g168 ( .A(n_158), .Y(n_168) );
INVx1_ASAP7_75t_L g557 ( .A(n_158), .Y(n_557) );
AND2x2_ASAP7_75t_L g390 ( .A(n_162), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g233 ( .A(n_163), .B(n_205), .Y(n_233) );
INVx2_ASAP7_75t_L g262 ( .A(n_163), .Y(n_262) );
AOI21x1_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_169), .B(n_181), .Y(n_163) );
NOR2xp67_ASAP7_75t_SL g164 ( .A(n_165), .B(n_167), .Y(n_164) );
INVx2_ASAP7_75t_L g523 ( .A(n_165), .Y(n_523) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AO31x2_ASAP7_75t_L g247 ( .A1(n_166), .A2(n_168), .A3(n_248), .B(n_254), .Y(n_247) );
NOR2xp33_ASAP7_75t_SL g536 ( .A(n_166), .B(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_166), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g517 ( .A(n_167), .Y(n_517) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AO31x2_ASAP7_75t_L g527 ( .A1(n_168), .A2(n_528), .A3(n_535), .B(n_536), .Y(n_527) );
AO31x2_ASAP7_75t_L g540 ( .A1(n_168), .A2(n_541), .A3(n_547), .B(n_548), .Y(n_540) );
AO31x2_ASAP7_75t_L g603 ( .A1(n_168), .A2(n_604), .A3(n_607), .B(n_608), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_175), .Y(n_169) );
INVx1_ASAP7_75t_L g227 ( .A(n_171), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVx2_ASAP7_75t_SL g573 ( .A(n_174), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_176), .A2(n_249), .B1(n_251), .B2(n_252), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_176), .A2(n_251), .B1(n_519), .B2(n_521), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_176), .A2(n_251), .B1(n_542), .B2(n_545), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_176), .A2(n_251), .B1(n_554), .B2(n_555), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_176), .A2(n_251), .B1(n_605), .B2(n_606), .Y(n_604) );
INVx2_ASAP7_75t_L g250 ( .A(n_179), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_179), .A2(n_276), .B(n_277), .Y(n_275) );
AND2x2_ASAP7_75t_L g427 ( .A(n_182), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OR2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_204), .Y(n_183) );
INVx1_ASAP7_75t_L g447 ( .A(n_184), .Y(n_447) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g285 ( .A(n_185), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g368 ( .A(n_185), .B(n_273), .Y(n_368) );
O2A1O1Ixp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_191), .C(n_193), .Y(n_187) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_192), .A2(n_209), .B(n_211), .Y(n_208) );
INVx1_ASAP7_75t_L g281 ( .A(n_192), .Y(n_281) );
INVx3_ASAP7_75t_L g520 ( .A(n_192), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_193), .A2(n_244), .B(n_245), .Y(n_243) );
INVx6_ASAP7_75t_L g251 ( .A(n_193), .Y(n_251) );
O2A1O1Ixp5_ASAP7_75t_L g583 ( .A1(n_193), .A2(n_533), .B(n_584), .C(n_585), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_199), .Y(n_194) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g543 ( .A(n_198), .Y(n_543) );
INVx2_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_200), .A2(n_226), .B1(n_227), .B2(n_228), .Y(n_225) );
INVx2_ASAP7_75t_L g607 ( .A(n_202), .Y(n_607) );
INVx4_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_SL g206 ( .A(n_203), .Y(n_206) );
INVx2_ASAP7_75t_L g238 ( .A(n_203), .Y(n_238) );
BUFx3_ASAP7_75t_L g547 ( .A(n_203), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_203), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_SL g581 ( .A(n_203), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_203), .B(n_597), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_203), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g294 ( .A(n_204), .B(n_232), .Y(n_294) );
INVxp67_ASAP7_75t_L g443 ( .A(n_204), .Y(n_443) );
OR2x2_ASAP7_75t_L g485 ( .A(n_204), .B(n_219), .Y(n_485) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g266 ( .A(n_205), .Y(n_266) );
OAI21x1_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_216), .Y(n_205) );
INVx1_ASAP7_75t_L g282 ( .A(n_210), .Y(n_282) );
INVx1_ASAP7_75t_SL g534 ( .A(n_210), .Y(n_534) );
INVx1_ASAP7_75t_L g575 ( .A(n_210), .Y(n_575) );
INVx1_ASAP7_75t_L g544 ( .A(n_214), .Y(n_544) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_230), .Y(n_217) );
INVx1_ASAP7_75t_L g340 ( .A(n_218), .Y(n_340) );
AND2x2_ASAP7_75t_L g494 ( .A(n_218), .B(n_390), .Y(n_494) );
BUFx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g265 ( .A(n_219), .Y(n_265) );
INVx4_ASAP7_75t_L g305 ( .A(n_219), .Y(n_305) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
OAI21x1_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_225), .B(n_229), .Y(n_221) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
AND2x2_ASAP7_75t_L g321 ( .A(n_231), .B(n_304), .Y(n_321) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g358 ( .A(n_232), .B(n_306), .Y(n_358) );
INVx2_ASAP7_75t_L g324 ( .A(n_233), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_233), .B(n_329), .Y(n_492) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_236), .B(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g477 ( .A(n_236), .Y(n_477) );
AND2x2_ASAP7_75t_L g491 ( .A(n_236), .B(n_313), .Y(n_491) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_247), .Y(n_236) );
INVx1_ASAP7_75t_L g271 ( .A(n_237), .Y(n_271) );
AND2x2_ASAP7_75t_L g426 ( .A(n_237), .B(n_333), .Y(n_426) );
OR2x2_ASAP7_75t_L g463 ( .A(n_237), .B(n_247), .Y(n_463) );
OAI21x1_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_246), .Y(n_237) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_238), .A2(n_274), .B(n_283), .Y(n_273) );
OA21x2_ASAP7_75t_L g286 ( .A1(n_238), .A2(n_274), .B(n_283), .Y(n_286) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_238), .A2(n_239), .B(n_246), .Y(n_289) );
AND2x2_ASAP7_75t_L g272 ( .A(n_247), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g287 ( .A(n_247), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g333 ( .A(n_247), .Y(n_333) );
OR2x2_ASAP7_75t_L g346 ( .A(n_247), .B(n_286), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_247), .B(n_286), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_251), .A2(n_529), .B1(n_532), .B2(n_534), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_251), .A2(n_572), .B1(n_574), .B2(n_575), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_251), .A2(n_587), .B(n_588), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_251), .A2(n_534), .B1(n_594), .B2(n_595), .Y(n_593) );
INVx1_ASAP7_75t_L g546 ( .A(n_253), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
BUFx2_ASAP7_75t_L g535 ( .A(n_256), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_267), .B(n_290), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AOI31xp33_ASAP7_75t_L g336 ( .A1(n_259), .A2(n_337), .A3(n_339), .B(n_342), .Y(n_336) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
AND2x2_ASAP7_75t_L g349 ( .A(n_260), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g359 ( .A(n_261), .Y(n_359) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_261), .Y(n_365) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g293 ( .A(n_262), .Y(n_293) );
AND2x2_ASAP7_75t_L g322 ( .A(n_262), .B(n_306), .Y(n_322) );
INVx2_ASAP7_75t_L g372 ( .A(n_262), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_263), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g397 ( .A(n_264), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g446 ( .A(n_264), .B(n_447), .Y(n_446) );
AOI33xp33_ASAP7_75t_L g501 ( .A1(n_264), .A2(n_331), .A3(n_341), .B1(n_368), .B2(n_477), .B3(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g306 ( .A(n_266), .Y(n_306) );
INVx1_ASAP7_75t_L g393 ( .A(n_266), .Y(n_393) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_284), .Y(n_268) );
INVx2_ASAP7_75t_L g301 ( .A(n_269), .Y(n_301) );
AND2x2_ASAP7_75t_L g382 ( .A(n_269), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
INVx1_ASAP7_75t_L g344 ( .A(n_270), .Y(n_344) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g412 ( .A(n_271), .B(n_299), .Y(n_412) );
AND2x2_ASAP7_75t_L g362 ( .A(n_272), .B(n_356), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_272), .B(n_380), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_272), .B(n_412), .Y(n_461) );
AND2x2_ASAP7_75t_L g298 ( .A(n_273), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g317 ( .A(n_273), .B(n_312), .Y(n_317) );
INVx1_ASAP7_75t_L g332 ( .A(n_273), .Y(n_332) );
AOI21x1_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B(n_282), .Y(n_278) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_L g387 ( .A(n_285), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_285), .B(n_480), .Y(n_482) );
AND2x2_ASAP7_75t_L g495 ( .A(n_285), .B(n_311), .Y(n_495) );
AND2x2_ASAP7_75t_L g313 ( .A(n_286), .B(n_299), .Y(n_313) );
INVx2_ASAP7_75t_L g295 ( .A(n_287), .Y(n_295) );
AND2x2_ASAP7_75t_L g409 ( .A(n_287), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g468 ( .A(n_287), .B(n_380), .Y(n_468) );
BUFx2_ASAP7_75t_L g450 ( .A(n_288), .Y(n_450) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx3_ASAP7_75t_L g312 ( .A(n_289), .Y(n_312) );
OAI32xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_295), .A3(n_296), .B1(n_301), .B2(n_302), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g398 ( .A(n_293), .Y(n_398) );
AND2x2_ASAP7_75t_L g428 ( .A(n_293), .B(n_350), .Y(n_428) );
AND2x2_ASAP7_75t_L g370 ( .A(n_294), .B(n_371), .Y(n_370) );
AND3x2_ASAP7_75t_L g377 ( .A(n_294), .B(n_304), .C(n_372), .Y(n_377) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_297), .A2(n_319), .B1(n_328), .B2(n_330), .Y(n_327) );
OAI322xp33_ASAP7_75t_L g475 ( .A1(n_297), .A2(n_396), .A3(n_476), .B1(n_477), .B2(n_478), .C1(n_479), .C2(n_482), .Y(n_475) );
INVx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g497 ( .A(n_298), .B(n_480), .Y(n_497) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_299), .Y(n_316) );
INVxp67_ASAP7_75t_SL g356 ( .A(n_299), .Y(n_356) );
BUFx3_ASAP7_75t_L g380 ( .A(n_299), .Y(n_380) );
INVx1_ASAP7_75t_L g406 ( .A(n_299), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_299), .Y(n_410) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g364 ( .A(n_303), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx1_ASAP7_75t_L g415 ( .A(n_304), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_304), .B(n_372), .Y(n_466) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2x1_ASAP7_75t_L g325 ( .A(n_305), .B(n_326), .Y(n_325) );
BUFx2_ASAP7_75t_L g329 ( .A(n_305), .Y(n_329) );
AND2x2_ASAP7_75t_L g371 ( .A(n_305), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g392 ( .A(n_305), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_306), .B(n_419), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_314), .B(n_318), .C(n_327), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AOI31xp33_ASAP7_75t_L g469 ( .A1(n_309), .A2(n_470), .A3(n_472), .B(n_473), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
AND2x4_ASAP7_75t_L g422 ( .A(n_310), .B(n_331), .Y(n_422) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_311), .Y(n_354) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp67_ASAP7_75t_L g438 ( .A(n_312), .B(n_332), .Y(n_438) );
BUFx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2x1_ASAP7_75t_L g318 ( .A(n_319), .B(n_323), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g478 ( .A(n_321), .Y(n_478) );
AND2x2_ASAP7_75t_L g338 ( .A(n_322), .B(n_329), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_323), .A2(n_408), .B1(n_411), .B2(n_413), .Y(n_407) );
OR2x6_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_SL g465 ( .A(n_326), .Y(n_465) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g435 ( .A(n_331), .B(n_380), .Y(n_435) );
INVx2_ASAP7_75t_L g481 ( .A(n_331), .Y(n_481) );
AND2x4_ASAP7_75t_L g489 ( .A(n_331), .B(n_410), .Y(n_489) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NAND3xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_351), .C(n_381), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_347), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_338), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AND2x4_ASAP7_75t_L g402 ( .A(n_340), .B(n_357), .Y(n_402) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_343), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AND2x2_ASAP7_75t_L g433 ( .A(n_345), .B(n_412), .Y(n_433) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_346), .Y(n_353) );
INVx1_ASAP7_75t_L g471 ( .A(n_346), .Y(n_471) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g500 ( .A(n_349), .Y(n_500) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_350), .Y(n_385) );
AOI211xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_357), .B(n_360), .C(n_373), .Y(n_351) );
NOR3x1_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .C(n_355), .Y(n_352) );
NAND2x1_ASAP7_75t_L g421 ( .A(n_355), .B(n_422), .Y(n_421) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2x1p5_ASAP7_75t_SL g357 ( .A(n_358), .B(n_359), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B1(n_366), .B2(n_369), .Y(n_360) );
INVxp67_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g454 ( .A(n_365), .Y(n_454) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g449 ( .A(n_368), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g503 ( .A(n_371), .Y(n_503) );
AOI21xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B(n_378), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g457 ( .A(n_378), .Y(n_457) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx2_ASAP7_75t_L g384 ( .A(n_380), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_380), .B(n_438), .Y(n_437) );
AOI21xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_385), .B(n_386), .Y(n_381) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_384), .B(n_471), .Y(n_470) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_394), .B2(n_396), .Y(n_386) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g414 ( .A(n_390), .B(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g431 ( .A(n_391), .Y(n_431) );
INVx1_ASAP7_75t_L g451 ( .A(n_392), .Y(n_451) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NOR2x1_ASAP7_75t_L g399 ( .A(n_400), .B(n_455), .Y(n_399) );
NAND3xp33_ASAP7_75t_SL g400 ( .A(n_401), .B(n_416), .C(n_429), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_407), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g462 ( .A(n_405), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2x1p5_ASAP7_75t_L g459 ( .A(n_414), .B(n_442), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .B1(n_423), .B2(n_427), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g472 ( .A(n_422), .Y(n_472) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI21xp33_ASAP7_75t_L g444 ( .A1(n_424), .A2(n_445), .B(n_448), .Y(n_444) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_440), .B1(n_444), .B2(n_452), .Y(n_429) );
OAI21xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B(n_434), .Y(n_430) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B(n_439), .Y(n_434) );
INVx1_ASAP7_75t_L g499 ( .A(n_435), .Y(n_499) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g488 ( .A(n_438), .Y(n_488) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_451), .Y(n_448) );
INVx2_ASAP7_75t_L g480 ( .A(n_450), .Y(n_480) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_474), .Y(n_455) );
AOI211xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B(n_460), .C(n_469), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B(n_464), .C(n_467), .Y(n_460) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_483), .C(n_498), .Y(n_474) );
OR2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_486), .B1(n_490), .B2(n_492), .C(n_493), .Y(n_483) );
NOR2xp67_ASAP7_75t_L g486 ( .A(n_487), .B(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_493) );
OAI21xp33_ASAP7_75t_SL g498 ( .A1(n_499), .A2(n_500), .B(n_501), .Y(n_498) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NOR2xp67_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_735), .Y(n_509) );
NOR2x1_ASAP7_75t_L g510 ( .A(n_511), .B(n_674), .Y(n_510) );
NAND4xp25_ASAP7_75t_L g511 ( .A(n_512), .B(n_625), .C(n_644), .D(n_655), .Y(n_511) );
O2A1O1Ixp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_560), .B(n_567), .C(n_598), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_538), .Y(n_513) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_514), .B(n_690), .C(n_691), .Y(n_689) );
AND2x2_ASAP7_75t_L g771 ( .A(n_514), .B(n_653), .Y(n_771) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_526), .Y(n_514) );
AND2x2_ASAP7_75t_L g615 ( .A(n_515), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g633 ( .A(n_515), .B(n_634), .Y(n_633) );
INVx3_ASAP7_75t_L g650 ( .A(n_515), .Y(n_650) );
AND2x2_ASAP7_75t_L g695 ( .A(n_515), .B(n_540), .Y(n_695) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g564 ( .A(n_516), .Y(n_564) );
AND2x4_ASAP7_75t_L g643 ( .A(n_516), .B(n_634), .Y(n_643) );
AO31x2_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .A3(n_523), .B(n_524), .Y(n_516) );
AO31x2_ASAP7_75t_L g592 ( .A1(n_517), .A2(n_535), .A3(n_593), .B(n_596), .Y(n_592) );
AO31x2_ASAP7_75t_L g552 ( .A1(n_523), .A2(n_553), .A3(n_556), .B(n_558), .Y(n_552) );
AND2x2_ASAP7_75t_L g565 ( .A(n_526), .B(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g618 ( .A(n_526), .B(n_619), .Y(n_618) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_526), .Y(n_641) );
INVx1_ASAP7_75t_L g652 ( .A(n_526), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_526), .B(n_550), .Y(n_661) );
INVx2_ASAP7_75t_L g668 ( .A(n_526), .Y(n_668) );
INVx4_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g613 ( .A(n_527), .B(n_540), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_527), .B(n_620), .Y(n_686) );
AND2x2_ASAP7_75t_L g694 ( .A(n_527), .B(n_552), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_527), .B(n_741), .Y(n_740) );
BUFx2_ASAP7_75t_L g747 ( .A(n_527), .Y(n_747) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g763 ( .A(n_539), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_550), .Y(n_539) );
INVx1_ASAP7_75t_L g566 ( .A(n_540), .Y(n_566) );
INVx1_ASAP7_75t_L g620 ( .A(n_540), .Y(n_620) );
INVx2_ASAP7_75t_L g654 ( .A(n_540), .Y(n_654) );
OR2x2_ASAP7_75t_L g658 ( .A(n_540), .B(n_552), .Y(n_658) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_540), .Y(n_707) );
AO31x2_ASAP7_75t_L g570 ( .A1(n_547), .A2(n_556), .A3(n_571), .B(n_576), .Y(n_570) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g680 ( .A(n_551), .B(n_564), .Y(n_680) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_552), .Y(n_616) );
INVx2_ASAP7_75t_L g634 ( .A(n_552), .Y(n_634) );
AND2x4_ASAP7_75t_L g653 ( .A(n_552), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g741 ( .A(n_552), .Y(n_741) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g589 ( .A(n_557), .Y(n_589) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g659 ( .A(n_563), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_563), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g722 ( .A(n_564), .Y(n_722) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2x1_ASAP7_75t_L g568 ( .A(n_569), .B(n_578), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_569), .B(n_579), .Y(n_672) );
INVx1_ASAP7_75t_L g770 ( .A(n_569), .Y(n_770) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g610 ( .A(n_570), .B(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g624 ( .A(n_570), .B(n_603), .Y(n_624) );
AND2x4_ASAP7_75t_L g647 ( .A(n_570), .B(n_591), .Y(n_647) );
INVx2_ASAP7_75t_L g664 ( .A(n_570), .Y(n_664) );
AND2x2_ASAP7_75t_L g690 ( .A(n_570), .B(n_592), .Y(n_690) );
INVx1_ASAP7_75t_L g755 ( .A(n_570), .Y(n_755) );
AND2x2_ASAP7_75t_L g715 ( .A(n_578), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_591), .Y(n_578) );
AND2x2_ASAP7_75t_L g681 ( .A(n_579), .B(n_638), .Y(n_681) );
AND2x4_ASAP7_75t_L g697 ( .A(n_579), .B(n_664), .Y(n_697) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx2_ASAP7_75t_L g691 ( .A(n_580), .Y(n_691) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B(n_590), .Y(n_580) );
OAI21x1_ASAP7_75t_L g612 ( .A1(n_581), .A2(n_582), .B(n_590), .Y(n_612) );
OAI21x1_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_586), .B(n_589), .Y(n_582) );
INVx2_ASAP7_75t_L g623 ( .A(n_591), .Y(n_623) );
INVx3_ASAP7_75t_L g629 ( .A(n_591), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_591), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_591), .B(n_758), .Y(n_757) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g663 ( .A(n_592), .B(n_664), .Y(n_663) );
BUFx2_ASAP7_75t_L g787 ( .A(n_592), .Y(n_787) );
OAI33xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_613), .A3(n_614), .B1(n_615), .B2(n_617), .B3(n_621), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_601), .B(n_610), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g721 ( .A(n_602), .B(n_722), .Y(n_721) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g630 ( .A(n_603), .B(n_612), .Y(n_630) );
INVx2_ASAP7_75t_L g638 ( .A(n_603), .Y(n_638) );
INVx1_ASAP7_75t_L g646 ( .A(n_603), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_610), .A2(n_666), .B1(n_669), .B2(n_673), .Y(n_665) );
OR2x2_ASAP7_75t_L g805 ( .A(n_610), .B(n_623), .Y(n_805) );
AND2x4_ASAP7_75t_L g709 ( .A(n_611), .B(n_671), .Y(n_709) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_612), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_613), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g673 ( .A(n_613), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_613), .B(n_649), .Y(n_751) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g724 ( .A(n_615), .Y(n_724) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g782 ( .A(n_618), .B(n_650), .Y(n_782) );
NAND2x1_ASAP7_75t_L g800 ( .A(n_618), .B(n_649), .Y(n_800) );
AND2x2_ASAP7_75t_L g824 ( .A(n_618), .B(n_643), .Y(n_824) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g814 ( .A(n_622), .B(n_691), .Y(n_814) );
NOR2x1p5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g748 ( .A(n_623), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g716 ( .A(n_624), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_631), .B1(n_635), .B2(n_639), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
AND2x2_ASAP7_75t_L g723 ( .A(n_628), .B(n_691), .Y(n_723) );
AND2x2_ASAP7_75t_L g760 ( .A(n_628), .B(n_709), .Y(n_760) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_L g635 ( .A(n_629), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_629), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g801 ( .A(n_629), .B(n_630), .Y(n_801) );
AND2x2_ASAP7_75t_L g662 ( .A(n_630), .B(n_663), .Y(n_662) );
AND2x4_ASAP7_75t_L g781 ( .A(n_630), .B(n_647), .Y(n_781) );
AND2x2_ASAP7_75t_L g825 ( .A(n_630), .B(n_690), .Y(n_825) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI222xp33_ASAP7_75t_L g759 ( .A1(n_635), .A2(n_760), .B1(n_761), .B2(n_764), .C1(n_766), .C2(n_767), .Y(n_759) );
AND2x2_ASAP7_75t_L g682 ( .A(n_636), .B(n_650), .Y(n_682) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g713 ( .A(n_637), .Y(n_713) );
INVxp67_ASAP7_75t_SL g758 ( .A(n_637), .Y(n_758) );
INVx2_ASAP7_75t_L g671 ( .A(n_638), .Y(n_671) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g728 ( .A(n_641), .Y(n_728) );
INVx2_ASAP7_75t_L g734 ( .A(n_642), .Y(n_734) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x4_ASAP7_75t_L g718 ( .A(n_643), .B(n_707), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_648), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
AND2x4_ASAP7_75t_L g749 ( .A(n_646), .B(n_697), .Y(n_749) );
INVx2_ASAP7_75t_L g796 ( .A(n_646), .Y(n_796) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVx4_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g739 ( .A(n_650), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g773 ( .A(n_650), .B(n_658), .Y(n_773) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g678 ( .A(n_652), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_653), .B(n_743), .Y(n_742) );
AND2x4_ASAP7_75t_L g785 ( .A(n_653), .B(n_701), .Y(n_785) );
O2A1O1Ixp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_660), .B(n_662), .C(n_665), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
OR2x2_ASAP7_75t_L g666 ( .A(n_658), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g702 ( .A(n_658), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_659), .B(n_694), .Y(n_798) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g774 ( .A(n_661), .B(n_743), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_663), .B(n_713), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_663), .A2(n_679), .B1(n_721), .B2(n_723), .Y(n_720) );
AND2x2_ASAP7_75t_L g726 ( .A(n_663), .B(n_691), .Y(n_726) );
AND2x2_ASAP7_75t_L g795 ( .A(n_663), .B(n_796), .Y(n_795) );
O2A1O1Ixp33_ASAP7_75t_L g788 ( .A1(n_666), .A2(n_768), .B(n_789), .C(n_792), .Y(n_788) );
INVx2_ASAP7_75t_L g701 ( .A(n_668), .Y(n_701) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx1_ASAP7_75t_L g779 ( .A(n_671), .Y(n_779) );
INVx1_ASAP7_75t_L g704 ( .A(n_672), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_673), .A2(n_720), .B1(n_724), .B2(n_725), .Y(n_719) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_687), .C(n_710), .Y(n_674) );
AO22x1_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_681), .B1(n_682), .B2(n_683), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_680), .Y(n_813) );
OR2x2_ASAP7_75t_L g820 ( .A(n_680), .B(n_701), .Y(n_820) );
AND2x2_ASAP7_75t_L g732 ( .A(n_681), .B(n_690), .Y(n_732) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g808 ( .A(n_686), .Y(n_808) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_692), .C(n_698), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g730 ( .A(n_690), .Y(n_730) );
AND2x4_ASAP7_75t_SL g766 ( .A(n_690), .B(n_709), .Y(n_766) );
INVx1_ASAP7_75t_SL g777 ( .A(n_690), .Y(n_777) );
OR2x2_ASAP7_75t_L g729 ( .A(n_691), .B(n_730), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_696), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
AND2x4_ASAP7_75t_L g706 ( .A(n_694), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g764 ( .A(n_695), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x4_ASAP7_75t_L g786 ( .A(n_697), .B(n_787), .Y(n_786) );
AND2x2_ASAP7_75t_L g811 ( .A(n_697), .B(n_791), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_703), .B1(n_705), .B2(n_708), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
AND2x4_ASAP7_75t_L g746 ( .A(n_702), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g768 ( .A(n_702), .Y(n_768) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g823 ( .A(n_706), .B(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_719), .C(n_727), .Y(n_710) );
AOI21xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .B(n_717), .Y(n_711) );
INVx1_ASAP7_75t_L g792 ( .A(n_713), .Y(n_792) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AOI222xp33_ASAP7_75t_L g815 ( .A1(n_718), .A2(n_816), .B1(n_819), .B2(n_821), .C1(n_823), .C2(n_825), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_721), .B(n_811), .Y(n_810) );
INVx3_ASAP7_75t_L g744 ( .A(n_722), .Y(n_744) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
O2A1O1Ixp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B(n_731), .C(n_733), .Y(n_727) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NOR2x1_ASAP7_75t_L g735 ( .A(n_736), .B(n_793), .Y(n_735) );
NAND4xp25_ASAP7_75t_L g736 ( .A(n_737), .B(n_759), .C(n_769), .D(n_780), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_748), .B1(n_750), .B2(n_752), .Y(n_737) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_742), .C(n_745), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_739), .B(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g765 ( .A(n_741), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_743), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AND2x4_ASAP7_75t_L g752 ( .A(n_753), .B(n_756), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
BUFx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g790 ( .A(n_755), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g804 ( .A(n_756), .Y(n_804) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_757), .Y(n_822) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx3_ASAP7_75t_L g817 ( .A(n_766), .Y(n_817) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
A2O1A1Ixp33_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B(n_772), .C(n_778), .Y(n_769) );
AOI21xp33_ASAP7_75t_SL g772 ( .A1(n_773), .A2(n_774), .B(n_775), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_773), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_782), .B1(n_783), .B2(n_786), .C(n_788), .Y(n_780) );
INVx1_ASAP7_75t_L g818 ( .A(n_781), .Y(n_818) );
AOI31xp33_ASAP7_75t_L g802 ( .A1(n_784), .A2(n_803), .A3(n_804), .B(n_805), .Y(n_802) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g791 ( .A(n_787), .Y(n_791) );
INVxp67_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NAND3xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_806), .C(n_815), .Y(n_793) );
AOI221xp5_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_797), .B1(n_799), .B2(n_801), .C(n_802), .Y(n_794) );
INVx2_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_SL g803 ( .A(n_801), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_809), .B1(n_812), .B2(n_814), .Y(n_806) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx6_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
AND2x6_ASAP7_75t_SL g830 ( .A(n_831), .B(n_833), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx3_ASAP7_75t_L g841 ( .A(n_832), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_832), .B(n_859), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_832), .B(n_872), .Y(n_879) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
AOI21xp5_ASAP7_75t_SL g839 ( .A1(n_840), .A2(n_842), .B(n_854), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_841), .B(n_870), .Y(n_869) );
INVxp33_ASAP7_75t_L g873 ( .A(n_842), .Y(n_873) );
OAI21xp5_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_848), .B(n_851), .Y(n_842) );
XNOR2x1_ASAP7_75t_L g843 ( .A(n_844), .B(n_847), .Y(n_843) );
INVx4_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
BUFx12f_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NOR2xp67_ASAP7_75t_SL g852 ( .A(n_850), .B(n_853), .Y(n_852) );
INVxp67_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
INVx6_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
BUFx10_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
OAI21xp33_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_873), .B(n_874), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_864), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_865), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_866), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_867), .Y(n_866) );
OR2x6_ASAP7_75t_L g867 ( .A(n_868), .B(n_872), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
OR2x4_ASAP7_75t_L g878 ( .A(n_870), .B(n_879), .Y(n_878) );
BUFx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx4_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
BUFx3_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
endmodule