module real_aes_8352_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
OAI22xp5_ASAP7_75t_SL g186 ( .A1(n_0), .A2(n_50), .B1(n_187), .B2(n_188), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_0), .Y(n_188) );
INVx1_ASAP7_75t_L g230 ( .A(n_1), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_2), .Y(n_172) );
AOI21xp33_ASAP7_75t_L g274 ( .A1(n_3), .A2(n_246), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g203 ( .A(n_4), .Y(n_203) );
AND2x6_ASAP7_75t_L g224 ( .A(n_4), .B(n_201), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_4), .B(n_530), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_5), .A2(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g280 ( .A(n_6), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_7), .B(n_309), .Y(n_308) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_8), .A2(n_26), .B1(n_90), .B2(n_91), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_9), .Y(n_167) );
INVx1_ASAP7_75t_L g216 ( .A(n_10), .Y(n_216) );
INVx1_ASAP7_75t_L g334 ( .A(n_11), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g114 ( .A1(n_12), .A2(n_20), .B1(n_115), .B2(n_122), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_13), .B(n_251), .Y(n_322) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_14), .A2(n_27), .B1(n_90), .B2(n_94), .Y(n_93) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_15), .A2(n_183), .B1(n_189), .B2(n_190), .Y(n_182) );
INVx1_ASAP7_75t_L g189 ( .A(n_15), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_15), .B(n_246), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_16), .B(n_258), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_17), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_18), .A2(n_332), .B(n_333), .C(n_335), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_19), .Y(n_130) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_21), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_22), .B(n_234), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_23), .Y(n_138) );
INVx1_ASAP7_75t_L g269 ( .A(n_24), .Y(n_269) );
INVx2_ASAP7_75t_L g222 ( .A(n_25), .Y(n_222) );
OAI221xp5_ASAP7_75t_L g194 ( .A1(n_27), .A2(n_40), .B1(n_47), .B2(n_195), .C(n_196), .Y(n_194) );
INVxp67_ASAP7_75t_L g197 ( .A(n_27), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g292 ( .A1(n_28), .A2(n_224), .B(n_226), .C(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g267 ( .A(n_29), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_30), .A2(n_80), .B1(n_180), .B2(n_181), .Y(n_79) );
INVx1_ASAP7_75t_L g180 ( .A(n_30), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_31), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_32), .B(n_234), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_33), .A2(n_54), .B1(n_142), .B2(n_146), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g270 ( .A(n_34), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_35), .B(n_246), .Y(n_311) );
AOI22xp5_ASAP7_75t_SL g525 ( .A1(n_35), .A2(n_80), .B1(n_181), .B2(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_35), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_36), .A2(n_226), .B1(n_236), .B2(n_265), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_37), .A2(n_76), .B1(n_151), .B2(n_156), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_38), .Y(n_301) );
CKINVDCx16_ASAP7_75t_R g218 ( .A(n_39), .Y(n_218) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_40), .A2(n_58), .B1(n_90), .B2(n_94), .Y(n_99) );
INVxp67_ASAP7_75t_L g198 ( .A(n_40), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_41), .A2(n_254), .B(n_278), .C(n_279), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_42), .Y(n_325) );
INVx1_ASAP7_75t_L g276 ( .A(n_43), .Y(n_276) );
INVx1_ASAP7_75t_L g201 ( .A(n_44), .Y(n_201) );
INVx1_ASAP7_75t_L g215 ( .A(n_45), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_46), .Y(n_195) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_47), .A2(n_64), .B1(n_90), .B2(n_91), .Y(n_97) );
A2O1A1Ixp33_ASAP7_75t_SL g250 ( .A1(n_48), .A2(n_251), .B(n_252), .C(n_254), .Y(n_250) );
INVxp67_ASAP7_75t_L g253 ( .A(n_49), .Y(n_253) );
CKINVDCx16_ASAP7_75t_R g187 ( .A(n_50), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_51), .A2(n_80), .B1(n_181), .B2(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_51), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_52), .Y(n_272) );
INVx1_ASAP7_75t_L g318 ( .A(n_53), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_55), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g319 ( .A1(n_56), .A2(n_224), .B(n_226), .C(n_320), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_57), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_59), .B(n_231), .Y(n_294) );
INVx2_ASAP7_75t_L g213 ( .A(n_60), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_61), .A2(n_184), .B1(n_185), .B2(n_186), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_61), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_62), .B(n_251), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_63), .A2(n_224), .B(n_226), .C(n_229), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_65), .B(n_241), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_66), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_67), .A2(n_224), .B(n_226), .C(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g534 ( .A(n_67), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_68), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_69), .Y(n_162) );
INVx1_ASAP7_75t_L g249 ( .A(n_70), .Y(n_249) );
CKINVDCx16_ASAP7_75t_R g330 ( .A(n_71), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_72), .B(n_231), .Y(n_307) );
INVx1_ASAP7_75t_L g90 ( .A(n_73), .Y(n_90) );
INVx1_ASAP7_75t_L g92 ( .A(n_73), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_74), .B(n_244), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_75), .A2(n_246), .B(n_247), .Y(n_245) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_191), .B1(n_204), .B2(n_520), .C(n_524), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_182), .Y(n_78) );
INVx2_ASAP7_75t_L g181 ( .A(n_80), .Y(n_181) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_139), .Y(n_80) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_106), .C(n_127), .Y(n_81) );
OAI22xp5_ASAP7_75t_SL g82 ( .A1(n_83), .A2(n_100), .B1(n_101), .B2(n_105), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
OR2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
INVx2_ASAP7_75t_L g149 ( .A(n_87), .Y(n_149) );
OR2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
AND2x2_ASAP7_75t_L g104 ( .A(n_88), .B(n_93), .Y(n_104) );
AND2x2_ASAP7_75t_L g145 ( .A(n_88), .B(n_120), .Y(n_145) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g110 ( .A(n_89), .B(n_93), .Y(n_110) );
AND2x2_ASAP7_75t_L g121 ( .A(n_89), .B(n_99), .Y(n_121) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g94 ( .A(n_92), .Y(n_94) );
INVx2_ASAP7_75t_L g120 ( .A(n_93), .Y(n_120) );
INVx1_ASAP7_75t_L g159 ( .A(n_93), .Y(n_159) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
NAND2x1p5_ASAP7_75t_L g103 ( .A(n_96), .B(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g175 ( .A(n_96), .B(n_145), .Y(n_175) );
AND2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_98), .Y(n_96) );
INVx1_ASAP7_75t_L g112 ( .A(n_97), .Y(n_112) );
INVx1_ASAP7_75t_L g119 ( .A(n_97), .Y(n_119) );
INVx1_ASAP7_75t_L g137 ( .A(n_97), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_97), .B(n_99), .Y(n_160) );
AND2x2_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g155 ( .A(n_99), .B(n_137), .Y(n_155) );
BUFx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g154 ( .A(n_104), .B(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g166 ( .A(n_104), .B(n_111), .Y(n_166) );
OAI21xp33_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_113), .B(n_114), .Y(n_106) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x6_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
AND2x2_ASAP7_75t_L g144 ( .A(n_111), .B(n_145), .Y(n_144) );
AND2x6_ASAP7_75t_L g148 ( .A(n_111), .B(n_149), .Y(n_148) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVx1_ASAP7_75t_L g126 ( .A(n_119), .Y(n_126) );
INVx1_ASAP7_75t_L g129 ( .A(n_120), .Y(n_129) );
AND2x4_ASAP7_75t_L g125 ( .A(n_121), .B(n_126), .Y(n_125) );
NAND2x1p5_ASAP7_75t_L g128 ( .A(n_121), .B(n_129), .Y(n_128) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx12f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp33_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_130), .B1(n_131), .B2(n_138), .Y(n_127) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g132 ( .A(n_133), .Y(n_132) );
OR2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR3xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_161), .C(n_171), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_150), .Y(n_140) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_145), .B(n_155), .Y(n_170) );
AND2x4_ASAP7_75t_L g178 ( .A(n_145), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx11_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx8_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx6_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
OR2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx1_ASAP7_75t_L g179 ( .A(n_160), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B1(n_167), .B2(n_168), .Y(n_161) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx6_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B1(n_176), .B2(n_177), .Y(n_171) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_183), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_193), .Y(n_192) );
AND3x1_ASAP7_75t_SL g193 ( .A(n_194), .B(n_199), .C(n_202), .Y(n_193) );
INVxp67_ASAP7_75t_L g530 ( .A(n_194), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_199), .A2(n_226), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g540 ( .A(n_199), .Y(n_540) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OAI322xp33_ASAP7_75t_L g524 ( .A1(n_200), .A2(n_525), .A3(n_527), .B1(n_531), .B2(n_534), .C1(n_535), .C2(n_537), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_200), .B(n_203), .Y(n_533) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_SL g539 ( .A(n_202), .B(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_203), .Y(n_202) );
OR4x1_ASAP7_75t_L g204 ( .A(n_205), .B(n_409), .C(n_469), .D(n_496), .Y(n_204) );
NAND4xp25_ASAP7_75t_SL g205 ( .A(n_206), .B(n_357), .C(n_388), .D(n_405), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_282), .B(n_284), .C(n_337), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_260), .Y(n_207) );
INVx1_ASAP7_75t_L g399 ( .A(n_208), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_208), .A2(n_440), .B1(n_488), .B2(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_242), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_209), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g350 ( .A(n_209), .B(n_262), .Y(n_350) );
AND2x2_ASAP7_75t_L g392 ( .A(n_209), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_209), .B(n_283), .Y(n_404) );
INVx1_ASAP7_75t_L g444 ( .A(n_209), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_209), .B(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g372 ( .A(n_210), .B(n_262), .Y(n_372) );
INVx3_ASAP7_75t_L g376 ( .A(n_210), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_210), .B(n_434), .Y(n_433) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_217), .B(n_238), .Y(n_210) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_211), .A2(n_263), .B(n_271), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_211), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g299 ( .A(n_211), .Y(n_299) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_212), .Y(n_244) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AND2x2_ASAP7_75t_SL g241 ( .A(n_213), .B(n_214), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_225), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g263 ( .A1(n_219), .A2(n_256), .B1(n_264), .B2(n_270), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_219), .A2(n_318), .B(n_319), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g219 ( .A(n_220), .B(n_224), .Y(n_219) );
AND2x4_ASAP7_75t_L g246 ( .A(n_220), .B(n_224), .Y(n_246) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_223), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g227 ( .A(n_222), .Y(n_227) );
INVx1_ASAP7_75t_L g237 ( .A(n_222), .Y(n_237) );
INVx1_ASAP7_75t_L g228 ( .A(n_223), .Y(n_228) );
INVx3_ASAP7_75t_L g232 ( .A(n_223), .Y(n_232) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_223), .Y(n_234) );
INVx1_ASAP7_75t_L g251 ( .A(n_223), .Y(n_251) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_223), .Y(n_266) );
INVx4_ASAP7_75t_SL g256 ( .A(n_224), .Y(n_256) );
BUFx3_ASAP7_75t_L g523 ( .A(n_224), .Y(n_523) );
INVx5_ASAP7_75t_L g248 ( .A(n_226), .Y(n_248) );
AND2x2_ASAP7_75t_L g522 ( .A(n_226), .B(n_523), .Y(n_522) );
AND2x6_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_227), .Y(n_255) );
BUFx3_ASAP7_75t_L g298 ( .A(n_227), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_233), .C(n_235), .Y(n_229) );
INVx5_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_232), .B(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_232), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g278 ( .A(n_234), .Y(n_278) );
INVx4_ASAP7_75t_L g309 ( .A(n_234), .Y(n_309) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_240), .B(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_240), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g303 ( .A(n_241), .Y(n_303) );
OA21x2_ASAP7_75t_L g326 ( .A1(n_241), .A2(n_327), .B(n_336), .Y(n_326) );
AND2x2_ASAP7_75t_L g463 ( .A(n_242), .B(n_273), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_242), .B(n_376), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_242), .B(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g283 ( .A(n_243), .B(n_262), .Y(n_283) );
INVx1_ASAP7_75t_L g345 ( .A(n_243), .Y(n_345) );
BUFx2_ASAP7_75t_L g349 ( .A(n_243), .Y(n_349) );
AND2x2_ASAP7_75t_L g393 ( .A(n_243), .B(n_261), .Y(n_393) );
OR2x2_ASAP7_75t_L g432 ( .A(n_243), .B(n_261), .Y(n_432) );
AND2x2_ASAP7_75t_L g457 ( .A(n_243), .B(n_273), .Y(n_457) );
AND2x2_ASAP7_75t_L g516 ( .A(n_243), .B(n_346), .Y(n_516) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_257), .Y(n_243) );
INVx4_ASAP7_75t_L g259 ( .A(n_244), .Y(n_259) );
BUFx2_ASAP7_75t_L g328 ( .A(n_246), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_250), .C(n_256), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g275 ( .A1(n_248), .A2(n_256), .B(n_276), .C(n_277), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_248), .A2(n_256), .B(n_330), .C(n_331), .Y(n_329) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_255), .Y(n_310) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_258), .A2(n_274), .B(n_281), .Y(n_273) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_SL g300 ( .A(n_259), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g491 ( .A(n_260), .Y(n_491) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_273), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_261), .B(n_273), .Y(n_377) );
AND2x2_ASAP7_75t_L g387 ( .A(n_261), .B(n_376), .Y(n_387) );
BUFx2_ASAP7_75t_L g398 ( .A(n_261), .Y(n_398) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g420 ( .A(n_262), .B(n_273), .Y(n_420) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_262), .Y(n_475) );
OAI22xp5_ASAP7_75t_SL g265 ( .A1(n_266), .A2(n_267), .B1(n_268), .B2(n_269), .Y(n_265) );
INVx2_ASAP7_75t_L g268 ( .A(n_266), .Y(n_268) );
INVx4_ASAP7_75t_L g332 ( .A(n_266), .Y(n_332) );
AND2x2_ASAP7_75t_SL g282 ( .A(n_273), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g346 ( .A(n_273), .Y(n_346) );
BUFx2_ASAP7_75t_L g371 ( .A(n_273), .Y(n_371) );
INVx2_ASAP7_75t_L g390 ( .A(n_273), .Y(n_390) );
AND2x2_ASAP7_75t_L g452 ( .A(n_273), .B(n_376), .Y(n_452) );
AOI321xp33_ASAP7_75t_L g471 ( .A1(n_282), .A2(n_472), .A3(n_473), .B1(n_474), .B2(n_476), .C(n_477), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_283), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_283), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g465 ( .A(n_283), .B(n_444), .Y(n_465) );
AND2x2_ASAP7_75t_L g498 ( .A(n_283), .B(n_390), .Y(n_498) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_314), .Y(n_285) );
OR2x2_ASAP7_75t_L g400 ( .A(n_286), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_302), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g352 ( .A(n_289), .Y(n_352) );
AND2x2_ASAP7_75t_L g362 ( .A(n_289), .B(n_316), .Y(n_362) );
AND2x2_ASAP7_75t_L g367 ( .A(n_289), .B(n_342), .Y(n_367) );
INVx1_ASAP7_75t_L g384 ( .A(n_289), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_289), .B(n_365), .Y(n_403) );
AND2x2_ASAP7_75t_L g408 ( .A(n_289), .B(n_341), .Y(n_408) );
OR2x2_ASAP7_75t_L g440 ( .A(n_289), .B(n_429), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_289), .B(n_353), .Y(n_479) );
AND2x2_ASAP7_75t_L g513 ( .A(n_289), .B(n_339), .Y(n_513) );
OR2x6_ASAP7_75t_L g289 ( .A(n_290), .B(n_300), .Y(n_289) );
AOI21xp5_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_292), .B(n_299), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B(n_296), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_296), .A2(n_321), .B(n_322), .Y(n_320) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g335 ( .A(n_298), .Y(n_335) );
INVx1_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
INVx1_ASAP7_75t_L g340 ( .A(n_302), .Y(n_340) );
INVx2_ASAP7_75t_L g355 ( .A(n_302), .Y(n_355) );
AND2x2_ASAP7_75t_L g395 ( .A(n_302), .B(n_366), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_302), .B(n_342), .Y(n_417) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_312), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_311), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B(n_310), .Y(n_306) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g501 ( .A(n_315), .B(n_352), .Y(n_501) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_326), .Y(n_315) );
INVx2_ASAP7_75t_L g342 ( .A(n_316), .Y(n_342) );
AND2x2_ASAP7_75t_L g495 ( .A(n_316), .B(n_355), .Y(n_495) );
AO21x2_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_323), .B(n_324), .Y(n_316) );
AND2x2_ASAP7_75t_L g341 ( .A(n_326), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g356 ( .A(n_326), .Y(n_356) );
INVx1_ASAP7_75t_L g366 ( .A(n_326), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_332), .B(n_334), .Y(n_333) );
OAI22xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_343), .B1(n_347), .B2(n_351), .Y(n_337) );
OAI22xp33_ASAP7_75t_L g492 ( .A1(n_338), .A2(n_456), .B1(n_493), .B2(n_494), .Y(n_492) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g407 ( .A(n_340), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_341), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g402 ( .A(n_342), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_342), .B(n_355), .Y(n_429) );
INVx1_ASAP7_75t_L g445 ( .A(n_342), .Y(n_445) );
AND2x2_ASAP7_75t_L g386 ( .A(n_344), .B(n_387), .Y(n_386) );
INVx3_ASAP7_75t_SL g425 ( .A(n_344), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_344), .B(n_350), .Y(n_502) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g511 ( .A(n_347), .Y(n_511) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_348), .B(n_444), .Y(n_486) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx3_ASAP7_75t_SL g391 ( .A(n_350), .Y(n_391) );
NAND2x1_ASAP7_75t_SL g351 ( .A(n_352), .B(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_L g412 ( .A(n_352), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g419 ( .A(n_352), .B(n_356), .Y(n_419) );
AND2x2_ASAP7_75t_L g424 ( .A(n_352), .B(n_365), .Y(n_424) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_352), .Y(n_473) );
OAI311xp33_ASAP7_75t_L g496 ( .A1(n_353), .A2(n_497), .A3(n_499), .B1(n_500), .C1(n_510), .Y(n_496) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g509 ( .A(n_354), .B(n_382), .Y(n_509) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
AND2x2_ASAP7_75t_L g365 ( .A(n_355), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g413 ( .A(n_355), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g468 ( .A(n_355), .Y(n_468) );
INVx1_ASAP7_75t_L g361 ( .A(n_356), .Y(n_361) );
INVx1_ASAP7_75t_L g381 ( .A(n_356), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_356), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g414 ( .A(n_356), .Y(n_414) );
AOI221xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_360), .B1(n_368), .B2(n_373), .C(n_378), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_363), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx4_ASAP7_75t_L g382 ( .A(n_362), .Y(n_382) );
AND2x2_ASAP7_75t_L g476 ( .A(n_362), .B(n_395), .Y(n_476) );
AND2x2_ASAP7_75t_L g483 ( .A(n_362), .B(n_365), .Y(n_483) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_365), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g394 ( .A(n_367), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_370), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g519 ( .A(n_372), .B(n_463), .Y(n_519) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g504 ( .A(n_376), .B(n_432), .Y(n_504) );
OAI211xp5_ASAP7_75t_L g469 ( .A1(n_377), .A2(n_470), .B(n_471), .C(n_484), .Y(n_469) );
AOI21xp33_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_383), .B(n_385), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp67_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g448 ( .A(n_382), .Y(n_448) );
OAI221xp5_ASAP7_75t_L g477 ( .A1(n_383), .A2(n_478), .B1(n_479), .B2(n_480), .C(n_481), .Y(n_477) );
AND2x2_ASAP7_75t_L g454 ( .A(n_384), .B(n_395), .Y(n_454) );
AND2x2_ASAP7_75t_L g507 ( .A(n_384), .B(n_402), .Y(n_507) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_387), .B(n_425), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_392), .B(n_394), .C(n_396), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AND2x2_ASAP7_75t_L g435 ( .A(n_390), .B(n_393), .Y(n_435) );
OR2x2_ASAP7_75t_L g478 ( .A(n_390), .B(n_432), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_391), .B(n_457), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_391), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g422 ( .A(n_392), .Y(n_422) );
INVx1_ASAP7_75t_L g488 ( .A(n_395), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .B1(n_403), .B2(n_404), .Y(n_396) );
INVx1_ASAP7_75t_L g411 ( .A(n_397), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_398), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g474 ( .A(n_399), .B(n_475), .Y(n_474) );
INVxp67_ASAP7_75t_L g460 ( .A(n_401), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_402), .B(n_488), .Y(n_487) );
OAI22xp33_ASAP7_75t_L g461 ( .A1(n_403), .A2(n_462), .B1(n_464), .B2(n_466), .Y(n_461) );
INVx1_ASAP7_75t_L g470 ( .A(n_406), .Y(n_470) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
AND2x2_ASAP7_75t_L g512 ( .A(n_407), .B(n_507), .Y(n_512) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_408), .A2(n_442), .B1(n_445), .B2(n_446), .C1(n_449), .C2(n_450), .Y(n_441) );
NAND4xp25_ASAP7_75t_SL g409 ( .A(n_410), .B(n_430), .C(n_441), .D(n_453), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B1(n_415), .B2(n_420), .C(n_421), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_413), .B(n_448), .Y(n_447) );
INVxp67_ASAP7_75t_L g439 ( .A(n_414), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_415), .A2(n_485), .B1(n_487), .B2(n_489), .C(n_492), .Y(n_484) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g427 ( .A(n_419), .B(n_428), .Y(n_427) );
OAI21xp33_ASAP7_75t_L g481 ( .A1(n_420), .A2(n_482), .B(n_483), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_425), .B2(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI21xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B(n_436), .Y(n_430) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g472 ( .A(n_443), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_444), .B(n_463), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_444), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_448), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g480 ( .A(n_452), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B1(n_458), .B2(n_460), .C(n_461), .Y(n_453) );
INVxp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AOI222xp33_ASAP7_75t_L g500 ( .A1(n_463), .A2(n_501), .B1(n_502), .B2(n_503), .C1(n_505), .C2(n_508), .Y(n_500) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_467), .B(n_507), .Y(n_506) );
INVxp67_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g499 ( .A(n_473), .Y(n_499) );
INVxp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVxp33_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_513), .B2(n_514), .C(n_517), .Y(n_510) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVxp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_529), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
endmodule