module fake_jpeg_17971_n_84 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_84);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_84;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx8_ASAP7_75t_SL g10 ( 
.A(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx4f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_13),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_29),
.B1(n_20),
.B2(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_4),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_13),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_36),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_21),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_39),
.B(n_14),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_20),
.B1(n_15),
.B2(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_19),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_17),
.B1(n_19),
.B2(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_29),
.C(n_26),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_52),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_10),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_53),
.A2(n_54),
.B(n_34),
.Y(n_55)
);

AND2x4_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_27),
.Y(n_54)
);

AO22x1_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_54),
.B1(n_53),
.B2(n_50),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_62),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_54),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_68),
.Y(n_69)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_52),
.Y(n_68)
);

OAI322xp33_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_55),
.A3(n_61),
.B1(n_43),
.B2(n_33),
.C1(n_56),
.C2(n_59),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

AOI321xp33_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_71),
.A3(n_64),
.B1(n_73),
.B2(n_33),
.C(n_14),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_71),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_78),
.Y(n_81)
);

NOR2xp67_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_74),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_81),
.Y(n_83)
);

AOI221xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_7),
.B1(n_9),
.B2(n_44),
.C(n_57),
.Y(n_84)
);


endmodule