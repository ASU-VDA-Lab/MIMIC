module fake_jpeg_3747_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_6),
.B(n_0),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_15),
.B(n_18),
.Y(n_29)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVxp67_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_7),
.B(n_5),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_11),
.A2(n_2),
.B1(n_3),
.B2(n_10),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_19),
.A2(n_20),
.B1(n_13),
.B2(n_14),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_11),
.A2(n_2),
.B1(n_12),
.B2(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_8),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_14),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_12),
.A2(n_13),
.B(n_14),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_15),
.B(n_16),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_31),
.B(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_18),
.C(n_17),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_39),
.B(n_26),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_42),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_26),
.B(n_29),
.Y(n_43)
);

AOI322xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_24),
.A3(n_32),
.B1(n_34),
.B2(n_38),
.C1(n_39),
.C2(n_41),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_44),
.Y(n_47)
);


endmodule