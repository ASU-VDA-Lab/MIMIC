module fake_ariane_234_n_1848 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1848);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1848;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1603;
wire n_1370;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_36),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_61),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_130),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_2),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_42),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_95),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_116),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_78),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_29),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_174),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_49),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_34),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_93),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_176),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_59),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_109),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_77),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_84),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_72),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_73),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_61),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_7),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_115),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_28),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_27),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_53),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_79),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_128),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_119),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_178),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_90),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_173),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_24),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_38),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_53),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_9),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_143),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_16),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_131),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_87),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_24),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_14),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_76),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_144),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_100),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_2),
.Y(n_233)
);

INVx4_ASAP7_75t_R g234 ( 
.A(n_17),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_26),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_44),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_32),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_65),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_81),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_31),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_37),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_133),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_145),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_89),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_179),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_88),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_169),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_12),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_170),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_122),
.Y(n_250)
);

BUFx8_ASAP7_75t_SL g251 ( 
.A(n_161),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_107),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_49),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_12),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_18),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_28),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_38),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_62),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_135),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_41),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_5),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_30),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_82),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_151),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_42),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_83),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_44),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_0),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_152),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_99),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_71),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_129),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_180),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_134),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_41),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_137),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_62),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_157),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_64),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_58),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_111),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_13),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_146),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_171),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_69),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_16),
.Y(n_286)
);

BUFx8_ASAP7_75t_SL g287 ( 
.A(n_21),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_155),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_108),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_33),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_181),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_9),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_29),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_125),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_57),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_8),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_40),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_50),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_4),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_15),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_85),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_167),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_66),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_114),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_75),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_63),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_20),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_64),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_91),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_43),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_43),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_36),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_20),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_58),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_80),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_0),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_165),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_5),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_150),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_45),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_159),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_94),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_126),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_57),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_14),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_3),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_3),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_31),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_56),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_96),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_59),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_148),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_11),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_17),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_177),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_175),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_113),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_22),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_60),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_13),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_30),
.Y(n_341)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_1),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_98),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_45),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_92),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_52),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_74),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_156),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_106),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_67),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_48),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_104),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_86),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_34),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_37),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_118),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_8),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_55),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_154),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_39),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_121),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_138),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_15),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_50),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_287),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_1),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_262),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_325),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_287),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_262),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_262),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_215),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_262),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_251),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_257),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_262),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_262),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_251),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_262),
.Y(n_379)
);

INVxp33_ASAP7_75t_SL g380 ( 
.A(n_282),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_231),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_191),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_182),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_189),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_258),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_191),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_190),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_284),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_209),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_342),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_342),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_218),
.B(n_4),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_192),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_258),
.Y(n_396)
);

INVxp33_ASAP7_75t_SL g397 ( 
.A(n_194),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_342),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_235),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_342),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_237),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_192),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_342),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_245),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_241),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_258),
.Y(n_408)
);

INVxp33_ASAP7_75t_SL g409 ( 
.A(n_194),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_219),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_196),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_185),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_219),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_248),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_274),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_256),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_261),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_219),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_219),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_254),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_229),
.B(n_6),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_265),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_245),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_222),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_270),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_278),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_222),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_275),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_286),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_222),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_184),
.B(n_6),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_222),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_227),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_227),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_227),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_227),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_240),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_292),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_240),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_296),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_260),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_260),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_267),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_267),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_254),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_280),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_312),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_297),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_280),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_278),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_210),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_298),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_210),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_323),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_228),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_228),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_284),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_323),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_374),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_385),
.B(n_187),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_367),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_396),
.B(n_198),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_420),
.B(n_205),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_382),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_365),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_386),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_367),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_370),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_378),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_395),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_370),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_371),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_369),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_212),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_403),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_405),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_397),
.B(n_201),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_383),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_423),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_373),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_426),
.Y(n_481)
);

INVxp33_ASAP7_75t_SL g482 ( 
.A(n_384),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_371),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_373),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_376),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_387),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_376),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_450),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_389),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_377),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_377),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_379),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_390),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_411),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_L g496 ( 
.A(n_366),
.B(n_299),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_399),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_401),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_406),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_390),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_414),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_392),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_392),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_451),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_393),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_393),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_398),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_398),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_400),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_372),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_402),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_402),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_404),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_404),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_453),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_416),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_454),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_417),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_422),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

OA21x2_ASAP7_75t_L g522 ( 
.A1(n_431),
.A2(n_223),
.B(n_214),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_454),
.Y(n_523)
);

BUFx8_ASAP7_75t_L g524 ( 
.A(n_366),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_388),
.B(n_225),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_388),
.B(n_232),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_457),
.B(n_337),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_429),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_458),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_455),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_456),
.A2(n_255),
.B1(n_354),
.B2(n_277),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_458),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_408),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_457),
.B(n_238),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_R g535 ( 
.A(n_438),
.B(n_196),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_425),
.B(n_372),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_522),
.A2(n_394),
.B1(n_421),
.B2(n_368),
.Y(n_537)
);

AND2x6_ASAP7_75t_L g538 ( 
.A(n_461),
.B(n_337),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_533),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_487),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_533),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_518),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_513),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_461),
.B(n_319),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_463),
.B(n_447),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_513),
.B(n_381),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_513),
.B(n_515),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_522),
.A2(n_380),
.B1(n_211),
.B2(n_224),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_519),
.B(n_425),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_461),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_489),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_477),
.B(n_409),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_467),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_519),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_474),
.B(n_447),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_522),
.A2(n_220),
.B1(n_236),
.B2(n_233),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_487),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_468),
.B(n_415),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_513),
.B(n_440),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_521),
.B(n_412),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_483),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_497),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_515),
.B(n_448),
.Y(n_563)
);

BUFx8_ASAP7_75t_SL g564 ( 
.A(n_504),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_484),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_521),
.B(n_452),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_523),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_515),
.B(n_468),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_527),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_515),
.B(n_239),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_511),
.B(n_375),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_471),
.B(n_480),
.Y(n_572)
);

NOR3xp33_ASAP7_75t_L g573 ( 
.A(n_495),
.B(n_221),
.C(n_279),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_529),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g575 ( 
.A(n_536),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_482),
.A2(n_200),
.B1(n_206),
.B2(n_197),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_471),
.B(n_447),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_480),
.B(n_244),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_498),
.B(n_391),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_483),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_487),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_484),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_460),
.B(n_408),
.Y(n_583)
);

AO22x2_ASAP7_75t_L g584 ( 
.A1(n_524),
.A2(n_407),
.B1(n_201),
.B2(n_289),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_529),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_532),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_467),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_524),
.A2(n_289),
.B1(n_268),
.B2(n_364),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_499),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_532),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_522),
.A2(n_341),
.B1(n_307),
.B2(n_308),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_490),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_516),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_484),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_501),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_490),
.Y(n_596)
);

OR2x6_ASAP7_75t_L g597 ( 
.A(n_459),
.B(n_437),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_467),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_491),
.B(n_410),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_491),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_527),
.A2(n_363),
.B1(n_333),
.B2(n_290),
.Y(n_601)
);

AND2x6_ASAP7_75t_L g602 ( 
.A(n_472),
.B(n_319),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_517),
.B(n_197),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_494),
.B(n_250),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_472),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_528),
.B(n_255),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_494),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_500),
.B(n_252),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_472),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_485),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_469),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_500),
.B(n_264),
.Y(n_612)
);

NAND2x1p5_ASAP7_75t_L g613 ( 
.A(n_459),
.B(n_186),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_478),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_486),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_520),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_462),
.B(n_437),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_475),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_479),
.B(n_200),
.Y(n_619)
);

INVx6_ASAP7_75t_L g620 ( 
.A(n_487),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_503),
.B(n_272),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_481),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_485),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_485),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_503),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_505),
.B(n_283),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_493),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_493),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_530),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_487),
.Y(n_630)
);

INVx6_ASAP7_75t_L g631 ( 
.A(n_487),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_493),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_483),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_465),
.B(n_439),
.Y(n_634)
);

BUFx10_ASAP7_75t_L g635 ( 
.A(n_473),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_492),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_505),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_502),
.Y(n_638)
);

INVx4_ASAP7_75t_SL g639 ( 
.A(n_527),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_508),
.B(n_410),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_525),
.B(n_206),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_502),
.B(n_506),
.Y(n_642)
);

BUFx4f_ASAP7_75t_L g643 ( 
.A(n_527),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_535),
.A2(n_354),
.B1(n_277),
.B2(n_314),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_508),
.B(n_439),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_526),
.B(n_441),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_502),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_L g648 ( 
.A(n_492),
.B(n_263),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_464),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_466),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_506),
.Y(n_651)
);

OR2x6_ASAP7_75t_L g652 ( 
.A(n_531),
.B(n_441),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_492),
.Y(n_653)
);

NOR3xp33_ASAP7_75t_L g654 ( 
.A(n_496),
.B(n_355),
.C(n_300),
.Y(n_654)
);

OR2x6_ASAP7_75t_L g655 ( 
.A(n_531),
.B(n_442),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_509),
.B(n_510),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_509),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_534),
.B(n_355),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_527),
.A2(n_331),
.B1(n_324),
.B2(n_295),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_527),
.B(n_312),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_506),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_510),
.B(n_514),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_507),
.Y(n_663)
);

INVxp33_ASAP7_75t_L g664 ( 
.A(n_470),
.Y(n_664)
);

OR2x6_ASAP7_75t_L g665 ( 
.A(n_524),
.B(n_442),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_476),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_483),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_514),
.B(n_413),
.Y(n_668)
);

AND3x2_ASAP7_75t_L g669 ( 
.A(n_524),
.B(n_234),
.C(n_443),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_492),
.B(n_285),
.Y(n_670)
);

AND2x6_ASAP7_75t_L g671 ( 
.A(n_507),
.B(n_362),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_507),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_488),
.B(n_443),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_492),
.Y(n_674)
);

OAI22xp33_ASAP7_75t_L g675 ( 
.A1(n_483),
.A2(n_314),
.B1(n_306),
.B2(n_310),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_492),
.Y(n_676)
);

AND2x6_ASAP7_75t_L g677 ( 
.A(n_512),
.B(n_362),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_512),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_512),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_512),
.B(n_413),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_512),
.B(n_288),
.Y(n_681)
);

INVx5_ASAP7_75t_L g682 ( 
.A(n_527),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_527),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_461),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_592),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_579),
.B(n_195),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_561),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_649),
.Y(n_688)
);

BUFx5_ASAP7_75t_L g689 ( 
.A(n_642),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_552),
.B(n_311),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_550),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_548),
.A2(n_309),
.B1(n_301),
.B2(n_273),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_552),
.B(n_313),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_583),
.B(n_294),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_546),
.B(n_318),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_546),
.B(n_320),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_558),
.B(n_326),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_596),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_583),
.B(n_322),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_600),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_559),
.B(n_327),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_537),
.A2(n_548),
.B1(n_543),
.B2(n_607),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_625),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_550),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_556),
.A2(n_309),
.B1(n_301),
.B2(n_273),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_545),
.B(n_555),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_549),
.B(n_185),
.Y(n_707)
);

INVx8_ASAP7_75t_L g708 ( 
.A(n_665),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_572),
.A2(n_315),
.B(n_304),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_553),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_637),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_545),
.B(n_336),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_537),
.A2(n_563),
.B1(n_559),
.B2(n_555),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_566),
.B(n_540),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_593),
.Y(n_715)
);

BUFx12f_ASAP7_75t_L g716 ( 
.A(n_551),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_545),
.B(n_343),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_553),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_665),
.B(n_618),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_555),
.B(n_199),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_563),
.A2(n_204),
.B1(n_203),
.B2(n_202),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_641),
.B(n_328),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_657),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_551),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_540),
.B(n_199),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_571),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_540),
.B(n_202),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_617),
.B(n_203),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_617),
.B(n_204),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_646),
.B(n_353),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_665),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_658),
.B(n_329),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_669),
.B(n_597),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_587),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_673),
.B(n_649),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_547),
.B(n_334),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_587),
.Y(n_737)
);

NAND2x1p5_ASAP7_75t_L g738 ( 
.A(n_643),
.B(n_317),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_SL g739 ( 
.A(n_611),
.B(n_562),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_554),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_598),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_581),
.B(n_353),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_560),
.B(n_185),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_539),
.B(n_338),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_541),
.B(n_339),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_597),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_542),
.B(n_340),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_567),
.B(n_344),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_581),
.B(n_335),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_547),
.B(n_574),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_654),
.A2(n_347),
.B1(n_352),
.B2(n_359),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_585),
.B(n_346),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_586),
.B(n_357),
.Y(n_753)
);

NAND2x1_ASAP7_75t_L g754 ( 
.A(n_642),
.B(n_183),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_634),
.A2(n_361),
.B1(n_188),
.B2(n_193),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_590),
.B(n_360),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_568),
.B(n_675),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_645),
.B(n_316),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_597),
.B(n_207),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_568),
.A2(n_418),
.B(n_419),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_603),
.B(n_207),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_599),
.Y(n_762)
);

CKINVDCx11_ASAP7_75t_R g763 ( 
.A(n_551),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_640),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_668),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_565),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_598),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_656),
.A2(n_316),
.B1(n_208),
.B2(n_213),
.Y(n_768)
);

NAND3xp33_ASAP7_75t_L g769 ( 
.A(n_576),
.B(n_305),
.C(n_217),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_642),
.B(n_611),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_556),
.A2(n_309),
.B1(n_301),
.B2(n_273),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_645),
.A2(n_433),
.B(n_419),
.C(n_424),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_581),
.B(n_263),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_662),
.A2(n_330),
.B(n_216),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_582),
.B(n_226),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_594),
.B(n_230),
.Y(n_776)
);

AND2x6_ASAP7_75t_SL g777 ( 
.A(n_652),
.B(n_444),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_636),
.B(n_263),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_636),
.B(n_653),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_627),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_636),
.B(n_263),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_561),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_653),
.B(n_263),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_614),
.B(n_207),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_584),
.A2(n_321),
.B1(n_249),
.B2(n_259),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_627),
.B(n_242),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_605),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_647),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_647),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_591),
.B(n_243),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_653),
.B(n_678),
.Y(n_791)
);

NOR2xp67_ASAP7_75t_L g792 ( 
.A(n_615),
.B(n_444),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_616),
.B(n_449),
.C(n_446),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_561),
.B(n_263),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_591),
.B(n_246),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_561),
.B(n_263),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_605),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_629),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_578),
.B(n_247),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_578),
.B(n_266),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_580),
.B(n_269),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_589),
.B(n_253),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_595),
.B(n_253),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_609),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_613),
.B(n_253),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_613),
.B(n_635),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_L g807 ( 
.A(n_642),
.B(n_269),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_609),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_604),
.B(n_271),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_619),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_604),
.B(n_276),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_L g812 ( 
.A(n_642),
.B(n_269),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_678),
.B(n_293),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_610),
.Y(n_814)
);

AND2x2_ASAP7_75t_SL g815 ( 
.A(n_601),
.B(n_183),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_608),
.B(n_281),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_612),
.B(n_291),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_577),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_672),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_684),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_621),
.B(n_626),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_635),
.B(n_293),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_674),
.B(n_293),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_684),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_621),
.B(n_626),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_650),
.B(n_449),
.Y(n_826)
);

INVxp67_ASAP7_75t_SL g827 ( 
.A(n_580),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_635),
.B(n_446),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_666),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_610),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_623),
.B(n_303),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_623),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_624),
.B(n_332),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_624),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_584),
.A2(n_270),
.B1(n_435),
.B2(n_434),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_628),
.B(n_632),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_584),
.A2(n_436),
.B1(n_435),
.B2(n_434),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_628),
.B(n_345),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_632),
.A2(n_436),
.B(n_433),
.C(n_432),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_674),
.B(n_7),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_570),
.A2(n_356),
.B1(n_348),
.B2(n_349),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_570),
.A2(n_350),
.B1(n_430),
.B2(n_427),
.Y(n_842)
);

AND2x4_ASAP7_75t_SL g843 ( 
.A(n_652),
.B(n_183),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_638),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_638),
.B(n_432),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_660),
.A2(n_430),
.B1(n_427),
.B2(n_424),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_SL g847 ( 
.A(n_569),
.B(n_183),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_651),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_564),
.Y(n_849)
);

O2A1O1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_690),
.A2(n_693),
.B(n_729),
.C(n_728),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_743),
.B(n_622),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_750),
.A2(n_663),
.B(n_661),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_690),
.B(n_651),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_693),
.B(n_622),
.C(n_606),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_726),
.B(n_575),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_707),
.B(n_575),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_815),
.A2(n_606),
.B1(n_588),
.B2(n_644),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_815),
.A2(n_588),
.B1(n_573),
.B2(n_660),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_779),
.A2(n_676),
.B(n_679),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_708),
.Y(n_860)
);

AOI21x1_ASAP7_75t_L g861 ( 
.A1(n_773),
.A2(n_661),
.B(n_663),
.Y(n_861)
);

AND2x2_ASAP7_75t_SL g862 ( 
.A(n_843),
.B(n_601),
.Y(n_862)
);

NOR3xp33_ASAP7_75t_L g863 ( 
.A(n_732),
.B(n_681),
.C(n_670),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_694),
.B(n_588),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_699),
.B(n_557),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_691),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_685),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_697),
.B(n_557),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_687),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_698),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_735),
.B(n_664),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_697),
.B(n_630),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_750),
.A2(n_778),
.B(n_773),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_732),
.B(n_659),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_791),
.A2(n_648),
.B(n_580),
.Y(n_875)
);

O2A1O1Ixp33_ASAP7_75t_SL g876 ( 
.A1(n_725),
.A2(n_681),
.B(n_670),
.C(n_680),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_784),
.B(n_652),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_722),
.B(n_762),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_722),
.B(n_659),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_764),
.B(n_660),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_714),
.A2(n_655),
.B(n_683),
.C(n_418),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_778),
.A2(n_633),
.B(n_667),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_SL g883 ( 
.A(n_739),
.B(n_564),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_781),
.A2(n_643),
.B(n_538),
.Y(n_884)
);

AOI22x1_ASAP7_75t_L g885 ( 
.A1(n_818),
.A2(n_700),
.B1(n_711),
.B2(n_703),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_814),
.Y(n_886)
);

INVx11_ASAP7_75t_L g887 ( 
.A(n_716),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_723),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_765),
.B(n_633),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_781),
.A2(n_633),
.B(n_667),
.Y(n_890)
);

AOI21x1_ASAP7_75t_L g891 ( 
.A1(n_783),
.A2(n_796),
.B(n_794),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_701),
.B(n_706),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_783),
.A2(n_667),
.B(n_682),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_757),
.A2(n_664),
.B(n_667),
.C(n_682),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_763),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_836),
.A2(n_796),
.B(n_794),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_725),
.A2(n_742),
.B(n_727),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_687),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_712),
.B(n_620),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_691),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_742),
.A2(n_682),
.B(n_620),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_713),
.A2(n_757),
.B1(n_702),
.B2(n_714),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_801),
.A2(n_538),
.B(n_671),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_SL g904 ( 
.A1(n_840),
.A2(n_10),
.B(n_11),
.C(n_18),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_717),
.B(n_631),
.Y(n_905)
);

INVx4_ASAP7_75t_L g906 ( 
.A(n_708),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_687),
.Y(n_907)
);

INVx4_ASAP7_75t_L g908 ( 
.A(n_708),
.Y(n_908)
);

NOR2x1_ASAP7_75t_L g909 ( 
.A(n_724),
.B(n_655),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_761),
.A2(n_631),
.B1(n_655),
.B2(n_671),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_761),
.B(n_631),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_828),
.B(n_671),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_SL g913 ( 
.A(n_716),
.B(n_677),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_782),
.A2(n_639),
.B(n_677),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_695),
.A2(n_671),
.B1(n_677),
.B2(n_538),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_819),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_832),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_827),
.A2(n_639),
.B(n_677),
.Y(n_918)
);

AOI21x1_ASAP7_75t_L g919 ( 
.A1(n_801),
.A2(n_538),
.B(n_544),
.Y(n_919)
);

AOI21x1_ASAP7_75t_L g920 ( 
.A1(n_834),
.A2(n_538),
.B(n_544),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_766),
.A2(n_639),
.B(n_677),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_788),
.A2(n_10),
.B1(n_19),
.B2(n_21),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_798),
.Y(n_923)
);

OAI321xp33_ASAP7_75t_L g924 ( 
.A1(n_692),
.A2(n_785),
.A3(n_751),
.B1(n_835),
.B2(n_705),
.C(n_771),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_780),
.A2(n_671),
.B(n_602),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_730),
.B(n_602),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_802),
.B(n_602),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_789),
.A2(n_602),
.B(n_544),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_704),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_788),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_689),
.B(n_302),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_749),
.A2(n_302),
.B(n_269),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_814),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_760),
.A2(n_302),
.B(n_269),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_731),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_736),
.B(n_23),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_821),
.A2(n_302),
.B(n_269),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_775),
.A2(n_302),
.B(n_269),
.Y(n_938)
);

NAND3xp33_ASAP7_75t_L g939 ( 
.A(n_740),
.B(n_25),
.C(n_26),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_710),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_776),
.A2(n_302),
.B(n_103),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_830),
.A2(n_102),
.B(n_166),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_843),
.A2(n_795),
.B1(n_790),
.B2(n_837),
.Y(n_943)
);

OAI22xp33_ASAP7_75t_L g944 ( 
.A1(n_825),
.A2(n_25),
.B1(n_27),
.B2(n_32),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_736),
.A2(n_117),
.B(n_160),
.Y(n_945)
);

AO21x1_ASAP7_75t_L g946 ( 
.A1(n_738),
.A2(n_110),
.B(n_158),
.Y(n_946)
);

OR2x6_ASAP7_75t_SL g947 ( 
.A(n_769),
.B(n_33),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_687),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_710),
.Y(n_949)
);

NAND3xp33_ASAP7_75t_SL g950 ( 
.A(n_721),
.B(n_35),
.C(n_39),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_810),
.A2(n_35),
.B1(n_40),
.B2(n_46),
.Y(n_951)
);

BUFx12f_ASAP7_75t_L g952 ( 
.A(n_733),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_695),
.B(n_46),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_786),
.A2(n_120),
.B(n_153),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_830),
.A2(n_101),
.B(n_149),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_731),
.B(n_47),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_696),
.B(n_47),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_686),
.B(n_48),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_844),
.A2(n_123),
.B(n_147),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_844),
.A2(n_97),
.B(n_142),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_848),
.A2(n_70),
.B(n_141),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_686),
.A2(n_51),
.B(n_52),
.C(n_54),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_848),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_831),
.A2(n_833),
.B(n_838),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_718),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_718),
.Y(n_966)
);

AO21x1_ASAP7_75t_L g967 ( 
.A1(n_738),
.A2(n_840),
.B(n_812),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_734),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_734),
.A2(n_124),
.B(n_140),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_803),
.B(n_51),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_696),
.B(n_813),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_737),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_813),
.B(n_54),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_754),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_720),
.B(n_758),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_823),
.B(n_55),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_746),
.B(n_56),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_805),
.B(n_60),
.Y(n_978)
);

AND2x2_ASAP7_75t_SL g979 ( 
.A(n_733),
.B(n_63),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_737),
.A2(n_68),
.B(n_127),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_724),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_741),
.Y(n_982)
);

CKINVDCx11_ASAP7_75t_R g983 ( 
.A(n_849),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_741),
.A2(n_132),
.B(n_136),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_823),
.B(n_139),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_767),
.A2(n_172),
.B(n_797),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_792),
.B(n_753),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_744),
.B(n_748),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_767),
.A2(n_797),
.B(n_824),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_745),
.B(n_747),
.Y(n_990)
);

AOI21x1_ASAP7_75t_L g991 ( 
.A1(n_787),
.A2(n_808),
.B(n_804),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_822),
.B(n_759),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_752),
.B(n_756),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_689),
.B(n_733),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_715),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_770),
.A2(n_793),
.B1(n_806),
.B2(n_755),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_787),
.B(n_808),
.Y(n_997)
);

AND2x6_ASAP7_75t_SL g998 ( 
.A(n_719),
.B(n_688),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_689),
.B(n_804),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_820),
.B(n_824),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_820),
.A2(n_774),
.B(n_807),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_709),
.A2(n_816),
.B(n_817),
.C(n_811),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_845),
.A2(n_809),
.B(n_800),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_799),
.A2(n_772),
.B(n_839),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_829),
.Y(n_1005)
);

OAI321xp33_ASAP7_75t_L g1006 ( 
.A1(n_826),
.A2(n_768),
.A3(n_719),
.B1(n_842),
.B2(n_846),
.C(n_841),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_719),
.A2(n_777),
.B(n_689),
.C(n_847),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_690),
.B(n_693),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_689),
.B(n_815),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_779),
.A2(n_543),
.B(n_791),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_779),
.A2(n_543),
.B(n_791),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_715),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_779),
.A2(n_543),
.B(n_791),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_779),
.A2(n_543),
.B(n_791),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_690),
.B(n_693),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_779),
.A2(n_543),
.B(n_791),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_750),
.A2(n_547),
.B(n_568),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_690),
.A2(n_693),
.B(n_552),
.C(n_728),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_779),
.A2(n_543),
.B(n_791),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_685),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_690),
.A2(n_693),
.B1(n_815),
.B2(n_552),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_779),
.A2(n_543),
.B(n_791),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_716),
.Y(n_1023)
);

AOI21x1_ASAP7_75t_L g1024 ( 
.A1(n_773),
.A2(n_781),
.B(n_778),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_690),
.B(n_693),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_690),
.B(n_693),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_779),
.A2(n_543),
.B(n_791),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_687),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_779),
.A2(n_543),
.B(n_791),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_SL g1030 ( 
.A1(n_690),
.A2(n_693),
.B(n_727),
.C(n_725),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1018),
.C(n_1025),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_891),
.A2(n_1024),
.B(n_920),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_999),
.A2(n_852),
.B(n_919),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1015),
.B(n_878),
.Y(n_1035)
);

NAND2x1_ASAP7_75t_L g1036 ( 
.A(n_869),
.B(n_1028),
.Y(n_1036)
);

AO21x2_ASAP7_75t_L g1037 ( 
.A1(n_937),
.A2(n_902),
.B(n_894),
.Y(n_1037)
);

AO221x1_ASAP7_75t_L g1038 ( 
.A1(n_1021),
.A2(n_944),
.B1(n_922),
.B2(n_930),
.C(n_951),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_851),
.B(n_979),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_971),
.B(n_892),
.Y(n_1040)
);

AOI21x1_ASAP7_75t_L g1041 ( 
.A1(n_985),
.A2(n_967),
.B(n_897),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_867),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_898),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_850),
.B(n_975),
.Y(n_1044)
);

AOI21x1_ASAP7_75t_SL g1045 ( 
.A1(n_976),
.A2(n_973),
.B(n_957),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_874),
.B(n_879),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_887),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_988),
.B(n_990),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1017),
.A2(n_873),
.B(n_1002),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_860),
.Y(n_1050)
);

NAND2x1_ASAP7_75t_L g1051 ( 
.A(n_869),
.B(n_1028),
.Y(n_1051)
);

AOI21xp33_ASAP7_75t_L g1052 ( 
.A1(n_953),
.A2(n_936),
.B(n_958),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_993),
.B(n_853),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_SL g1054 ( 
.A1(n_885),
.A2(n_945),
.B(n_1007),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_958),
.A2(n_857),
.B1(n_854),
.B2(n_862),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_964),
.A2(n_1030),
.B(n_872),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_860),
.B(n_906),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_931),
.A2(n_1003),
.B(n_890),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1002),
.A2(n_1001),
.B(n_1010),
.Y(n_1059)
);

AND3x4_ASAP7_75t_L g1060 ( 
.A(n_1023),
.B(n_909),
.C(n_956),
.Y(n_1060)
);

OR2x6_ASAP7_75t_L g1061 ( 
.A(n_952),
.B(n_994),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_906),
.B(n_908),
.Y(n_1062)
);

AND3x1_ASAP7_75t_SL g1063 ( 
.A(n_870),
.B(n_1020),
.C(n_888),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_908),
.B(n_935),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_882),
.A2(n_896),
.B(n_928),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_1011),
.A2(n_1016),
.B(n_1029),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1030),
.A2(n_868),
.B(n_875),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_911),
.A2(n_1027),
.B(n_1022),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1013),
.A2(n_1019),
.B(n_1014),
.Y(n_1069)
);

AO31x2_ASAP7_75t_L g1070 ( 
.A1(n_894),
.A2(n_946),
.A3(n_864),
.B(n_938),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_950),
.A2(n_944),
.B(n_962),
.C(n_904),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_978),
.B(n_856),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_935),
.B(n_994),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_862),
.B(n_916),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_L g1075 ( 
.A(n_863),
.B(n_978),
.C(n_904),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_880),
.B(n_917),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_889),
.A2(n_865),
.B(n_859),
.Y(n_1077)
);

AO21x1_ASAP7_75t_L g1078 ( 
.A1(n_1009),
.A2(n_934),
.B(n_863),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_979),
.B(n_877),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_923),
.B(n_992),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_925),
.A2(n_986),
.B(n_921),
.Y(n_1081)
);

NAND3xp33_ASAP7_75t_SL g1082 ( 
.A(n_883),
.B(n_871),
.C(n_981),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_942),
.A2(n_959),
.B(n_893),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_926),
.A2(n_876),
.B(n_987),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1004),
.A2(n_941),
.B(n_932),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_881),
.A2(n_996),
.B(n_924),
.C(n_1006),
.Y(n_1086)
);

OR2x6_ASAP7_75t_L g1087 ( 
.A(n_1012),
.B(n_1023),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_903),
.A2(n_884),
.B(n_914),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_963),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_918),
.A2(n_1000),
.B(n_997),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_910),
.A2(n_858),
.B(n_970),
.C(n_977),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_1005),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_876),
.A2(n_901),
.B(n_954),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_898),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_855),
.B(n_995),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1009),
.A2(n_905),
.B(n_899),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_995),
.B(n_977),
.Y(n_1097)
);

INVx3_ASAP7_75t_SL g1098 ( 
.A(n_895),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_956),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_898),
.A2(n_948),
.B(n_907),
.Y(n_1100)
);

OAI21xp33_ASAP7_75t_SL g1101 ( 
.A1(n_943),
.A2(n_915),
.B(n_912),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_927),
.B(n_913),
.Y(n_1102)
);

AO31x2_ASAP7_75t_L g1103 ( 
.A1(n_900),
.A2(n_949),
.A3(n_982),
.B(n_966),
.Y(n_1103)
);

OR2x6_ASAP7_75t_L g1104 ( 
.A(n_886),
.B(n_933),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_929),
.A2(n_961),
.B(n_984),
.Y(n_1105)
);

AOI21xp33_ASAP7_75t_L g1106 ( 
.A1(n_943),
.A2(n_965),
.B(n_972),
.Y(n_1106)
);

NAND2x1_ASAP7_75t_L g1107 ( 
.A(n_898),
.B(n_907),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_907),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_907),
.Y(n_1109)
);

AO31x2_ASAP7_75t_L g1110 ( 
.A1(n_968),
.A2(n_940),
.A3(n_960),
.B(n_955),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_948),
.B(n_974),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_947),
.B(n_983),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_948),
.B(n_998),
.Y(n_1113)
);

BUFx4f_ASAP7_75t_L g1114 ( 
.A(n_948),
.Y(n_1114)
);

INVx6_ASAP7_75t_L g1115 ( 
.A(n_983),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_939),
.B(n_974),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_974),
.B(n_969),
.Y(n_1117)
);

AO21x1_ASAP7_75t_L g1118 ( 
.A1(n_980),
.A2(n_1026),
.B(n_1008),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_974),
.A2(n_1026),
.B(n_1008),
.C(n_1025),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1021),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1021),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_983),
.Y(n_1124)
);

OAI21xp33_ASAP7_75t_SL g1125 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1025),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1025),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1021),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_851),
.B(n_743),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_861),
.A2(n_991),
.B(n_989),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_861),
.A2(n_991),
.B(n_989),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_861),
.A2(n_991),
.B(n_989),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_866),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1025),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_866),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1021),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1018),
.C(n_1025),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_866),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1143)
);

NAND2x1p5_ASAP7_75t_L g1144 ( 
.A(n_860),
.B(n_906),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1012),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_861),
.A2(n_991),
.B(n_989),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1025),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_983),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_861),
.A2(n_991),
.B(n_989),
.Y(n_1151)
);

NAND2x1p5_ASAP7_75t_L g1152 ( 
.A(n_860),
.B(n_906),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_861),
.A2(n_991),
.B(n_989),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1025),
.Y(n_1155)
);

NOR2xp67_ASAP7_75t_L g1156 ( 
.A(n_995),
.B(n_562),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1008),
.A2(n_1026),
.B1(n_1021),
.B2(n_1025),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1025),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_861),
.A2(n_991),
.B(n_989),
.Y(n_1161)
);

NAND2x1p5_ASAP7_75t_L g1162 ( 
.A(n_860),
.B(n_906),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_860),
.B(n_906),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_866),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_SL g1165 ( 
.A1(n_1021),
.A2(n_1025),
.B(n_1015),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_902),
.A2(n_967),
.A3(n_894),
.B(n_1002),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_861),
.A2(n_991),
.B(n_989),
.Y(n_1167)
);

AOI21x1_ASAP7_75t_SL g1168 ( 
.A1(n_1015),
.A2(n_1025),
.B(n_976),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_861),
.A2(n_991),
.B(n_989),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_R g1170 ( 
.A(n_981),
.B(n_649),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_SL g1172 ( 
.A1(n_1021),
.A2(n_902),
.B(n_1008),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1018),
.C(n_1025),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1005),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1177)
);

INVx5_ASAP7_75t_L g1178 ( 
.A(n_1061),
.Y(n_1178)
);

AOI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_1149),
.A2(n_1174),
.B1(n_1140),
.B2(n_1141),
.C(n_1122),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1057),
.B(n_1062),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1039),
.B(n_1128),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1122),
.A2(n_1177),
.B1(n_1159),
.B2(n_1158),
.Y(n_1182)
);

O2A1O1Ixp5_ASAP7_75t_L g1183 ( 
.A1(n_1120),
.A2(n_1135),
.B(n_1127),
.C(n_1123),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1042),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1145),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_1148),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1172),
.A2(n_1123),
.B(n_1120),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1177),
.B(n_1140),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1127),
.A2(n_1135),
.B(n_1133),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_L g1190 ( 
.A(n_1157),
.B(n_1147),
.C(n_1126),
.Y(n_1190)
);

NAND2x1_ASAP7_75t_L g1191 ( 
.A(n_1043),
.B(n_1094),
.Y(n_1191)
);

OAI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1034),
.A2(n_1142),
.B1(n_1173),
.B2(n_1136),
.Y(n_1192)
);

INVxp67_ASAP7_75t_L g1193 ( 
.A(n_1176),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1095),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1143),
.B(n_1141),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1155),
.A2(n_1160),
.B(n_1138),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1079),
.B(n_1048),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1031),
.A2(n_1175),
.B(n_1154),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1170),
.Y(n_1199)
);

NAND2xp33_ASAP7_75t_L g1200 ( 
.A(n_1150),
.B(n_1154),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1150),
.B(n_1158),
.Y(n_1201)
);

NAND2x1p5_ASAP7_75t_L g1202 ( 
.A(n_1114),
.B(n_1064),
.Y(n_1202)
);

OA21x2_ASAP7_75t_L g1203 ( 
.A1(n_1059),
.A2(n_1056),
.B(n_1066),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1092),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1159),
.A2(n_1125),
.B(n_1119),
.C(n_1052),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1087),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1121),
.A2(n_1137),
.B(n_1171),
.C(n_1052),
.Y(n_1207)
);

NAND2x1p5_ASAP7_75t_L g1208 ( 
.A(n_1114),
.B(n_1064),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1080),
.B(n_1099),
.Y(n_1209)
);

AND2x2_ASAP7_75t_SL g1210 ( 
.A(n_1074),
.B(n_1112),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_1057),
.B(n_1062),
.Y(n_1211)
);

INVx4_ASAP7_75t_L g1212 ( 
.A(n_1047),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1061),
.B(n_1050),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_1111),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1061),
.B(n_1050),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1087),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1040),
.B(n_1035),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1097),
.A2(n_1055),
.B1(n_1074),
.B2(n_1072),
.Y(n_1218)
);

AOI221x1_ASAP7_75t_L g1219 ( 
.A1(n_1086),
.A2(n_1075),
.B1(n_1055),
.B2(n_1165),
.C(n_1049),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1040),
.A2(n_1071),
.B(n_1075),
.C(n_1044),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1073),
.B(n_1113),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1044),
.A2(n_1091),
.B(n_1053),
.C(n_1054),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1053),
.B(n_1046),
.Y(n_1223)
);

NAND2x1p5_ASAP7_75t_L g1224 ( 
.A(n_1073),
.B(n_1107),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1089),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1132),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_SL g1227 ( 
.A(n_1060),
.B(n_1082),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1134),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1124),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1047),
.B(n_1104),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1104),
.B(n_1156),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1043),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_1111),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1115),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1098),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1139),
.Y(n_1236)
);

INVxp67_ASAP7_75t_L g1237 ( 
.A(n_1104),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1067),
.A2(n_1085),
.B(n_1068),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1144),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_1116),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1076),
.A2(n_1049),
.B1(n_1046),
.B2(n_1085),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1069),
.A2(n_1059),
.B(n_1118),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1043),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1101),
.A2(n_1076),
.B(n_1084),
.C(n_1106),
.Y(n_1244)
);

BUFx12f_ASAP7_75t_L g1245 ( 
.A(n_1094),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1152),
.Y(n_1246)
);

AND2x6_ASAP7_75t_L g1247 ( 
.A(n_1094),
.B(n_1108),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1108),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1037),
.B(n_1164),
.Y(n_1249)
);

AO21x1_ASAP7_75t_L g1250 ( 
.A1(n_1106),
.A2(n_1096),
.B(n_1093),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1108),
.Y(n_1251)
);

AOI21x1_ASAP7_75t_SL g1252 ( 
.A1(n_1117),
.A2(n_1168),
.B(n_1045),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_1109),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1093),
.A2(n_1078),
.B(n_1037),
.C(n_1077),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1117),
.A2(n_1033),
.B(n_1088),
.C(n_1102),
.Y(n_1255)
);

CKINVDCx8_ASAP7_75t_R g1256 ( 
.A(n_1063),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1152),
.B(n_1162),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1163),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1163),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1036),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1051),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1103),
.B(n_1166),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1038),
.B(n_1166),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1166),
.B(n_1103),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1100),
.B(n_1041),
.Y(n_1265)
);

NAND2xp33_ASAP7_75t_L g1266 ( 
.A(n_1070),
.B(n_1065),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1058),
.A2(n_1081),
.B(n_1105),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1090),
.B(n_1110),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1110),
.B(n_1032),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1129),
.B(n_1151),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1130),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1131),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1083),
.A2(n_1169),
.B(n_1153),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1146),
.A2(n_1161),
.B(n_1167),
.Y(n_1274)
);

INVxp67_ASAP7_75t_SL g1275 ( 
.A(n_1149),
.Y(n_1275)
);

NOR2xp67_ASAP7_75t_L g1276 ( 
.A(n_1047),
.B(n_562),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1149),
.A2(n_1008),
.B1(n_1026),
.B2(n_531),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1114),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1176),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1176),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1149),
.B(n_1174),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1172),
.A2(n_1123),
.B(n_1120),
.Y(n_1282)
);

INVx3_ASAP7_75t_SL g1283 ( 
.A(n_1148),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1176),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1039),
.B(n_1128),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1042),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1170),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1039),
.B(n_1128),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1149),
.A2(n_1026),
.B(n_1008),
.C(n_1174),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1176),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1114),
.B(n_731),
.Y(n_1291)
);

OR2x6_ASAP7_75t_L g1292 ( 
.A(n_1061),
.B(n_708),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1122),
.B(n_1141),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1057),
.B(n_1062),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1172),
.A2(n_1123),
.B(n_1120),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1149),
.B(n_1174),
.Y(n_1296)
);

NAND2xp33_ASAP7_75t_L g1297 ( 
.A(n_1120),
.B(n_1123),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1172),
.A2(n_1123),
.B(n_1120),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1039),
.B(n_1128),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1172),
.A2(n_1123),
.B(n_1120),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1122),
.B(n_1141),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1172),
.A2(n_1123),
.B(n_1120),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1149),
.A2(n_1174),
.B1(n_1122),
.B2(n_1141),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1042),
.Y(n_1304)
);

INVxp67_ASAP7_75t_L g1305 ( 
.A(n_1176),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1120),
.A2(n_1127),
.B(n_1123),
.Y(n_1306)
);

INVx5_ASAP7_75t_L g1307 ( 
.A(n_1061),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1176),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1149),
.B(n_1174),
.Y(n_1309)
);

AND2x2_ASAP7_75t_SL g1310 ( 
.A(n_1149),
.B(n_815),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1149),
.B(n_1008),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1145),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1114),
.Y(n_1313)
);

NOR2x1_ASAP7_75t_SL g1314 ( 
.A(n_1061),
.B(n_1104),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1149),
.A2(n_1008),
.B(n_1026),
.C(n_1174),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1122),
.B(n_1141),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1114),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1149),
.A2(n_1026),
.B(n_1008),
.C(n_1174),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1145),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1042),
.Y(n_1320)
);

OR2x6_ASAP7_75t_SL g1321 ( 
.A(n_1148),
.B(n_649),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1122),
.B(n_1141),
.Y(n_1322)
);

NOR2xp67_ASAP7_75t_L g1323 ( 
.A(n_1047),
.B(n_562),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1310),
.A2(n_1227),
.B1(n_1281),
.B2(n_1309),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1184),
.Y(n_1325)
);

AO21x1_ASAP7_75t_L g1326 ( 
.A1(n_1187),
.A2(n_1295),
.B(n_1282),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1192),
.B(n_1179),
.Y(n_1327)
);

AO21x1_ASAP7_75t_L g1328 ( 
.A1(n_1298),
.A2(n_1302),
.B(n_1300),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1296),
.B(n_1195),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1277),
.A2(n_1179),
.B1(n_1227),
.B2(n_1311),
.Y(n_1330)
);

BUFx10_ASAP7_75t_L g1331 ( 
.A(n_1199),
.Y(n_1331)
);

AO21x2_ASAP7_75t_L g1332 ( 
.A1(n_1274),
.A2(n_1273),
.B(n_1264),
.Y(n_1332)
);

OR2x6_ASAP7_75t_L g1333 ( 
.A(n_1292),
.B(n_1249),
.Y(n_1333)
);

CKINVDCx6p67_ASAP7_75t_R g1334 ( 
.A(n_1321),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1275),
.A2(n_1303),
.B1(n_1197),
.B2(n_1181),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1303),
.A2(n_1210),
.B1(n_1182),
.B2(n_1306),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1245),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1286),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1201),
.B(n_1217),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1229),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1180),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1203),
.Y(n_1342)
);

AOI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1267),
.A2(n_1242),
.B(n_1238),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1185),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1304),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1247),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1320),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1315),
.A2(n_1289),
.B1(n_1318),
.B2(n_1306),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1194),
.A2(n_1218),
.B1(n_1299),
.B2(n_1285),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1194),
.A2(n_1288),
.B1(n_1223),
.B2(n_1182),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1225),
.Y(n_1351)
);

INVx3_ASAP7_75t_SL g1352 ( 
.A(n_1235),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1254),
.A2(n_1268),
.B(n_1270),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1223),
.A2(n_1198),
.B1(n_1297),
.B2(n_1217),
.Y(n_1354)
);

INVxp67_ASAP7_75t_SL g1355 ( 
.A(n_1222),
.Y(n_1355)
);

BUFx8_ASAP7_75t_L g1356 ( 
.A(n_1287),
.Y(n_1356)
);

AO21x1_ASAP7_75t_SL g1357 ( 
.A1(n_1263),
.A2(n_1198),
.B(n_1268),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1264),
.Y(n_1358)
);

INVx6_ASAP7_75t_L g1359 ( 
.A(n_1180),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1262),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1203),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1263),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1219),
.A2(n_1270),
.B(n_1189),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1226),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1228),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1196),
.A2(n_1252),
.B(n_1271),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1271),
.A2(n_1272),
.B(n_1269),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1236),
.Y(n_1368)
);

AO21x1_ASAP7_75t_SL g1369 ( 
.A1(n_1183),
.A2(n_1293),
.B(n_1322),
.Y(n_1369)
);

BUFx8_ASAP7_75t_L g1370 ( 
.A(n_1186),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1214),
.B(n_1233),
.Y(n_1371)
);

INVx4_ASAP7_75t_SL g1372 ( 
.A(n_1292),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1248),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1314),
.A2(n_1190),
.B1(n_1200),
.B2(n_1178),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1214),
.B(n_1233),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1240),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1240),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1221),
.A2(n_1188),
.B1(n_1293),
.B2(n_1322),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1221),
.A2(n_1188),
.B1(n_1301),
.B2(n_1316),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1205),
.B(n_1241),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1312),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1248),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1241),
.B(n_1316),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1206),
.Y(n_1384)
);

AO21x1_ASAP7_75t_SL g1385 ( 
.A1(n_1301),
.A2(n_1190),
.B(n_1257),
.Y(n_1385)
);

AOI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1250),
.A2(n_1260),
.B(n_1191),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1319),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1209),
.A2(n_1231),
.B1(n_1307),
.B2(n_1216),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1248),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1237),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1220),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1290),
.B(n_1308),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1244),
.A2(n_1255),
.B(n_1265),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1256),
.A2(n_1308),
.B1(n_1290),
.B2(n_1307),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1224),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1231),
.A2(n_1204),
.B1(n_1280),
.B2(n_1284),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1193),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1230),
.A2(n_1305),
.B1(n_1215),
.B2(n_1213),
.Y(n_1398)
);

AOI21xp33_ASAP7_75t_L g1399 ( 
.A1(n_1207),
.A2(n_1266),
.B(n_1261),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1232),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1294),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1243),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1251),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1234),
.A2(n_1317),
.B1(n_1313),
.B2(n_1278),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1259),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1283),
.A2(n_1253),
.B1(n_1212),
.B2(n_1211),
.Y(n_1406)
);

BUFx2_ASAP7_75t_R g1407 ( 
.A(n_1239),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1323),
.A2(n_1276),
.B1(n_1208),
.B2(n_1202),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1258),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1258),
.B(n_1246),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1313),
.A2(n_1317),
.B1(n_1291),
.B2(n_1212),
.Y(n_1411)
);

AO21x1_ASAP7_75t_L g1412 ( 
.A1(n_1187),
.A2(n_1021),
.B(n_1008),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1310),
.A2(n_1277),
.B1(n_1008),
.B2(n_1026),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1249),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1249),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1184),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1279),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1249),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1315),
.A2(n_1174),
.B1(n_1149),
.B2(n_1026),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1247),
.Y(n_1420)
);

AOI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1267),
.A2(n_1242),
.B(n_1238),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1306),
.B(n_1197),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1199),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1184),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1290),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1203),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1184),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1203),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1279),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1184),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1199),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1274),
.A2(n_1273),
.B(n_1264),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1203),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1315),
.A2(n_1174),
.B1(n_1149),
.B2(n_1026),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_1340),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1329),
.B(n_1339),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1422),
.B(n_1357),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1358),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1352),
.B(n_1324),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1386),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1354),
.B(n_1422),
.Y(n_1441)
);

INVx6_ASAP7_75t_L g1442 ( 
.A(n_1356),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1414),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1413),
.A2(n_1327),
.B1(n_1330),
.B2(n_1419),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1414),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1342),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1415),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1415),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1417),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1429),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1362),
.B(n_1360),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1418),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1343),
.A2(n_1421),
.B(n_1366),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1353),
.A2(n_1328),
.B(n_1326),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1386),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1418),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1412),
.A2(n_1361),
.B(n_1343),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1357),
.B(n_1383),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1425),
.B(n_1391),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1378),
.B(n_1379),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1362),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1336),
.A2(n_1434),
.B1(n_1380),
.B2(n_1376),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1372),
.B(n_1333),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1348),
.A2(n_1355),
.B1(n_1380),
.B2(n_1350),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1367),
.A2(n_1328),
.B(n_1326),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1383),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1325),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1374),
.A2(n_1399),
.B(n_1392),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1335),
.B(n_1397),
.Y(n_1469)
);

BUFx8_ASAP7_75t_SL g1470 ( 
.A(n_1340),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1342),
.B(n_1426),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1431),
.Y(n_1472)
);

INVx1_ASAP7_75t_SL g1473 ( 
.A(n_1344),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1403),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1403),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1431),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1400),
.B(n_1405),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1338),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1345),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1347),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1351),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1344),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1402),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1416),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1371),
.B(n_1375),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1424),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1393),
.A2(n_1408),
.B(n_1394),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1384),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1405),
.B(n_1427),
.Y(n_1489)
);

OA21x2_ASAP7_75t_L g1490 ( 
.A1(n_1412),
.A2(n_1361),
.B(n_1367),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1430),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1428),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1371),
.B(n_1375),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1433),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1433),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1349),
.B(n_1377),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1396),
.B(n_1368),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1369),
.B(n_1363),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1364),
.Y(n_1499)
);

OAI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1393),
.A2(n_1411),
.B(n_1363),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1365),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1390),
.Y(n_1502)
);

AO21x2_ASAP7_75t_L g1503 ( 
.A1(n_1332),
.A2(n_1432),
.B(n_1395),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1393),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1332),
.B(n_1432),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1346),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1369),
.B(n_1385),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1458),
.B(n_1385),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1482),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1466),
.B(n_1373),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1437),
.B(n_1373),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1507),
.B(n_1372),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1492),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1467),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1471),
.B(n_1389),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1471),
.B(n_1389),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1467),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1498),
.B(n_1382),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1461),
.B(n_1382),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1485),
.B(n_1334),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1492),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1446),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1485),
.B(n_1493),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1498),
.B(n_1334),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1461),
.B(n_1420),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1446),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1454),
.B(n_1346),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1454),
.B(n_1381),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1494),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1493),
.B(n_1387),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1474),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_L g1532 ( 
.A(n_1444),
.B(n_1398),
.C(n_1356),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1454),
.B(n_1387),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1482),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1443),
.B(n_1409),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1454),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1464),
.B(n_1406),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1495),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1503),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1490),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1462),
.A2(n_1359),
.B1(n_1341),
.B2(n_1401),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1490),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1505),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1451),
.B(n_1410),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1451),
.B(n_1410),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1473),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1514),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1528),
.B(n_1504),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_SL g1549 ( 
.A1(n_1537),
.A2(n_1439),
.B(n_1468),
.Y(n_1549)
);

NAND3xp33_ASAP7_75t_L g1550 ( 
.A(n_1537),
.B(n_1469),
.C(n_1500),
.Y(n_1550)
);

OAI21xp33_ASAP7_75t_L g1551 ( 
.A1(n_1528),
.A2(n_1441),
.B(n_1459),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1531),
.B(n_1449),
.Y(n_1552)
);

AOI211xp5_ASAP7_75t_L g1553 ( 
.A1(n_1528),
.A2(n_1487),
.B(n_1436),
.C(n_1489),
.Y(n_1553)
);

OAI21xp5_ASAP7_75t_SL g1554 ( 
.A1(n_1508),
.A2(n_1475),
.B(n_1477),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1533),
.B(n_1504),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1531),
.B(n_1450),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1533),
.B(n_1506),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1532),
.A2(n_1460),
.B1(n_1496),
.B2(n_1497),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1546),
.B(n_1502),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1546),
.B(n_1483),
.Y(n_1560)
);

NAND3xp33_ASAP7_75t_L g1561 ( 
.A(n_1540),
.B(n_1488),
.C(n_1445),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1508),
.B(n_1506),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1523),
.B(n_1438),
.Y(n_1563)
);

NOR3xp33_ASAP7_75t_L g1564 ( 
.A(n_1536),
.B(n_1455),
.C(n_1440),
.Y(n_1564)
);

NAND3xp33_ASAP7_75t_L g1565 ( 
.A(n_1540),
.B(n_1447),
.C(n_1456),
.Y(n_1565)
);

NAND3xp33_ASAP7_75t_L g1566 ( 
.A(n_1542),
.B(n_1447),
.C(n_1456),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1508),
.B(n_1506),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1544),
.B(n_1448),
.Y(n_1568)
);

OAI21xp33_ASAP7_75t_L g1569 ( 
.A1(n_1542),
.A2(n_1525),
.B(n_1536),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1515),
.B(n_1478),
.Y(n_1570)
);

NOR3xp33_ASAP7_75t_SL g1571 ( 
.A(n_1519),
.B(n_1472),
.C(n_1476),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1514),
.Y(n_1572)
);

OA21x2_ASAP7_75t_L g1573 ( 
.A1(n_1539),
.A2(n_1465),
.B(n_1453),
.Y(n_1573)
);

NOR3xp33_ASAP7_75t_L g1574 ( 
.A(n_1536),
.B(n_1440),
.C(n_1455),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1541),
.A2(n_1442),
.B1(n_1435),
.B2(n_1388),
.Y(n_1575)
);

NAND3xp33_ASAP7_75t_L g1576 ( 
.A(n_1525),
.B(n_1452),
.C(n_1448),
.Y(n_1576)
);

NOR3xp33_ASAP7_75t_L g1577 ( 
.A(n_1536),
.B(n_1455),
.C(n_1440),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_L g1578 ( 
.A(n_1519),
.B(n_1452),
.C(n_1499),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_SL g1579 ( 
.A1(n_1524),
.A2(n_1505),
.B(n_1404),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1517),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_L g1581 ( 
.A(n_1536),
.B(n_1499),
.C(n_1501),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1544),
.B(n_1545),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1517),
.Y(n_1583)
);

NAND3xp33_ASAP7_75t_L g1584 ( 
.A(n_1513),
.B(n_1501),
.C(n_1484),
.Y(n_1584)
);

NOR3xp33_ASAP7_75t_L g1585 ( 
.A(n_1535),
.B(n_1465),
.C(n_1479),
.Y(n_1585)
);

AND2x2_ASAP7_75t_SL g1586 ( 
.A(n_1512),
.B(n_1463),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1516),
.B(n_1479),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1545),
.B(n_1480),
.Y(n_1588)
);

OAI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1520),
.A2(n_1480),
.B1(n_1481),
.B2(n_1491),
.C(n_1486),
.Y(n_1589)
);

NAND3xp33_ASAP7_75t_L g1590 ( 
.A(n_1513),
.B(n_1491),
.C(n_1486),
.Y(n_1590)
);

NAND4xp25_ASAP7_75t_L g1591 ( 
.A(n_1522),
.B(n_1526),
.C(n_1524),
.D(n_1538),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1516),
.B(n_1457),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1547),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1572),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1557),
.B(n_1522),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1549),
.B(n_1352),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1580),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1583),
.Y(n_1598)
);

NOR4xp25_ASAP7_75t_L g1599 ( 
.A(n_1550),
.B(n_1530),
.C(n_1510),
.D(n_1543),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1584),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1553),
.B(n_1509),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1592),
.B(n_1521),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1548),
.Y(n_1603)
);

NOR2x1_ASAP7_75t_L g1604 ( 
.A(n_1591),
.B(n_1509),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1590),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1582),
.B(n_1529),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1581),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1563),
.B(n_1529),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1578),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1585),
.B(n_1529),
.Y(n_1610)
);

NAND2x1_ASAP7_75t_L g1611 ( 
.A(n_1555),
.B(n_1538),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1565),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1588),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1573),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1573),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1573),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1570),
.B(n_1511),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1576),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1562),
.B(n_1526),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1562),
.B(n_1527),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1587),
.B(n_1527),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1568),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1586),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1567),
.B(n_1527),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1618),
.B(n_1609),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1620),
.B(n_1587),
.Y(n_1626)
);

OAI21xp33_ASAP7_75t_L g1627 ( 
.A1(n_1607),
.A2(n_1569),
.B(n_1556),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1618),
.B(n_1609),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1604),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1620),
.B(n_1554),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1620),
.B(n_1567),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1593),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1600),
.B(n_1552),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1620),
.B(n_1564),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1600),
.B(n_1566),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1605),
.B(n_1612),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1614),
.Y(n_1637)
);

NAND2xp33_ASAP7_75t_L g1638 ( 
.A(n_1604),
.B(n_1571),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1614),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1605),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1593),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1624),
.B(n_1574),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1606),
.B(n_1559),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1614),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1624),
.B(n_1534),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1594),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1594),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1615),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1624),
.B(n_1577),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1606),
.B(n_1560),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1607),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1597),
.Y(n_1652)
);

OAI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1623),
.A2(n_1612),
.B1(n_1601),
.B2(n_1579),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1608),
.B(n_1561),
.Y(n_1654)
);

AND2x4_ASAP7_75t_SL g1655 ( 
.A(n_1623),
.B(n_1512),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1621),
.B(n_1603),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1615),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1621),
.B(n_1518),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1597),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1621),
.B(n_1518),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1598),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1611),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1632),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1632),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1633),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1641),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1641),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1625),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1653),
.A2(n_1596),
.B1(n_1558),
.B2(n_1603),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1640),
.A2(n_1558),
.B1(n_1551),
.B2(n_1575),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1637),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1646),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1646),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1637),
.Y(n_1674)
);

NAND4xp25_ASAP7_75t_L g1675 ( 
.A(n_1636),
.B(n_1651),
.C(n_1628),
.D(n_1625),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1628),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1651),
.B(n_1599),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1636),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1635),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1635),
.Y(n_1680)
);

INVx1_ASAP7_75t_SL g1681 ( 
.A(n_1633),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1630),
.B(n_1617),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1647),
.Y(n_1683)
);

NAND2x1_ASAP7_75t_L g1684 ( 
.A(n_1629),
.B(n_1619),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1647),
.Y(n_1685)
);

NAND2x1_ASAP7_75t_L g1686 ( 
.A(n_1629),
.B(n_1619),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1652),
.Y(n_1687)
);

NAND2x1p5_ASAP7_75t_L g1688 ( 
.A(n_1662),
.B(n_1586),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1640),
.B(n_1470),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1638),
.A2(n_1599),
.B(n_1610),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1630),
.B(n_1617),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1630),
.A2(n_1610),
.B1(n_1611),
.B2(n_1595),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1652),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1655),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1659),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1656),
.B(n_1595),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1659),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1627),
.B(n_1613),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1627),
.B(n_1613),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1637),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1643),
.B(n_1472),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1626),
.B(n_1656),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1661),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1639),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1661),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1682),
.B(n_1656),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1702),
.Y(n_1707)
);

NOR2x1_ASAP7_75t_L g1708 ( 
.A(n_1675),
.B(n_1634),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1676),
.B(n_1654),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1689),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1663),
.Y(n_1711)
);

NOR2x1_ASAP7_75t_L g1712 ( 
.A(n_1676),
.B(n_1634),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1664),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1688),
.B(n_1662),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1666),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1677),
.A2(n_1639),
.B1(n_1644),
.B2(n_1657),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1681),
.B(n_1654),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1665),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1679),
.B(n_1643),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1689),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1701),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_1694),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1667),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1682),
.B(n_1634),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_L g1725 ( 
.A(n_1690),
.B(n_1616),
.C(n_1615),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1672),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1691),
.B(n_1642),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1701),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1673),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1691),
.B(n_1642),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1683),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1702),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1680),
.B(n_1678),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1696),
.B(n_1642),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1698),
.B(n_1650),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1668),
.B(n_1370),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1685),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1687),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1688),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1693),
.Y(n_1740)
);

OAI21x1_ASAP7_75t_L g1741 ( 
.A1(n_1684),
.A2(n_1644),
.B(n_1639),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1718),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1708),
.A2(n_1669),
.B(n_1699),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1712),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1711),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1725),
.A2(n_1670),
.B1(n_1674),
.B2(n_1671),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1709),
.B(n_1695),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1724),
.B(n_1694),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1711),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1713),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1713),
.Y(n_1751)
);

NAND3xp33_ASAP7_75t_L g1752 ( 
.A(n_1712),
.B(n_1705),
.C(n_1703),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1708),
.A2(n_1717),
.B1(n_1688),
.B2(n_1707),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1717),
.B(n_1697),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1741),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1719),
.B(n_1626),
.Y(n_1756)
);

O2A1O1Ixp33_ASAP7_75t_SL g1757 ( 
.A1(n_1710),
.A2(n_1684),
.B(n_1686),
.C(n_1662),
.Y(n_1757)
);

AOI32xp33_ASAP7_75t_L g1758 ( 
.A1(n_1739),
.A2(n_1692),
.A3(n_1649),
.B1(n_1616),
.B2(n_1696),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1736),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1724),
.B(n_1696),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1741),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1714),
.A2(n_1686),
.B(n_1649),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1707),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1719),
.B(n_1626),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1727),
.B(n_1649),
.Y(n_1765)
);

INVx1_ASAP7_75t_SL g1766 ( 
.A(n_1720),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1715),
.Y(n_1767)
);

AO22x1_ASAP7_75t_L g1768 ( 
.A1(n_1753),
.A2(n_1728),
.B1(n_1739),
.B2(n_1721),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1766),
.B(n_1727),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1745),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1760),
.B(n_1734),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1745),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1760),
.B(n_1734),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1765),
.B(n_1730),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1748),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1750),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1750),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1748),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1763),
.B(n_1733),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1767),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1765),
.B(n_1730),
.Y(n_1781)
);

AOI222xp33_ASAP7_75t_L g1782 ( 
.A1(n_1752),
.A2(n_1716),
.B1(n_1739),
.B2(n_1728),
.C1(n_1616),
.C2(n_1674),
.Y(n_1782)
);

INVx2_ASAP7_75t_SL g1783 ( 
.A(n_1763),
.Y(n_1783)
);

NAND2x1p5_ASAP7_75t_L g1784 ( 
.A(n_1742),
.B(n_1337),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1744),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1759),
.B(n_1728),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1754),
.B(n_1733),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_R g1788 ( 
.A(n_1786),
.B(n_1423),
.Y(n_1788)
);

OAI21xp33_ASAP7_75t_L g1789 ( 
.A1(n_1778),
.A2(n_1743),
.B(n_1769),
.Y(n_1789)
);

AOI322xp5_ASAP7_75t_L g1790 ( 
.A1(n_1783),
.A2(n_1746),
.A3(n_1785),
.B1(n_1744),
.B2(n_1772),
.C1(n_1777),
.C2(n_1776),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1775),
.A2(n_1758),
.B1(n_1732),
.B2(n_1762),
.Y(n_1791)
);

AOI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1768),
.A2(n_1747),
.B1(n_1761),
.B2(n_1755),
.C(n_1767),
.Y(n_1792)
);

NAND3xp33_ASAP7_75t_SL g1793 ( 
.A(n_1782),
.B(n_1786),
.C(n_1784),
.Y(n_1793)
);

AOI21xp33_ASAP7_75t_SL g1794 ( 
.A1(n_1784),
.A2(n_1722),
.B(n_1749),
.Y(n_1794)
);

AOI221xp5_ASAP7_75t_L g1795 ( 
.A1(n_1783),
.A2(n_1779),
.B1(n_1787),
.B2(n_1755),
.C(n_1761),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1779),
.Y(n_1796)
);

OAI32xp33_ASAP7_75t_L g1797 ( 
.A1(n_1787),
.A2(n_1735),
.A3(n_1764),
.B1(n_1756),
.B2(n_1732),
.Y(n_1797)
);

AOI322xp5_ASAP7_75t_L g1798 ( 
.A1(n_1770),
.A2(n_1780),
.A3(n_1781),
.B1(n_1774),
.B2(n_1775),
.C1(n_1751),
.C2(n_1773),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_SL g1799 ( 
.A(n_1771),
.B(n_1735),
.C(n_1706),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1771),
.B(n_1722),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1773),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1794),
.B(n_1789),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1801),
.Y(n_1803)
);

NOR3xp33_ASAP7_75t_L g1804 ( 
.A(n_1793),
.B(n_1757),
.C(n_1723),
.Y(n_1804)
);

NAND4xp75_ASAP7_75t_L g1805 ( 
.A(n_1795),
.B(n_1706),
.C(n_1740),
.D(n_1729),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1788),
.B(n_1715),
.Y(n_1806)
);

NAND3xp33_ASAP7_75t_L g1807 ( 
.A(n_1790),
.B(n_1792),
.C(n_1798),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1796),
.Y(n_1808)
);

NOR3xp33_ASAP7_75t_L g1809 ( 
.A(n_1791),
.B(n_1757),
.C(n_1726),
.Y(n_1809)
);

NOR2x1_ASAP7_75t_L g1810 ( 
.A(n_1800),
.B(n_1423),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1799),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1797),
.Y(n_1812)
);

NAND4xp25_ASAP7_75t_L g1813 ( 
.A(n_1789),
.B(n_1740),
.C(n_1738),
.D(n_1723),
.Y(n_1813)
);

AO22x2_ASAP7_75t_L g1814 ( 
.A1(n_1796),
.A2(n_1738),
.B1(n_1737),
.B2(n_1726),
.Y(n_1814)
);

NOR3xp33_ASAP7_75t_L g1815 ( 
.A(n_1807),
.B(n_1731),
.C(n_1729),
.Y(n_1815)
);

INVxp67_ASAP7_75t_L g1816 ( 
.A(n_1802),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1806),
.B(n_1731),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1804),
.B(n_1737),
.Y(n_1818)
);

AOI211xp5_ASAP7_75t_L g1819 ( 
.A1(n_1809),
.A2(n_1370),
.B(n_1476),
.C(n_1337),
.Y(n_1819)
);

OAI221xp5_ASAP7_75t_SL g1820 ( 
.A1(n_1812),
.A2(n_1811),
.B1(n_1808),
.B2(n_1813),
.C(n_1803),
.Y(n_1820)
);

NOR2x1_ASAP7_75t_L g1821 ( 
.A(n_1818),
.B(n_1805),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1817),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1816),
.Y(n_1823)
);

AOI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1815),
.A2(n_1810),
.B1(n_1814),
.B2(n_1648),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1819),
.B(n_1370),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1820),
.B(n_1814),
.Y(n_1826)
);

NAND3xp33_ASAP7_75t_SL g1827 ( 
.A(n_1815),
.B(n_1700),
.C(n_1671),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1821),
.B(n_1631),
.Y(n_1828)
);

NOR2x1_ASAP7_75t_L g1829 ( 
.A(n_1826),
.B(n_1331),
.Y(n_1829)
);

NOR3xp33_ASAP7_75t_L g1830 ( 
.A(n_1823),
.B(n_1704),
.C(n_1700),
.Y(n_1830)
);

NOR3xp33_ASAP7_75t_L g1831 ( 
.A(n_1822),
.B(n_1704),
.C(n_1648),
.Y(n_1831)
);

INVxp33_ASAP7_75t_L g1832 ( 
.A(n_1825),
.Y(n_1832)
);

OAI211xp5_ASAP7_75t_L g1833 ( 
.A1(n_1824),
.A2(n_1331),
.B(n_1631),
.C(n_1645),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1828),
.A2(n_1827),
.B(n_1648),
.Y(n_1834)
);

BUFx3_ASAP7_75t_L g1835 ( 
.A(n_1832),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1830),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1835),
.Y(n_1837)
);

NOR3xp33_ASAP7_75t_SL g1838 ( 
.A(n_1837),
.B(n_1836),
.C(n_1834),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1838),
.B(n_1829),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1838),
.A2(n_1833),
.B(n_1831),
.Y(n_1840)
);

XNOR2xp5_ASAP7_75t_L g1841 ( 
.A(n_1839),
.B(n_1331),
.Y(n_1841)
);

OA21x2_ASAP7_75t_L g1842 ( 
.A1(n_1840),
.A2(n_1650),
.B(n_1644),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1842),
.Y(n_1843)
);

NAND3xp33_ASAP7_75t_L g1844 ( 
.A(n_1841),
.B(n_1356),
.C(n_1657),
.Y(n_1844)
);

OAI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1843),
.A2(n_1844),
.B(n_1657),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1845),
.A2(n_1645),
.B1(n_1407),
.B2(n_1631),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1846),
.A2(n_1655),
.B1(n_1602),
.B2(n_1589),
.C(n_1622),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1847),
.A2(n_1655),
.B1(n_1660),
.B2(n_1658),
.Y(n_1848)
);


endmodule