module real_jpeg_25980_n_16 (n_5, n_4, n_8, n_0, n_12, n_351, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_351;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g87 ( 
.A(n_3),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_4),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_4),
.B(n_91),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_4),
.B(n_30),
.C(n_46),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_4),
.A2(n_48),
.B1(n_49),
.B2(n_81),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_4),
.B(n_74),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_4),
.A2(n_27),
.B1(n_167),
.B2(n_170),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_5),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_5),
.A2(n_51),
.B1(n_65),
.B2(n_68),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_5),
.A2(n_51),
.B1(n_80),
.B2(n_90),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_6),
.A2(n_38),
.B1(n_48),
.B2(n_49),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_6),
.A2(n_38),
.B1(n_65),
.B2(n_68),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_6),
.A2(n_38),
.B1(n_83),
.B2(n_285),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_7),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_7),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_7),
.A2(n_67),
.B1(n_80),
.B2(n_90),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_67),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_67),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_9),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_9),
.A2(n_35),
.B1(n_65),
.B2(n_68),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_9),
.A2(n_35),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_10),
.A2(n_61),
.B1(n_65),
.B2(n_68),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_61),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_10),
.A2(n_61),
.B1(n_89),
.B2(n_90),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_11),
.A2(n_65),
.B1(n_68),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_11),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_76),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_76),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_11),
.A2(n_76),
.B1(n_89),
.B2(n_90),
.Y(n_232)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_12),
.B(n_68),
.C(n_87),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_13),
.A2(n_80),
.B1(n_83),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_13),
.A2(n_65),
.B1(n_68),
.B2(n_94),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_94),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_94),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_15),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_343),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_330),
.B(n_342),
.Y(n_17)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_293),
.A3(n_323),
.B1(n_328),
.B2(n_329),
.C(n_351),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_266),
.B(n_292),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_238),
.B(n_265),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_129),
.B(n_217),
.C(n_237),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_115),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_23),
.B(n_115),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_95),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_58),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_25),
.B(n_58),
.C(n_95),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_43),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_26),
.B(n_43),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_36),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_27),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_27),
.A2(n_40),
.B1(n_160),
.B2(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_27),
.A2(n_36),
.B(n_149),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_27),
.A2(n_149),
.B(n_174),
.Y(n_244)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_28),
.A2(n_34),
.B1(n_39),
.B2(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_28),
.B(n_37),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_28),
.A2(n_39),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_29),
.B(n_173),
.Y(n_172)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_32),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_42),
.A2(n_111),
.B(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g147 ( 
.A(n_42),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B(n_52),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_57),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_44),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_44),
.A2(n_54),
.B1(n_142),
.B2(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_44),
.B(n_81),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_44),
.A2(n_54),
.B(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_45),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_47),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_49),
.B1(n_71),
.B2(n_72),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_48),
.A2(n_72),
.B(n_183),
.C(n_185),
.Y(n_182)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_49),
.B(n_137),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_L g185 ( 
.A(n_49),
.B(n_68),
.C(n_71),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_52),
.B(n_207),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_60),
.B(n_62),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_53),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_53),
.A2(n_140),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_53),
.A2(n_140),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_54),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_54),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.C(n_77),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_63),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_60),
.B(n_140),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_60),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_62),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_63)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_68),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_65),
.A2(n_82),
.B(n_86),
.C(n_113),
.Y(n_112)
);

HAxp5_ASAP7_75t_SL g184 ( 
.A(n_65),
.B(n_81),
.CON(n_184),
.SN(n_184)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_69),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_69),
.A2(n_74),
.B1(n_127),
.B2(n_184),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_69),
.A2(n_106),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_69),
.B(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_69),
.A2(n_74),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_69),
.A2(n_234),
.B(n_273),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_69),
.A2(n_74),
.B(n_106),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_73),
.A2(n_104),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_73),
.B(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_73),
.A2(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_84),
.B1(n_91),
.B2(n_92),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B(n_82),
.Y(n_78)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_79),
.Y(n_285)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_80),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_81),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_81),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_84),
.A2(n_91),
.B1(n_101),
.B2(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_84),
.B(n_284),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_84),
.A2(n_91),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_84),
.A2(n_318),
.B(n_337),
.Y(n_336)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_93),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_85),
.A2(n_298),
.B(n_299),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_91),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_91),
.B(n_284),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_107),
.B2(n_114),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_98),
.B(n_102),
.C(n_114),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_99),
.A2(n_253),
.B(n_254),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_99),
.A2(n_282),
.B(n_283),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B(n_105),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_105),
.B(n_259),
.Y(n_315)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.C(n_120),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_116),
.B(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_118),
.B(n_120),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.C(n_125),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_121),
.A2(n_123),
.B1(n_124),
.B2(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_122),
.B(n_146),
.Y(n_223)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_125),
.B(n_200),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_216),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_211),
.B(n_215),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_195),
.B(n_210),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_178),
.B(n_194),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_156),
.B(n_177),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_143),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_143),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_138),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_150),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_144),
.B(n_151),
.C(n_154),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_163),
.B(n_176),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_162),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_168),
.B(n_175),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_166),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_193),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_193),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_188),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_189),
.C(n_190),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_186),
.B2(n_187),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_197),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_202),
.B2(n_203),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_205),
.C(n_208),
.Y(n_214)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_203)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_214),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_219),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_236),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_228),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_228),
.C(n_236),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_227),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_227),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_226),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_231),
.C(n_233),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_239),
.B(n_240),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_264),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_249),
.B1(n_262),
.B2(n_263),
.Y(n_241)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_263),
.C(n_264),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_248),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_243),
.A2(n_244),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_243),
.A2(n_277),
.B(n_281),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_245),
.Y(n_278)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_256),
.C(n_261),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_256),
.B1(n_257),
.B2(n_261),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_254),
.B(n_299),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_267),
.B(n_268),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_268)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_276),
.B1(n_287),
.B2(n_288),
.Y(n_269)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

OAI21xp33_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_274),
.B(n_275),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_274),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_275),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_275),
.A2(n_295),
.B1(n_307),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_287),
.C(n_291),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_286),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_283),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_289),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_309),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_309),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_307),
.C(n_308),
.Y(n_294)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_295),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_300),
.B2(n_301),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_297),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_302),
.C(n_306),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_312),
.C(n_322),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_298),
.Y(n_317)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_302),
.A2(n_303),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_303),
.B(n_314),
.C(n_316),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_322),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

INVx8_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_332),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_340),
.B2(n_341),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_338),
.B2(n_339),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_335),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_336),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_338),
.C(n_340),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_348),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_345),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_349),
.Y(n_348)
);


endmodule