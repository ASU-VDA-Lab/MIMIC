module real_aes_7740_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_1), .A2(n_146), .B(n_151), .C(n_188), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_2), .A2(n_141), .B(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g458 ( .A(n_3), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_4), .B(n_165), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_5), .A2(n_15), .B1(n_721), .B2(n_722), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_5), .Y(n_722) );
AOI21xp33_ASAP7_75t_L g475 ( .A1(n_6), .A2(n_141), .B(n_476), .Y(n_475) );
AND2x6_ASAP7_75t_L g146 ( .A(n_7), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g175 ( .A(n_8), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_9), .B(n_44), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_9), .B(n_44), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_10), .A2(n_253), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_11), .B(n_156), .Y(n_192) );
INVx1_ASAP7_75t_L g480 ( .A(n_12), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_13), .B(n_155), .Y(n_528) );
INVx1_ASAP7_75t_L g139 ( .A(n_14), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_15), .Y(n_721) );
INVx1_ASAP7_75t_L g540 ( .A(n_16), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_17), .A2(n_176), .B(n_201), .C(n_203), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_18), .B(n_165), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_19), .B(n_469), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_20), .B(n_141), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_21), .B(n_261), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_22), .A2(n_155), .B(n_157), .C(n_161), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_23), .B(n_165), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_24), .B(n_156), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_25), .A2(n_159), .B(n_203), .C(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_26), .B(n_156), .Y(n_237) );
CKINVDCx16_ASAP7_75t_R g221 ( .A(n_27), .Y(n_221) );
INVx1_ASAP7_75t_L g235 ( .A(n_28), .Y(n_235) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_29), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_30), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_31), .B(n_156), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_32), .A2(n_104), .B1(n_114), .B2(n_733), .Y(n_103) );
INVx1_ASAP7_75t_L g258 ( .A(n_33), .Y(n_258) );
INVx1_ASAP7_75t_L g493 ( .A(n_34), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_35), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g144 ( .A(n_36), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_37), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_38), .A2(n_155), .B(n_214), .C(n_216), .Y(n_213) );
INVxp67_ASAP7_75t_L g259 ( .A(n_39), .Y(n_259) );
CKINVDCx14_ASAP7_75t_R g212 ( .A(n_40), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_41), .A2(n_151), .B(n_234), .C(n_240), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_42), .A2(n_146), .B(n_151), .C(n_508), .Y(n_507) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_43), .A2(n_92), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_43), .Y(n_125) );
INVx1_ASAP7_75t_L g492 ( .A(n_45), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_46), .A2(n_173), .B(n_174), .C(n_177), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_47), .B(n_156), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_48), .A2(n_122), .B1(n_434), .B2(n_435), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_48), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_49), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_50), .Y(n_255) );
INVx1_ASAP7_75t_L g149 ( .A(n_51), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_52), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_53), .B(n_141), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_54), .A2(n_151), .B1(n_161), .B2(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_55), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g455 ( .A(n_56), .Y(n_455) );
CKINVDCx14_ASAP7_75t_R g171 ( .A(n_57), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_58), .A2(n_173), .B(n_216), .C(n_479), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_59), .Y(n_521) );
INVx1_ASAP7_75t_L g477 ( .A(n_60), .Y(n_477) );
INVx1_ASAP7_75t_L g147 ( .A(n_61), .Y(n_147) );
INVx1_ASAP7_75t_L g138 ( .A(n_62), .Y(n_138) );
INVx1_ASAP7_75t_SL g215 ( .A(n_63), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_64), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_65), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g224 ( .A(n_66), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_SL g468 ( .A1(n_67), .A2(n_216), .B(n_469), .C(n_470), .Y(n_468) );
INVxp67_ASAP7_75t_L g471 ( .A(n_68), .Y(n_471) );
INVx1_ASAP7_75t_L g113 ( .A(n_69), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_70), .A2(n_141), .B(n_170), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_71), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_72), .A2(n_141), .B(n_198), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_73), .Y(n_496) );
INVx1_ASAP7_75t_L g515 ( .A(n_74), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_75), .A2(n_253), .B(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g199 ( .A(n_76), .Y(n_199) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_77), .Y(n_232) );
AOI222xp33_ASAP7_75t_L g445 ( .A1(n_78), .A2(n_446), .B1(n_718), .B2(n_724), .C1(n_728), .C2(n_729), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_79), .A2(n_146), .B(n_151), .C(n_517), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_80), .A2(n_141), .B(n_148), .Y(n_140) );
INVx1_ASAP7_75t_L g202 ( .A(n_81), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_82), .B(n_236), .Y(n_509) );
INVx2_ASAP7_75t_L g136 ( .A(n_83), .Y(n_136) );
INVx1_ASAP7_75t_L g189 ( .A(n_84), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_85), .B(n_469), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_86), .A2(n_146), .B(n_151), .C(n_457), .Y(n_456) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_87), .B(n_110), .C(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g438 ( .A(n_87), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g716 ( .A(n_87), .Y(n_716) );
OR2x2_ASAP7_75t_L g717 ( .A(n_87), .B(n_440), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_88), .A2(n_151), .B(n_223), .C(n_226), .Y(n_222) );
OAI22xp5_ASAP7_75t_SL g718 ( .A1(n_89), .A2(n_719), .B1(n_720), .B2(n_723), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_89), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_90), .B(n_168), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_91), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_92), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_93), .A2(n_146), .B(n_151), .C(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_94), .Y(n_532) );
INVx1_ASAP7_75t_L g467 ( .A(n_95), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_96), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_97), .B(n_236), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_98), .B(n_134), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_99), .B(n_134), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_100), .B(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g158 ( .A(n_101), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_102), .A2(n_141), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g733 ( .A(n_106), .Y(n_733) );
CKINVDCx12_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x2_ASAP7_75t_L g440 ( .A(n_110), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AO21x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_444), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g732 ( .A(n_117), .Y(n_732) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_436), .B(n_442), .Y(n_120) );
INVx1_ASAP7_75t_L g435 ( .A(n_122), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_126), .B1(n_432), .B2(n_433), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_123), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_126), .A2(n_715), .B1(n_725), .B2(n_726), .Y(n_724) );
BUFx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g433 ( .A(n_127), .Y(n_433) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_358), .Y(n_127) );
NOR4xp25_ASAP7_75t_L g128 ( .A(n_129), .B(n_300), .C(n_330), .D(n_340), .Y(n_128) );
OAI211xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_205), .B(n_263), .C(n_290), .Y(n_129) );
OAI222xp33_ASAP7_75t_L g385 ( .A1(n_130), .A2(n_305), .B1(n_386), .B2(n_387), .C1(n_388), .C2(n_389), .Y(n_385) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_180), .Y(n_130) );
AOI33xp33_ASAP7_75t_L g311 ( .A1(n_131), .A2(n_298), .A3(n_299), .B1(n_312), .B2(n_317), .B3(n_319), .Y(n_311) );
OAI211xp5_ASAP7_75t_SL g368 ( .A1(n_131), .A2(n_369), .B(n_371), .C(n_373), .Y(n_368) );
OR2x2_ASAP7_75t_L g384 ( .A(n_131), .B(n_370), .Y(n_384) );
INVx1_ASAP7_75t_L g417 ( .A(n_131), .Y(n_417) );
OR2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_167), .Y(n_131) );
INVx2_ASAP7_75t_L g294 ( .A(n_132), .Y(n_294) );
AND2x2_ASAP7_75t_L g310 ( .A(n_132), .B(n_196), .Y(n_310) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_132), .Y(n_345) );
AND2x2_ASAP7_75t_L g374 ( .A(n_132), .B(n_167), .Y(n_374) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_140), .B(n_164), .Y(n_132) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_133), .A2(n_197), .B(n_204), .Y(n_196) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_133), .A2(n_210), .B(n_218), .Y(n_209) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx4_ASAP7_75t_L g166 ( .A(n_134), .Y(n_166) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_134), .A2(n_465), .B(n_472), .Y(n_464) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g251 ( .A(n_135), .Y(n_251) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g168 ( .A(n_136), .B(n_137), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx2_ASAP7_75t_L g253 ( .A(n_141), .Y(n_253) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_142), .B(n_146), .Y(n_186) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx1_ASAP7_75t_L g239 ( .A(n_143), .Y(n_239) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
INVx1_ASAP7_75t_L g162 ( .A(n_144), .Y(n_162) );
INVx1_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_145), .Y(n_160) );
INVx3_ASAP7_75t_L g176 ( .A(n_145), .Y(n_176) );
INVx1_ASAP7_75t_L g469 ( .A(n_145), .Y(n_469) );
INVx4_ASAP7_75t_SL g163 ( .A(n_146), .Y(n_163) );
BUFx3_ASAP7_75t_L g240 ( .A(n_146), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g148 ( .A1(n_149), .A2(n_150), .B(n_154), .C(n_163), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_SL g170 ( .A1(n_150), .A2(n_163), .B(n_171), .C(n_172), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_SL g198 ( .A1(n_150), .A2(n_163), .B(n_199), .C(n_200), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_150), .A2(n_163), .B(n_212), .C(n_213), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_SL g254 ( .A1(n_150), .A2(n_163), .B(n_255), .C(n_256), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_150), .A2(n_163), .B(n_467), .C(n_468), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_150), .A2(n_163), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_150), .A2(n_163), .B(n_537), .C(n_538), .Y(n_536) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx3_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_152), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_155), .B(n_215), .Y(n_214) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g173 ( .A(n_156), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_159), .B(n_202), .Y(n_201) );
OAI22xp33_ASAP7_75t_L g257 ( .A1(n_159), .A2(n_236), .B1(n_258), .B2(n_259), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_159), .B(n_540), .Y(n_539) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g191 ( .A(n_160), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g491 ( .A1(n_160), .A2(n_191), .B1(n_492), .B2(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g460 ( .A(n_161), .Y(n_460) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g226 ( .A(n_163), .Y(n_226) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_163), .A2(n_186), .B1(n_490), .B2(n_494), .Y(n_489) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_165), .A2(n_475), .B(n_481), .Y(n_474) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_166), .B(n_195), .Y(n_194) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_166), .A2(n_220), .B(n_227), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_166), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_SL g511 ( .A(n_166), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g274 ( .A(n_167), .Y(n_274) );
BUFx3_ASAP7_75t_L g282 ( .A(n_167), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_167), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g293 ( .A(n_167), .B(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_167), .B(n_181), .Y(n_322) );
AND2x2_ASAP7_75t_L g391 ( .A(n_167), .B(n_325), .Y(n_391) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_179), .Y(n_167) );
INVx1_ASAP7_75t_L g183 ( .A(n_168), .Y(n_183) );
INVx2_ASAP7_75t_L g229 ( .A(n_168), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_168), .A2(n_186), .B(n_232), .C(n_233), .Y(n_231) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_168), .A2(n_535), .B(n_541), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
INVx5_ASAP7_75t_L g236 ( .A(n_176), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_176), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_176), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g193 ( .A(n_177), .Y(n_193) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g203 ( .A(n_178), .Y(n_203) );
INVx2_ASAP7_75t_SL g285 ( .A(n_180), .Y(n_285) );
OR2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_196), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_181), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g327 ( .A(n_181), .Y(n_327) );
AND2x2_ASAP7_75t_L g338 ( .A(n_181), .B(n_294), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_181), .B(n_323), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_181), .B(n_325), .Y(n_370) );
AND2x2_ASAP7_75t_L g429 ( .A(n_181), .B(n_374), .Y(n_429) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g299 ( .A(n_182), .B(n_196), .Y(n_299) );
AND2x2_ASAP7_75t_L g309 ( .A(n_182), .B(n_310), .Y(n_309) );
BUFx3_ASAP7_75t_L g331 ( .A(n_182), .Y(n_331) );
AND3x2_ASAP7_75t_L g390 ( .A(n_182), .B(n_391), .C(n_392), .Y(n_390) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_194), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_183), .B(n_462), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_183), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_183), .B(n_532), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_186), .A2(n_221), .B(n_222), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_186), .A2(n_455), .B(n_456), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_186), .A2(n_515), .B(n_516), .Y(n_514) );
O2A1O1Ixp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_192), .C(n_193), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_190), .A2(n_193), .B(n_224), .C(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_193), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_193), .A2(n_518), .B(n_519), .Y(n_517) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_196), .Y(n_281) );
INVx1_ASAP7_75t_SL g325 ( .A(n_196), .Y(n_325) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_196), .B(n_274), .C(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_243), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g360 ( .A1(n_206), .A2(n_309), .B(n_361), .C(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_208), .B(n_230), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_208), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_SL g377 ( .A(n_208), .Y(n_377) );
AND2x2_ASAP7_75t_L g398 ( .A(n_208), .B(n_245), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_208), .B(n_307), .Y(n_426) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_219), .Y(n_208) );
AND2x2_ASAP7_75t_L g271 ( .A(n_209), .B(n_262), .Y(n_271) );
INVx2_ASAP7_75t_L g278 ( .A(n_209), .Y(n_278) );
AND2x2_ASAP7_75t_L g298 ( .A(n_209), .B(n_245), .Y(n_298) );
AND2x2_ASAP7_75t_L g348 ( .A(n_209), .B(n_230), .Y(n_348) );
INVx1_ASAP7_75t_L g352 ( .A(n_209), .Y(n_352) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_217), .Y(n_529) );
INVx2_ASAP7_75t_SL g262 ( .A(n_219), .Y(n_262) );
BUFx2_ASAP7_75t_L g288 ( .A(n_219), .Y(n_288) );
AND2x2_ASAP7_75t_L g415 ( .A(n_219), .B(n_230), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g261 ( .A(n_229), .Y(n_261) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_229), .A2(n_524), .B(n_531), .Y(n_523) );
INVx3_ASAP7_75t_SL g245 ( .A(n_230), .Y(n_245) );
AND2x2_ASAP7_75t_L g270 ( .A(n_230), .B(n_271), .Y(n_270) );
AND2x4_ASAP7_75t_L g277 ( .A(n_230), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g307 ( .A(n_230), .B(n_267), .Y(n_307) );
OR2x2_ASAP7_75t_L g316 ( .A(n_230), .B(n_262), .Y(n_316) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_230), .Y(n_334) );
AND2x2_ASAP7_75t_L g339 ( .A(n_230), .B(n_292), .Y(n_339) );
AND2x2_ASAP7_75t_L g367 ( .A(n_230), .B(n_247), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_230), .B(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g405 ( .A(n_230), .B(n_246), .Y(n_405) );
OR2x6_ASAP7_75t_L g230 ( .A(n_231), .B(n_241), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_237), .C(n_238), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_236), .A2(n_458), .B(n_459), .C(n_460), .Y(n_457) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_239), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
AND2x2_ASAP7_75t_L g329 ( .A(n_245), .B(n_278), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_245), .B(n_271), .Y(n_357) );
AND2x2_ASAP7_75t_L g375 ( .A(n_245), .B(n_292), .Y(n_375) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_262), .Y(n_246) );
AND2x2_ASAP7_75t_L g276 ( .A(n_247), .B(n_262), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_247), .B(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g314 ( .A(n_247), .Y(n_314) );
OR2x2_ASAP7_75t_L g362 ( .A(n_247), .B(n_282), .Y(n_362) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_252), .B(n_260), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_249), .A2(n_268), .B(n_269), .Y(n_267) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_249), .A2(n_514), .B(n_520), .Y(n_513) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AOI21xp5_ASAP7_75t_SL g505 ( .A1(n_250), .A2(n_506), .B(n_507), .Y(n_505) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_251), .A2(n_454), .B(n_461), .Y(n_453) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_251), .A2(n_489), .B(n_495), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_251), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g268 ( .A(n_252), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_260), .Y(n_269) );
AND2x2_ASAP7_75t_L g297 ( .A(n_262), .B(n_267), .Y(n_297) );
INVx1_ASAP7_75t_L g305 ( .A(n_262), .Y(n_305) );
AND2x2_ASAP7_75t_L g400 ( .A(n_262), .B(n_278), .Y(n_400) );
AOI222xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_272), .B1(n_275), .B2(n_279), .C1(n_283), .C2(n_286), .Y(n_263) );
INVx1_ASAP7_75t_L g395 ( .A(n_264), .Y(n_395) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_270), .Y(n_264) );
AND2x2_ASAP7_75t_L g291 ( .A(n_265), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g302 ( .A(n_265), .B(n_271), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_265), .B(n_293), .Y(n_318) );
OAI222xp33_ASAP7_75t_L g340 ( .A1(n_265), .A2(n_341), .B1(n_346), .B2(n_347), .C1(n_355), .C2(n_357), .Y(n_340) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g328 ( .A(n_267), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_267), .B(n_348), .Y(n_388) );
AND2x2_ASAP7_75t_L g399 ( .A(n_267), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g407 ( .A(n_270), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_272), .B(n_323), .Y(n_386) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_274), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g344 ( .A(n_274), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx3_ASAP7_75t_L g289 ( .A(n_277), .Y(n_289) );
O2A1O1Ixp33_ASAP7_75t_L g379 ( .A1(n_277), .A2(n_380), .B(n_383), .C(n_385), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_277), .B(n_314), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_277), .B(n_297), .Y(n_419) );
AND2x2_ASAP7_75t_L g292 ( .A(n_278), .B(n_288), .Y(n_292) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g319 ( .A(n_281), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_282), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g371 ( .A(n_282), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g410 ( .A(n_282), .B(n_310), .Y(n_410) );
INVx1_ASAP7_75t_L g422 ( .A(n_282), .Y(n_422) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_285), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g403 ( .A(n_288), .Y(n_403) );
A2O1A1Ixp33_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_293), .B(n_295), .C(n_299), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_291), .A2(n_321), .B1(n_336), .B2(n_339), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_292), .B(n_306), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_292), .B(n_314), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_293), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g356 ( .A(n_293), .Y(n_356) );
AND2x2_ASAP7_75t_L g363 ( .A(n_293), .B(n_343), .Y(n_363) );
INVx2_ASAP7_75t_L g324 ( .A(n_294), .Y(n_324) );
INVxp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NOR4xp25_ASAP7_75t_L g301 ( .A(n_298), .B(n_302), .C(n_303), .D(n_306), .Y(n_301) );
INVx1_ASAP7_75t_SL g372 ( .A(n_299), .Y(n_372) );
AND2x2_ASAP7_75t_L g416 ( .A(n_299), .B(n_417), .Y(n_416) );
OAI211xp5_ASAP7_75t_SL g300 ( .A1(n_301), .A2(n_308), .B(n_311), .C(n_320), .Y(n_300) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_307), .B(n_377), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_309), .A2(n_428), .B1(n_429), .B2(n_430), .Y(n_427) );
INVx1_ASAP7_75t_SL g382 ( .A(n_310), .Y(n_382) );
AND2x2_ASAP7_75t_L g421 ( .A(n_310), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_314), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_318), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_319), .B(n_344), .Y(n_404) );
OAI21xp5_ASAP7_75t_SL g320 ( .A1(n_321), .A2(n_326), .B(n_328), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g396 ( .A(n_323), .Y(n_396) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx2_ASAP7_75t_L g424 ( .A(n_324), .Y(n_424) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_325), .Y(n_351) );
OAI21xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B(n_335), .Y(n_330) );
CKINVDCx16_ASAP7_75t_R g343 ( .A(n_331), .Y(n_343) );
OR2x2_ASAP7_75t_L g381 ( .A(n_331), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI21xp33_ASAP7_75t_SL g376 ( .A1(n_334), .A2(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_338), .A2(n_365), .B1(n_368), .B2(n_375), .C(n_376), .Y(n_364) );
INVx1_ASAP7_75t_SL g408 ( .A(n_339), .Y(n_408) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
OR2x2_ASAP7_75t_L g355 ( .A(n_343), .B(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g392 ( .A(n_345), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_352), .B2(n_353), .Y(n_347) );
INVx1_ASAP7_75t_L g387 ( .A(n_348), .Y(n_387) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_351), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR4xp25_ASAP7_75t_L g358 ( .A(n_359), .B(n_393), .C(n_406), .D(n_418), .Y(n_358) );
NAND3xp33_ASAP7_75t_SL g359 ( .A(n_360), .B(n_364), .C(n_379), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_362), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_369), .B(n_374), .Y(n_378) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI221xp5_ASAP7_75t_SL g406 ( .A1(n_381), .A2(n_407), .B1(n_408), .B2(n_409), .C(n_411), .Y(n_406) );
O2A1O1Ixp33_ASAP7_75t_L g397 ( .A1(n_383), .A2(n_398), .B(n_399), .C(n_401), .Y(n_397) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_384), .A2(n_402), .B1(n_404), .B2(n_405), .Y(n_401) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
A2O1A1Ixp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B(n_396), .C(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g412 ( .A(n_405), .Y(n_412) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI21xp5_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_413), .B(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g418 ( .A1(n_419), .A2(n_420), .B1(n_423), .B2(n_425), .C(n_427), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_433), .A2(n_447), .B1(n_715), .B2(n_717), .Y(n_446) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g443 ( .A(n_438), .Y(n_443) );
NOR2x2_ASAP7_75t_L g731 ( .A(n_439), .B(n_716), .Y(n_731) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g715 ( .A(n_440), .B(n_716), .Y(n_715) );
AOI21xp33_ASAP7_75t_SL g444 ( .A1(n_442), .A2(n_445), .B(n_732), .Y(n_444) );
INVx1_ASAP7_75t_L g725 ( .A(n_447), .Y(n_725) );
NAND2x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_631), .Y(n_447) );
NOR5xp2_ASAP7_75t_L g448 ( .A(n_449), .B(n_554), .C(n_586), .D(n_601), .E(n_618), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_482), .B(n_501), .C(n_542), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_463), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_451), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_451), .B(n_606), .Y(n_669) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_452), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_452), .B(n_498), .Y(n_555) );
AND2x2_ASAP7_75t_L g596 ( .A(n_452), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_452), .B(n_565), .Y(n_600) );
OR2x2_ASAP7_75t_L g637 ( .A(n_452), .B(n_488), .Y(n_637) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g487 ( .A(n_453), .B(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g545 ( .A(n_453), .Y(n_545) );
OR2x2_ASAP7_75t_L g708 ( .A(n_453), .B(n_548), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_463), .A2(n_611), .B1(n_612), .B2(n_615), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_463), .B(n_545), .Y(n_694) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_473), .Y(n_463) );
AND2x2_ASAP7_75t_L g500 ( .A(n_464), .B(n_488), .Y(n_500) );
AND2x2_ASAP7_75t_L g547 ( .A(n_464), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g552 ( .A(n_464), .Y(n_552) );
INVx3_ASAP7_75t_L g565 ( .A(n_464), .Y(n_565) );
OR2x2_ASAP7_75t_L g585 ( .A(n_464), .B(n_548), .Y(n_585) );
AND2x2_ASAP7_75t_L g604 ( .A(n_464), .B(n_474), .Y(n_604) );
BUFx2_ASAP7_75t_L g636 ( .A(n_464), .Y(n_636) );
AND2x4_ASAP7_75t_L g551 ( .A(n_473), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g486 ( .A(n_474), .Y(n_486) );
INVx2_ASAP7_75t_L g499 ( .A(n_474), .Y(n_499) );
OR2x2_ASAP7_75t_L g567 ( .A(n_474), .B(n_548), .Y(n_567) );
AND2x2_ASAP7_75t_L g597 ( .A(n_474), .B(n_488), .Y(n_597) );
AND2x2_ASAP7_75t_L g614 ( .A(n_474), .B(n_545), .Y(n_614) );
AND2x2_ASAP7_75t_L g654 ( .A(n_474), .B(n_565), .Y(n_654) );
AND2x2_ASAP7_75t_SL g690 ( .A(n_474), .B(n_500), .Y(n_690) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp33_ASAP7_75t_SL g483 ( .A(n_484), .B(n_497), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_485), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
OAI21xp33_ASAP7_75t_L g628 ( .A1(n_486), .A2(n_500), .B(n_629), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_486), .B(n_488), .Y(n_684) );
AND2x2_ASAP7_75t_L g620 ( .A(n_487), .B(n_621), .Y(n_620) );
INVx3_ASAP7_75t_L g548 ( .A(n_488), .Y(n_548) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_488), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_497), .B(n_545), .Y(n_713) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_498), .A2(n_656), .B1(n_657), .B2(n_662), .Y(n_655) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
AND2x2_ASAP7_75t_L g546 ( .A(n_499), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g584 ( .A(n_499), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_SL g621 ( .A(n_499), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_500), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g675 ( .A(n_500), .Y(n_675) );
CKINVDCx16_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_522), .Y(n_502) );
INVx4_ASAP7_75t_L g561 ( .A(n_503), .Y(n_561) );
AND2x2_ASAP7_75t_L g639 ( .A(n_503), .B(n_606), .Y(n_639) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_513), .Y(n_503) );
INVx3_ASAP7_75t_L g558 ( .A(n_504), .Y(n_558) );
AND2x2_ASAP7_75t_L g572 ( .A(n_504), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g576 ( .A(n_504), .Y(n_576) );
INVx2_ASAP7_75t_L g590 ( .A(n_504), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_504), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g647 ( .A(n_504), .B(n_642), .Y(n_647) );
AND2x2_ASAP7_75t_L g712 ( .A(n_504), .B(n_682), .Y(n_712) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_511), .Y(n_504) );
AND2x2_ASAP7_75t_L g553 ( .A(n_513), .B(n_534), .Y(n_553) );
INVx2_ASAP7_75t_L g573 ( .A(n_513), .Y(n_573) );
INVx1_ASAP7_75t_L g578 ( .A(n_522), .Y(n_578) );
AND2x2_ASAP7_75t_L g624 ( .A(n_522), .B(n_572), .Y(n_624) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_533), .Y(n_522) );
INVx2_ASAP7_75t_L g563 ( .A(n_523), .Y(n_563) );
INVx1_ASAP7_75t_L g571 ( .A(n_523), .Y(n_571) );
AND2x2_ASAP7_75t_L g589 ( .A(n_523), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_523), .B(n_573), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_530), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_529), .Y(n_526) );
AND2x2_ASAP7_75t_L g606 ( .A(n_533), .B(n_563), .Y(n_606) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g559 ( .A(n_534), .Y(n_559) );
AND2x2_ASAP7_75t_L g642 ( .A(n_534), .B(n_573), .Y(n_642) );
OAI21xp5_ASAP7_75t_SL g542 ( .A1(n_543), .A2(n_549), .B(n_553), .Y(n_542) );
INVx1_ASAP7_75t_SL g587 ( .A(n_543), .Y(n_587) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_544), .B(n_551), .Y(n_644) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g593 ( .A(n_545), .B(n_548), .Y(n_593) );
AND2x2_ASAP7_75t_L g622 ( .A(n_545), .B(n_566), .Y(n_622) );
OR2x2_ASAP7_75t_L g625 ( .A(n_545), .B(n_585), .Y(n_625) );
AOI222xp33_ASAP7_75t_L g689 ( .A1(n_546), .A2(n_638), .B1(n_690), .B2(n_691), .C1(n_693), .C2(n_695), .Y(n_689) );
BUFx2_ASAP7_75t_L g603 ( .A(n_548), .Y(n_603) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g592 ( .A(n_551), .B(n_593), .Y(n_592) );
INVx3_ASAP7_75t_SL g609 ( .A(n_551), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_551), .B(n_603), .Y(n_663) );
AND2x2_ASAP7_75t_L g598 ( .A(n_553), .B(n_558), .Y(n_598) );
INVx1_ASAP7_75t_L g617 ( .A(n_553), .Y(n_617) );
OAI221xp5_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_556), .B1(n_560), .B2(n_564), .C(n_568), .Y(n_554) );
OR2x2_ASAP7_75t_L g626 ( .A(n_556), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AND2x2_ASAP7_75t_L g611 ( .A(n_558), .B(n_581), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_558), .B(n_571), .Y(n_651) );
AND2x2_ASAP7_75t_L g656 ( .A(n_558), .B(n_606), .Y(n_656) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_558), .Y(n_666) );
NAND2x1_ASAP7_75t_SL g677 ( .A(n_558), .B(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g562 ( .A(n_559), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g582 ( .A(n_559), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_559), .B(n_577), .Y(n_608) );
INVx1_ASAP7_75t_L g674 ( .A(n_559), .Y(n_674) );
INVx1_ASAP7_75t_L g649 ( .A(n_560), .Y(n_649) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g661 ( .A(n_561), .Y(n_661) );
NOR2xp67_ASAP7_75t_L g673 ( .A(n_561), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g678 ( .A(n_562), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_562), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g581 ( .A(n_563), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_563), .B(n_573), .Y(n_594) );
INVx1_ASAP7_75t_L g660 ( .A(n_563), .Y(n_660) );
INVx1_ASAP7_75t_L g681 ( .A(n_564), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI21xp5_ASAP7_75t_SL g568 ( .A1(n_569), .A2(n_574), .B(n_583), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
AND2x2_ASAP7_75t_L g714 ( .A(n_570), .B(n_647), .Y(n_714) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g682 ( .A(n_571), .B(n_642), .Y(n_682) );
AOI32xp33_ASAP7_75t_L g595 ( .A1(n_572), .A2(n_578), .A3(n_596), .B1(n_598), .B2(n_599), .Y(n_595) );
AOI322xp5_ASAP7_75t_L g697 ( .A1(n_572), .A2(n_604), .A3(n_687), .B1(n_698), .B2(n_699), .C1(n_700), .C2(n_702), .Y(n_697) );
INVx2_ASAP7_75t_L g577 ( .A(n_573), .Y(n_577) );
INVx1_ASAP7_75t_L g687 ( .A(n_573), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_578), .B1(n_579), .B2(n_580), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_575), .B(n_581), .Y(n_630) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_576), .B(n_642), .Y(n_692) );
INVx1_ASAP7_75t_L g579 ( .A(n_577), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_577), .B(n_606), .Y(n_696) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_585), .B(n_680), .Y(n_679) );
OAI221xp5_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_588), .B1(n_591), .B2(n_594), .C(n_595), .Y(n_586) );
OR2x2_ASAP7_75t_L g607 ( .A(n_588), .B(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g616 ( .A(n_588), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g641 ( .A(n_589), .B(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g645 ( .A(n_599), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OAI221xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_605), .B1(n_607), .B2(n_609), .C(n_610), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_603), .A2(n_634), .B1(n_638), .B2(n_639), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_604), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g709 ( .A(n_604), .Y(n_709) );
INVx1_ASAP7_75t_L g703 ( .A(n_606), .Y(n_703) );
INVx1_ASAP7_75t_SL g638 ( .A(n_607), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_609), .B(n_637), .Y(n_699) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_614), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g680 ( .A(n_614), .Y(n_680) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
OAI221xp5_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_623), .B1(n_625), .B2(n_626), .C(n_628), .Y(n_618) );
NOR2xp33_ASAP7_75t_SL g619 ( .A(n_620), .B(n_622), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_620), .A2(n_638), .B1(n_684), .B2(n_685), .Y(n_683) );
CKINVDCx14_ASAP7_75t_R g623 ( .A(n_624), .Y(n_623) );
OAI21xp33_ASAP7_75t_L g702 ( .A1(n_625), .A2(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NOR3xp33_ASAP7_75t_SL g631 ( .A(n_632), .B(n_664), .C(n_688), .Y(n_631) );
NAND4xp25_ASAP7_75t_L g632 ( .A(n_633), .B(n_640), .C(n_648), .D(n_655), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g711 ( .A(n_636), .Y(n_711) );
INVx3_ASAP7_75t_SL g705 ( .A(n_637), .Y(n_705) );
OR2x2_ASAP7_75t_L g710 ( .A(n_637), .B(n_711), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B1(n_645), .B2(n_647), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_642), .B(n_660), .Y(n_701) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI21xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_650), .B(n_652), .Y(n_648) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI211xp5_ASAP7_75t_SL g664 ( .A1(n_665), .A2(n_667), .B(n_670), .C(n_683), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g698 ( .A(n_669), .Y(n_698) );
AOI222xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_675), .B1(n_676), .B2(n_679), .C1(n_681), .C2(n_682), .Y(n_670) );
INVxp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND4xp25_ASAP7_75t_SL g707 ( .A(n_680), .B(n_708), .C(n_709), .D(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND3xp33_ASAP7_75t_SL g688 ( .A(n_689), .B(n_697), .C(n_706), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_706) );
INVx1_ASAP7_75t_L g727 ( .A(n_717), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_718), .Y(n_728) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
endmodule