module fake_jpeg_14111_n_238 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_6),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_51),
.Y(n_88)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_60),
.Y(n_92)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_66),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_12),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_73),
.Y(n_77)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_14),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_76),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_41),
.Y(n_94)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_30),
.B1(n_42),
.B2(n_31),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_79),
.A2(n_90),
.B1(n_115),
.B2(n_0),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_46),
.A2(n_30),
.B1(n_42),
.B2(n_23),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_94),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_53),
.A2(n_41),
.B1(n_23),
.B2(n_27),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_96),
.A2(n_114),
.B1(n_117),
.B2(n_119),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_50),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_103),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_69),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_27),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_0),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_25),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_108),
.B(n_112),
.Y(n_136)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

BUFx2_ASAP7_75t_SL g135 ( 
.A(n_109),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_35),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_49),
.A2(n_35),
.B1(n_38),
.B2(n_37),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_54),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_56),
.A2(n_67),
.B1(n_55),
.B2(n_48),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_62),
.A2(n_39),
.B1(n_3),
.B2(n_4),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_121),
.B(n_134),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_107),
.B(n_85),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_125),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_14),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_3),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_4),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_139),
.Y(n_164)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_143),
.Y(n_149)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_141),
.A2(n_86),
.B1(n_99),
.B2(n_93),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_83),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_148),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_88),
.B(n_92),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_92),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_146),
.Y(n_154)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_96),
.B1(n_117),
.B2(n_111),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_133),
.B1(n_127),
.B2(n_125),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_116),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_150),
.A2(n_152),
.B1(n_100),
.B2(n_138),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_145),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_91),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_158),
.B(n_162),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_109),
.B(n_110),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_160),
.B(n_148),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_81),
.Y(n_162)
);

NAND2x1_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_86),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_84),
.C(n_146),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_159),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_170),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_148),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_181),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_176),
.A2(n_149),
.B(n_157),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_167),
.A2(n_122),
.B(n_132),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_170),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_139),
.C(n_120),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_180),
.C(n_161),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_136),
.B1(n_140),
.B2(n_87),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_182),
.B1(n_166),
.B2(n_172),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_129),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_130),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_128),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_183),
.B(n_184),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_156),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_156),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_187),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_189),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_150),
.B1(n_164),
.B2(n_165),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_177),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_196),
.C(n_180),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_164),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_168),
.A2(n_150),
.B1(n_161),
.B2(n_163),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_181),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_203),
.A2(n_198),
.B1(n_195),
.B2(n_193),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_186),
.A2(n_169),
.B(n_179),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_205),
.B(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

AOI22x1_ASAP7_75t_SL g210 ( 
.A1(n_186),
.A2(n_171),
.B1(n_174),
.B2(n_163),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_199),
.B1(n_190),
.B2(n_194),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_198),
.B(n_208),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_216),
.Y(n_222)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_203),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_201),
.C(n_200),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_220),
.C(n_223),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_200),
.C(n_191),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_218),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_204),
.C(n_209),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_210),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_209),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_226),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_213),
.Y(n_231)
);

NOR2xp67_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_231),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_222),
.C(n_225),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_212),
.Y(n_234)
);

AOI221xp5_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_235),
.B1(n_161),
.B2(n_141),
.C(n_124),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_217),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_106),
.Y(n_237)
);

NOR2xp67_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_135),
.Y(n_238)
);


endmodule