module fake_jpeg_1547_n_40 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_40);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_3),
.B(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_17),
.B(n_15),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_19),
.B(n_20),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_12),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_14),
.B1(n_13),
.B2(n_16),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_16),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_13),
.C(n_11),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_6),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_2),
.B(n_4),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_32),
.B(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_29),
.B(n_8),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_29),
.B(n_8),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_37),
.B1(n_9),
.B2(n_10),
.Y(n_39)
);

BUFx24_ASAP7_75t_SL g40 ( 
.A(n_39),
.Y(n_40)
);


endmodule