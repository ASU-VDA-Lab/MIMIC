module fake_jpeg_28435_n_158 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_158);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_45),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_5),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_47),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_20),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_24),
.Y(n_49)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_64),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_19),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_16),
.B1(n_18),
.B2(n_26),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_68),
.B1(n_29),
.B2(n_19),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_34),
.B1(n_27),
.B2(n_15),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_67),
.Y(n_74)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_30),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_16),
.B1(n_18),
.B2(n_27),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_69),
.B(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_14),
.Y(n_81)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NAND2x1_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_49),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_85),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_22),
.C(n_27),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_80),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_59),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_22),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_56),
.Y(n_84)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_17),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_8),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_89),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_24),
.B1(n_21),
.B2(n_2),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_91),
.B1(n_59),
.B2(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_7),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_53),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_101),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_61),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_9),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_9),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_102),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_72),
.C(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_93),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_116),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_80),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_88),
.B1(n_77),
.B2(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_107),
.B1(n_113),
.B2(n_13),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_106),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_129),
.B(n_130),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_127),
.B(n_128),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_81),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_132),
.A2(n_82),
.B1(n_115),
.B2(n_113),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_116),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_140),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_138),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_98),
.C(n_92),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_125),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_98),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_134),
.Y(n_149)
);

AOI322xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_129),
.A3(n_131),
.B1(n_100),
.B2(n_92),
.C1(n_85),
.C2(n_57),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_140),
.B1(n_136),
.B2(n_78),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_50),
.C(n_11),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_147),
.A2(n_145),
.B1(n_78),
.B2(n_71),
.Y(n_153)
);

OAI21x1_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_145),
.B(n_87),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_148),
.A2(n_136),
.B(n_141),
.C(n_146),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_151),
.A2(n_152),
.A3(n_153),
.B1(n_150),
.B2(n_149),
.C1(n_50),
.C2(n_57),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_11),
.A3(n_50),
.B1(n_4),
.B2(n_58),
.C1(n_63),
.C2(n_55),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_155),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_58),
.Y(n_158)
);


endmodule