module fake_jpeg_1423_n_432 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_432);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_432;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

AOI21xp33_ASAP7_75t_SL g38 ( 
.A1(n_15),
.A2(n_8),
.B(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_49),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_46),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_47),
.Y(n_140)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_50),
.Y(n_141)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_18),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_51),
.Y(n_114)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_14),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_65),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_23),
.Y(n_54)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_27),
.B(n_13),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_38),
.B(n_30),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_81),
.Y(n_122)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_27),
.B(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_83),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_29),
.B(n_13),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_86),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_43),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_26),
.B1(n_36),
.B2(n_42),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_90),
.A2(n_97),
.B1(n_81),
.B2(n_80),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_43),
.B1(n_37),
.B2(n_42),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_94),
.A2(n_115),
.B1(n_119),
.B2(n_142),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_42),
.B1(n_37),
.B2(n_39),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_111),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_33),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_55),
.A2(n_42),
.B1(n_39),
.B2(n_31),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_46),
.B(n_33),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_131),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_86),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_120),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_59),
.A2(n_39),
.B1(n_35),
.B2(n_31),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_35),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_52),
.B(n_38),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_0),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_64),
.B(n_40),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_57),
.B(n_28),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_132),
.B(n_139),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_74),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_138),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_84),
.A2(n_40),
.B1(n_32),
.B2(n_28),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_44),
.B1(n_2),
.B2(n_3),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_32),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_85),
.B(n_25),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_25),
.B1(n_78),
.B2(n_82),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_143),
.A2(n_185),
.B1(n_113),
.B2(n_141),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_0),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_147),
.B(n_168),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_148),
.B(n_151),
.Y(n_211)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_150),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_114),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_153),
.A2(n_190),
.B1(n_106),
.B2(n_121),
.Y(n_204)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_154),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_77),
.B1(n_44),
.B2(n_14),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_158),
.B1(n_161),
.B2(n_166),
.Y(n_199)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_156),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_157),
.A2(n_162),
.B(n_173),
.Y(n_237)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_97),
.A2(n_44),
.B1(n_11),
.B2(n_3),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_1),
.B(n_2),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_3),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_102),
.B(n_3),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_164),
.B(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_119),
.A2(n_44),
.B1(n_5),
.B2(n_6),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_98),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_193),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_101),
.B(n_4),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_90),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_169),
.A2(n_175),
.B1(n_176),
.B2(n_105),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_133),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_96),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_115),
.A2(n_8),
.B1(n_9),
.B2(n_94),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_92),
.A2(n_9),
.B1(n_127),
.B2(n_104),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_108),
.B(n_96),
.C(n_91),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_188),
.C(n_157),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_93),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_133),
.A2(n_100),
.B1(n_89),
.B2(n_107),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_89),
.A2(n_100),
.B(n_107),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_123),
.B(n_91),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_93),
.A2(n_130),
.B1(n_121),
.B2(n_141),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_142),
.Y(n_186)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_88),
.Y(n_187)
);

BUFx2_ASAP7_75t_SL g239 ( 
.A(n_187),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_127),
.B(n_95),
.C(n_109),
.Y(n_188)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_142),
.B(n_88),
.CI(n_103),
.CON(n_189),
.SN(n_189)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_192),
.Y(n_196)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_140),
.Y(n_191)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_106),
.B(n_103),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_194),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_105),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_204),
.A2(n_226),
.B1(n_229),
.B2(n_231),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_205),
.B(n_224),
.C(n_216),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_146),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_206),
.B(n_222),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_212),
.A2(n_189),
.B1(n_150),
.B2(n_182),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_186),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_168),
.B(n_145),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_219),
.B(n_230),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_157),
.B(n_147),
.C(n_188),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_144),
.B(n_159),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_225),
.B(n_160),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_155),
.A2(n_161),
.B1(n_176),
.B2(n_158),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_163),
.A2(n_159),
.B1(n_183),
.B2(n_190),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_172),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_163),
.A2(n_190),
.B1(n_177),
.B2(n_174),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_165),
.B(n_171),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_240),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_190),
.A2(n_173),
.B1(n_154),
.B2(n_184),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_234),
.A2(n_221),
.B1(n_228),
.B2(n_210),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_148),
.B(n_151),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_179),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_149),
.B(n_152),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_231),
.A2(n_167),
.B1(n_191),
.B2(n_173),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_241),
.A2(n_271),
.B1(n_257),
.B2(n_270),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_259),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_184),
.B1(n_180),
.B2(n_156),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_243),
.A2(n_252),
.B1(n_242),
.B2(n_269),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_230),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_244),
.B(n_264),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_211),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_245),
.B(n_255),
.Y(n_291)
);

OAI22x1_ASAP7_75t_L g246 ( 
.A1(n_196),
.A2(n_189),
.B1(n_193),
.B2(n_195),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_247),
.B(n_256),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_248),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_249),
.B(n_251),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_203),
.A2(n_197),
.B1(n_220),
.B2(n_212),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_219),
.B(n_207),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_220),
.B1(n_226),
.B2(n_217),
.Y(n_252)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_254),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_201),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_207),
.B(n_205),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_214),
.Y(n_257)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g259 ( 
.A1(n_209),
.A2(n_199),
.B(n_197),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_233),
.B(n_215),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_261),
.B(n_263),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_209),
.A2(n_203),
.B(n_237),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_262),
.A2(n_239),
.B(n_235),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_215),
.B(n_224),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_209),
.A2(n_208),
.B(n_199),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_198),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_265),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_201),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_279),
.Y(n_302)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_223),
.B(n_202),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_269),
.B(n_272),
.Y(n_304)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_236),
.B(n_200),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_278),
.C(n_280),
.Y(n_313)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_276),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_198),
.B(n_213),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_200),
.B(n_210),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_227),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_227),
.B(n_213),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_281),
.A2(n_300),
.B(n_304),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_235),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_283),
.B(n_287),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_258),
.Y(n_287)
);

AND2x6_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_275),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_276),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_251),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_246),
.C(n_274),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_245),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_293),
.B(n_311),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_297),
.A2(n_305),
.B1(n_298),
.B2(n_310),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_259),
.B(n_252),
.Y(n_300)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_301),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_260),
.A2(n_243),
.B1(n_242),
.B2(n_271),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_305),
.A2(n_310),
.B1(n_254),
.B2(n_273),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_253),
.Y(n_306)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_306),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_247),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_307),
.B(n_279),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_278),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_260),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_315),
.Y(n_343)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_308),
.Y(n_316)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_316),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_317),
.B(n_318),
.C(n_319),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_311),
.C(n_288),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_259),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_308),
.Y(n_321)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_241),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_331),
.C(n_335),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_323),
.B(n_314),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_325),
.A2(n_309),
.B1(n_314),
.B2(n_282),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_327),
.A2(n_338),
.B1(n_296),
.B2(n_303),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_291),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_329),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_291),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_290),
.Y(n_331)
);

NOR2x1p5_ASAP7_75t_SL g332 ( 
.A(n_285),
.B(n_298),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_332),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_300),
.A2(n_285),
.B(n_281),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_333),
.A2(n_284),
.B(n_304),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_306),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_336),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_303),
.B(n_287),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_302),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_337),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_297),
.A2(n_293),
.B1(n_296),
.B2(n_283),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_282),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_342),
.A2(n_333),
.B(n_332),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_338),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_346),
.B(n_357),
.Y(n_383)
);

XNOR2x1_ASAP7_75t_L g366 ( 
.A(n_347),
.B(n_365),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_348),
.A2(n_340),
.B1(n_337),
.B2(n_316),
.Y(n_373)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_349),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_353),
.A2(n_327),
.B1(n_315),
.B2(n_322),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_312),
.Y(n_354)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_354),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_282),
.Y(n_356)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_356),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_324),
.B(n_302),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_319),
.B(n_292),
.C(n_289),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_358),
.B(n_360),
.C(n_339),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_299),
.C(n_294),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_364),
.B(n_320),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_368),
.A2(n_346),
.B1(n_343),
.B2(n_362),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_317),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_374),
.Y(n_398)
);

MAJx2_ASAP7_75t_L g370 ( 
.A(n_352),
.B(n_331),
.C(n_341),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_372),
.Y(n_395)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_371),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_350),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_341),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_324),
.C(n_315),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_381),
.C(n_382),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_315),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_380),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_345),
.A2(n_294),
.B1(n_340),
.B2(n_321),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_379),
.B(n_350),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_294),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_330),
.C(n_301),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_354),
.B(n_301),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_359),
.C(n_354),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_347),
.C(n_364),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_384),
.B(n_359),
.Y(n_385)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_385),
.Y(n_403)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_387),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_390),
.A2(n_393),
.B1(n_394),
.B2(n_396),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_391),
.A2(n_378),
.B(n_366),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_363),
.C(n_353),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_370),
.C(n_376),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_372),
.B(n_363),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_367),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_381),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_399),
.A2(n_380),
.B1(n_369),
.B2(n_377),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_385),
.A2(n_366),
.B(n_382),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_400),
.A2(n_357),
.B(n_349),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_388),
.A2(n_383),
.B(n_368),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_405),
.Y(n_411)
);

AOI31xp33_ASAP7_75t_L g417 ( 
.A1(n_406),
.A2(n_397),
.A3(n_343),
.B(n_355),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_398),
.C(n_395),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_408),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_398),
.C(n_395),
.Y(n_408)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_410),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_403),
.A2(n_404),
.B1(n_409),
.B2(n_402),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_412),
.B(n_413),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_402),
.A2(n_387),
.B1(n_392),
.B2(n_391),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_414),
.B(n_417),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_400),
.B(n_397),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_418),
.B(n_405),
.C(n_407),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_421),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_415),
.B(n_408),
.C(n_348),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_422),
.B(n_423),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_411),
.B(n_361),
.Y(n_423)
);

OA21x2_ASAP7_75t_SL g424 ( 
.A1(n_419),
.A2(n_416),
.B(n_418),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_424),
.B(n_420),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_427),
.B(n_428),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_426),
.B(n_414),
.C(n_355),
.Y(n_428)
);

XNOR2x2_ASAP7_75t_SL g430 ( 
.A(n_429),
.B(n_425),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_344),
.C(n_361),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_431),
.B(n_344),
.Y(n_432)
);


endmodule