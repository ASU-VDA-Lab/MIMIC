module fake_jpeg_23977_n_272 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_19),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_21),
.B1(n_15),
.B2(n_13),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_13),
.B1(n_19),
.B2(n_21),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_46),
.B1(n_52),
.B2(n_32),
.Y(n_61)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_47),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_13),
.B1(n_15),
.B2(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_50),
.Y(n_70)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

AO22x1_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_31),
.B1(n_29),
.B2(n_34),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_49),
.B1(n_54),
.B2(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_62),
.B1(n_34),
.B2(n_54),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_53),
.A2(n_37),
.B1(n_36),
.B2(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_37),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_64),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_37),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_17),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_71),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_28),
.B(n_33),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_73),
.Y(n_87)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_17),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_78),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_74),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_82),
.B1(n_69),
.B2(n_39),
.Y(n_116)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_84),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_36),
.B1(n_49),
.B2(n_34),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_57),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_39),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_65),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_56),
.B1(n_69),
.B2(n_64),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_116),
.B1(n_29),
.B2(n_74),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_108),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_87),
.B1(n_63),
.B2(n_83),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_111),
.B1(n_110),
.B2(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_63),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_109),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_67),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_66),
.B(n_71),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_61),
.B1(n_67),
.B2(n_62),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_60),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_114),
.B(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_60),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_87),
.B1(n_83),
.B2(n_90),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_122),
.B1(n_127),
.B2(n_129),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_60),
.B1(n_84),
.B2(n_64),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_80),
.B1(n_59),
.B2(n_73),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_72),
.B(n_64),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_116),
.B(n_97),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_28),
.C(n_88),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_59),
.B1(n_86),
.B2(n_106),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_138),
.B(n_115),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_107),
.B1(n_111),
.B2(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_59),
.B1(n_86),
.B2(n_46),
.Y(n_134)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_136),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_25),
.B1(n_22),
.B2(n_16),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_147),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_140),
.A2(n_136),
.B1(n_120),
.B2(n_121),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_100),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_29),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_143),
.B(n_145),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_101),
.B(n_102),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_150),
.B1(n_138),
.B2(n_125),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_137),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_102),
.B(n_104),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_97),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_161),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_99),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_155),
.B(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_162),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_27),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_130),
.A2(n_98),
.B(n_103),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_168),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_131),
.C(n_119),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_176),
.C(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_154),
.A2(n_134),
.B1(n_16),
.B2(n_22),
.Y(n_171)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_24),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_174),
.B(n_183),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_25),
.B1(n_26),
.B2(n_18),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_75),
.C(n_74),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_29),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_179),
.C(n_181),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_27),
.C(n_24),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_27),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_139),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_27),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_147),
.C(n_161),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_24),
.B1(n_20),
.B2(n_14),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_149),
.B1(n_162),
.B2(n_157),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_27),
.B1(n_20),
.B2(n_14),
.Y(n_211)
);

AO221x1_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_144),
.B1(n_153),
.B2(n_150),
.C(n_20),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_191),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_140),
.B(n_160),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_199),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_202),
.C(n_20),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_27),
.C(n_24),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_0),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_201),
.B(n_166),
.CI(n_165),
.CON(n_205),
.SN(n_205)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_198),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_211),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_181),
.B1(n_179),
.B2(n_178),
.Y(n_208)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_177),
.B1(n_174),
.B2(n_184),
.Y(n_209)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

NOR3xp33_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_12),
.C(n_11),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_219),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_189),
.C(n_2),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_0),
.C(n_1),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_220),
.C(n_1),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_10),
.B(n_2),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_1),
.C(n_2),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

OAI221xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_192),
.B1(n_203),
.B2(n_200),
.C(n_198),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_215),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_189),
.C(n_202),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_227),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_232),
.C(n_7),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_218),
.B(n_10),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_234),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_231),
.A2(n_219),
.B1(n_208),
.B2(n_210),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_1),
.C(n_3),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_3),
.B(n_4),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_227),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_213),
.B(n_209),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_237),
.A2(n_225),
.B(n_224),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_206),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_242),
.C(n_245),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_223),
.A2(n_220),
.B1(n_205),
.B2(n_5),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_205),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_3),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_3),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_234),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_251),
.B(n_253),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_252),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_4),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_4),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_255),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_250),
.B(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_235),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_258),
.A2(n_261),
.B(n_260),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_238),
.B(n_246),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_SL g262 ( 
.A(n_251),
.B(n_245),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_256),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_264),
.B(n_266),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_265),
.B(n_259),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_268),
.A2(n_263),
.B(n_6),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_267),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_5),
.C(n_7),
.Y(n_272)
);


endmodule