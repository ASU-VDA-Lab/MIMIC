module fake_jpeg_30983_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx2_ASAP7_75t_SL g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx5_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_1),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_14),
.B(n_16),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_11),
.A2(n_1),
.B(n_3),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_18),
.C(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_6),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_8),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_6),
.B1(n_10),
.B2(n_12),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_21),
.A2(n_10),
.B1(n_13),
.B2(n_9),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_27),
.B1(n_22),
.B2(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_20),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_19),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_23),
.C(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_32),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_28),
.B(n_30),
.Y(n_34)
);

AO221x1_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_27),
.B1(n_17),
.B2(n_5),
.C(n_3),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_33),
.C(n_5),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_9),
.B1(n_1),
.B2(n_13),
.Y(n_37)
);


endmodule