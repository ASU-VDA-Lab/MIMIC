module fake_netlist_1_5271_n_31 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_31);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
BUFx8_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
INVxp33_ASAP7_75t_SL g16 ( .A(n_1), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_4), .B(n_1), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_13), .B(n_0), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_16), .B(n_2), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_18), .B(n_17), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_19), .B(n_14), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_14), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AOI22xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_21), .B1(n_15), .B2(n_6), .Y(n_25) );
AOI21xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_3), .B(n_5), .Y(n_26) );
INVxp67_ASAP7_75t_SL g27 ( .A(n_25), .Y(n_27) );
OAI221xp5_ASAP7_75t_R g28 ( .A1(n_27), .A2(n_7), .B1(n_10), .B2(n_11), .C(n_12), .Y(n_28) );
AND2x4_ASAP7_75t_L g29 ( .A(n_28), .B(n_26), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
INVxp67_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
endmodule