module real_jpeg_23154_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_1),
.B(n_80),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_1),
.A2(n_35),
.B1(n_60),
.B2(n_61),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_1),
.A2(n_42),
.B(n_98),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_1),
.B(n_115),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_1),
.A2(n_88),
.B1(n_176),
.B2(n_179),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_1),
.A2(n_37),
.B(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_2),
.A2(n_27),
.B1(n_37),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_2),
.A2(n_60),
.B1(n_61),
.B2(n_69),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_69),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_3),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_26),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_5),
.A2(n_27),
.B1(n_37),
.B2(n_73),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_5),
.A2(n_60),
.B1(n_61),
.B2(n_73),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_73),
.Y(n_176)
);

INVx8_ASAP7_75t_SL g32 ( 
.A(n_6),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_8),
.A2(n_27),
.B1(n_37),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_66),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_8),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_9),
.A2(n_48),
.B1(n_60),
.B2(n_61),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_11),
.A2(n_72),
.B1(n_78),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_11),
.A2(n_27),
.B1(n_37),
.B2(n_83),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_83),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_83),
.Y(n_166)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_13),
.A2(n_60),
.B1(n_61),
.B2(n_95),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_15),
.Y(n_93)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_15),
.Y(n_169)
);

XNOR2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_135),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_117),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_20),
.B(n_117),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_84),
.B1(n_85),
.B2(n_116),
.Y(n_20)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_21),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_55),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_23),
.A2(n_38),
.B1(n_39),
.B2(n_121),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_23),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.A3(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_23)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_27),
.A2(n_37),
.B1(n_59),
.B2(n_63),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_27),
.A2(n_30),
.B1(n_31),
.B2(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_27),
.B(n_35),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_30),
.A2(n_31),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_33),
.A2(n_35),
.B(n_72),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_35),
.A2(n_61),
.B(n_100),
.C(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_35),
.B(n_97),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_35),
.B(n_93),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_37),
.A2(n_59),
.A3(n_61),
.B1(n_192),
.B2(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_49),
.B2(n_53),
.Y(n_39)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_40),
.B(n_94),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_40),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_41),
.A2(n_42),
.B1(n_98),
.B2(n_100),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_41),
.B(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_47),
.A2(n_130),
.B(n_132),
.Y(n_129)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_50),
.A2(n_88),
.B1(n_166),
.B2(n_176),
.Y(n_175)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_70),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_65),
.B(n_67),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_57),
.A2(n_65),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_57),
.A2(n_114),
.B1(n_115),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_57),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_64),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_58),
.A2(n_126),
.B1(n_190),
.B2(n_193),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_58)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_60),
.A2(n_61),
.B1(n_98),
.B2(n_100),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_60),
.B(n_63),
.Y(n_200)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_80),
.B2(n_81),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_74),
.B1(n_80),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_76),
.Y(n_80)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_107),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_96),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B(n_90),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_88),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_88),
.A2(n_90),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_101),
.B(n_102),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_104),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_142)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

BUFx24_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_105),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_146),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_105),
.A2(n_154),
.B1(n_155),
.B2(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.C(n_113),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_113),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_109),
.B(n_154),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.C(n_122),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_118),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_120),
.Y(n_226)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.C(n_128),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_124),
.B(n_211),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_222),
.B(n_227),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_206),
.B(n_221),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_185),
.B(n_205),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_162),
.B(n_184),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_149),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_140),
.B(n_149),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_147),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_142),
.B1(n_147),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_144),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_147),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_157),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_156),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_156),
.C(n_157),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_158),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_172),
.B(n_183),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_164),
.B(n_170),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_177),
.B(n_182),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_174),
.B(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_186),
.B(n_187),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_198),
.B1(n_203),
.B2(n_204),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_188)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_194),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_197),
.C(n_203),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_201),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_207),
.B(n_208),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_216),
.C(n_219),
.Y(n_223)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_214)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);


endmodule