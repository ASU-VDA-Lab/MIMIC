module fake_jpeg_9738_n_251 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_41),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_56),
.Y(n_81)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_36),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_33),
.B(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_20),
.B(n_35),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_30),
.B(n_22),
.C(n_37),
.Y(n_93)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

AO22x1_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_45),
.B1(n_17),
.B2(n_42),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_64),
.B1(n_67),
.B2(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_62),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_20),
.B1(n_33),
.B2(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_37),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_20),
.B1(n_17),
.B2(n_32),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_24),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_72),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_26),
.B1(n_36),
.B2(n_29),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_31),
.B(n_30),
.Y(n_92)
);

OAI32xp33_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_26),
.A3(n_29),
.B1(n_39),
.B2(n_22),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_103),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_SL g113 ( 
.A1(n_76),
.A2(n_101),
.B(n_64),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_77),
.B(n_90),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_79),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_28),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_80),
.A2(n_92),
.B1(n_9),
.B2(n_10),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_87),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_89),
.B1(n_96),
.B2(n_97),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_1),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_93),
.B(n_95),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_27),
.B1(n_30),
.B2(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_27),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_1),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_30),
.B1(n_22),
.B2(n_37),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_48),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_9),
.B(n_10),
.Y(n_129)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_105),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_48),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_103),
.B1(n_11),
.B2(n_13),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_6),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_54),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_85),
.Y(n_138)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_118),
.Y(n_142)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_131),
.B1(n_135),
.B2(n_82),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_116),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_65),
.B1(n_66),
.B2(n_50),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_125),
.B1(n_127),
.B2(n_129),
.Y(n_158)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_81),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_50),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_120),
.B(n_123),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_59),
.B1(n_69),
.B2(n_72),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_78),
.B1(n_84),
.B2(n_94),
.Y(n_139)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_59),
.B1(n_16),
.B2(n_11),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_10),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_130),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_80),
.Y(n_149)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_79),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_133),
.C(n_105),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_144),
.B1(n_145),
.B2(n_151),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_95),
.B(n_88),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_140),
.A2(n_146),
.B(n_147),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_134),
.A2(n_79),
.B1(n_75),
.B2(n_97),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_96),
.B1(n_95),
.B2(n_88),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_90),
.B(n_102),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_105),
.B(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_154),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_86),
.B1(n_82),
.B2(n_106),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_153),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_155),
.B(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_159),
.Y(n_165)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_14),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_135),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_163),
.B(n_173),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_124),
.Y(n_164)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_118),
.Y(n_167)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_177),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_109),
.B1(n_132),
.B2(n_131),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_171),
.A2(n_175),
.B1(n_153),
.B2(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_122),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_174),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_148),
.A2(n_109),
.B1(n_128),
.B2(n_123),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_129),
.B(n_117),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_178),
.B(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_157),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_148),
.A2(n_117),
.B(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_141),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_86),
.Y(n_180)
);

NOR2x1_ASAP7_75t_SL g181 ( 
.A(n_144),
.B(n_125),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_181),
.A2(n_172),
.B(n_145),
.C(n_175),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_146),
.C(n_140),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_192),
.C(n_197),
.Y(n_205)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_195),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_152),
.B1(n_158),
.B2(n_139),
.Y(n_190)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_165),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_191),
.B(n_198),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_151),
.Y(n_192)
);

BUFx24_ASAP7_75t_SL g195 ( 
.A(n_179),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_150),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_180),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_199),
.A2(n_162),
.B1(n_181),
.B2(n_171),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_199),
.B1(n_208),
.B2(n_209),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_166),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_210),
.C(n_184),
.Y(n_218)
);

AOI321xp33_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_196),
.A3(n_192),
.B1(n_176),
.B2(n_194),
.C(n_187),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_207),
.A2(n_186),
.B(n_196),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_213),
.Y(n_221)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_177),
.Y(n_224)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_200),
.C(n_162),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_216),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_173),
.B1(n_199),
.B2(n_191),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_194),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_218),
.C(n_219),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_204),
.B(n_199),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_222),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_201),
.A2(n_199),
.B(n_178),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_223),
.B(n_163),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_208),
.C(n_202),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_193),
.C(n_136),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_206),
.C(n_160),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_210),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_228),
.B(n_229),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_233),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_232),
.A2(n_221),
.B(n_215),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_180),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_217),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_227),
.B(n_231),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_236),
.A2(n_233),
.B(n_145),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_238),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_242),
.Y(n_245)
);

O2A1O1Ixp33_ASAP7_75t_SL g241 ( 
.A1(n_239),
.A2(n_143),
.B(n_159),
.C(n_15),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_15),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_100),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_243),
.B(n_235),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_246),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_245),
.Y(n_250)
);

HAxp5_ASAP7_75t_SL g251 ( 
.A(n_250),
.B(n_247),
.CON(n_251),
.SN(n_251)
);


endmodule