module real_jpeg_31521_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

NAND2x1p5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_12),
.Y(n_11)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_2),
.B(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g10 ( 
.A1(n_4),
.A2(n_11),
.B(n_13),
.Y(n_10)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_14),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_17),
.B1(n_26),
.B2(n_27),
.Y(n_6)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

NAND2x1_ASAP7_75t_SL g7 ( 
.A(n_8),
.B(n_16),
.Y(n_7)
);

NAND2xp67_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_15),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_15),
.B(n_22),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_22),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_20),
.B(n_24),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_18),
.A2(n_20),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_20),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

INVx2_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);


endmodule