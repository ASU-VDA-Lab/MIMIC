module fake_jpeg_12336_n_91 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_91);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_91;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_9),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_0),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_27),
.Y(n_31)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_41),
.Y(n_42)
);

CKINVDCx12_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_13),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_22),
.A2(n_18),
.B1(n_11),
.B2(n_21),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_47),
.Y(n_56)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_11),
.B(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_34),
.B(n_41),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_25),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_41),
.B1(n_32),
.B2(n_37),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_57),
.B1(n_44),
.B2(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_16),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_41),
.B1(n_31),
.B2(n_30),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_62),
.B(n_50),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_67),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_49),
.C(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_68),
.B(n_70),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_62),
.B1(n_53),
.B2(n_59),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_74),
.B1(n_68),
.B2(n_64),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_55),
.B1(n_34),
.B2(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_79),
.Y(n_82)
);

AOI221xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_76),
.B1(n_73),
.B2(n_71),
.C(n_75),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_78),
.A2(n_80),
.B(n_66),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_70),
.C(n_54),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_74),
.B(n_65),
.Y(n_80)
);

OAI21x1_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_17),
.B(n_23),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_7),
.C(n_5),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_14),
.A3(n_16),
.B1(n_17),
.B2(n_6),
.C1(n_7),
.C2(n_5),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_86),
.Y(n_88)
);

AOI21x1_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_23),
.B(n_14),
.Y(n_87)
);

OAI321xp33_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_1),
.A3(n_2),
.B1(n_28),
.B2(n_39),
.C(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_89),
.B(n_1),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_2),
.Y(n_91)
);


endmodule