module fake_jpeg_5569_n_347 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_8),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_20),
.Y(n_55)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_8),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_47),
.Y(n_72)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_0),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_17),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_55),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_53),
.Y(n_85)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_57),
.B(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_24),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_70),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

AO22x1_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_47),
.B1(n_32),
.B2(n_45),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_79),
.Y(n_106)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_21),
.B1(n_29),
.B2(n_32),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_40),
.B1(n_42),
.B2(n_29),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_52),
.B1(n_69),
.B2(n_47),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_90),
.B1(n_91),
.B2(n_52),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_92),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_93),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_42),
.B1(n_40),
.B2(n_21),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_32),
.B1(n_37),
.B2(n_41),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_49),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_69),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_55),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_20),
.B1(n_25),
.B2(n_24),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_62),
.B(n_49),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_75),
.Y(n_105)
);

OR2x4_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_108),
.Y(n_151)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_110),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_61),
.Y(n_108)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_111),
.A2(n_102),
.B1(n_79),
.B2(n_78),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_122),
.B1(n_101),
.B2(n_102),
.Y(n_152)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_117),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_128),
.Y(n_141)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_38),
.Y(n_118)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_37),
.B(n_97),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_25),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_125),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_96),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_72),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_90),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_133),
.Y(n_160)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_89),
.Y(n_142)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_144),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_87),
.B1(n_92),
.B2(n_104),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_113),
.B1(n_109),
.B2(n_122),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_126),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_77),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_36),
.Y(n_184)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_150),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_77),
.C(n_93),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_147),
.B(n_35),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_56),
.B1(n_53),
.B2(n_98),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_153),
.B1(n_105),
.B2(n_129),
.Y(n_169)
);

FAx1_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_36),
.CI(n_39),
.CON(n_149),
.SN(n_149)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_129),
.B(n_120),
.Y(n_164)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_130),
.B1(n_101),
.B2(n_95),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_118),
.Y(n_163)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_159),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_108),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_160),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_161),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_162),
.A2(n_164),
.B1(n_169),
.B2(n_178),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_138),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_118),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_155),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_166),
.B(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_171),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_154),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_133),
.B1(n_110),
.B2(n_132),
.Y(n_178)
);

OAI32xp33_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_109),
.A3(n_113),
.B1(n_128),
.B2(n_116),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_30),
.Y(n_214)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_183),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_182),
.B1(n_153),
.B2(n_149),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_115),
.B1(n_71),
.B2(n_63),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_187),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_60),
.B(n_31),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_186),
.B(n_140),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_31),
.B(n_97),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_175),
.A2(n_149),
.B1(n_155),
.B2(n_159),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_192),
.B(n_195),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_197),
.Y(n_215)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_196),
.Y(n_218)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_136),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_199),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_138),
.C(n_139),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_36),
.Y(n_240)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_210),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_27),
.B(n_30),
.Y(n_235)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_R g211 ( 
.A(n_181),
.B(n_139),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_164),
.B(n_43),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_150),
.Y(n_212)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_163),
.A2(n_158),
.B1(n_145),
.B2(n_63),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_213),
.A2(n_176),
.B1(n_161),
.B2(n_187),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_169),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_181),
.B1(n_170),
.B2(n_183),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_184),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_217),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_236),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_180),
.B1(n_179),
.B2(n_186),
.Y(n_225)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_231),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_238),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_197),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_185),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_26),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_234),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_27),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_199),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_26),
.B(n_33),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_205),
.Y(n_239)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_193),
.C(n_203),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_244),
.C(n_254),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_216),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_198),
.C(n_200),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_246),
.B(n_248),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_219),
.Y(n_248)
);

AO22x1_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_208),
.B1(n_192),
.B2(n_189),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_253),
.A2(n_256),
.B1(n_247),
.B2(n_245),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_223),
.C(n_225),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_210),
.C(n_206),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_257),
.C(n_260),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_231),
.B1(n_217),
.B2(n_238),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_188),
.C(n_204),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_201),
.C(n_191),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_222),
.Y(n_267)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_227),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_263),
.B(n_235),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_260),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_265),
.A2(n_252),
.B1(n_19),
.B2(n_18),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_228),
.B1(n_230),
.B2(n_229),
.Y(n_266)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_278),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_270),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_224),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_SL g286 ( 
.A1(n_271),
.A2(n_261),
.B(n_256),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_249),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_274),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_230),
.B1(n_220),
.B2(n_144),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_282),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_258),
.B(n_257),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_277),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_254),
.B(n_33),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_SL g299 ( 
.A(n_279),
.B(n_281),
.C(n_26),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_135),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_26),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_263),
.B(n_33),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_250),
.A2(n_123),
.B1(n_88),
.B2(n_19),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_88),
.C(n_65),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_19),
.C(n_39),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_291),
.B(n_297),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_255),
.B1(n_283),
.B2(n_259),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_287),
.A2(n_268),
.B1(n_33),
.B2(n_2),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_34),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_39),
.C(n_26),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_296),
.C(n_279),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_275),
.B(n_11),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_270),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_281),
.B(n_271),
.Y(n_301)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_302),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_304),
.C(n_306),
.Y(n_314)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_264),
.Y(n_303)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_285),
.B(n_293),
.Y(n_305)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_305),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_286),
.C(n_4),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_284),
.B(n_33),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_311),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_288),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_4),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_34),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_312),
.B(n_291),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_1),
.C(n_2),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_296),
.C(n_3),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_315),
.A2(n_324),
.B(n_308),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_54),
.B(n_1),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_320),
.B(n_5),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_5),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_5),
.C(n_6),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_316),
.Y(n_326)
);

OAI32xp33_ASAP7_75t_L g338 ( 
.A1(n_326),
.A2(n_321),
.A3(n_34),
.B1(n_23),
.B2(n_12),
.Y(n_338)
);

AOI322xp5_ASAP7_75t_L g335 ( 
.A1(n_327),
.A2(n_328),
.A3(n_332),
.B1(n_315),
.B2(n_324),
.C1(n_10),
.C2(n_12),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_323),
.A2(n_304),
.B1(n_301),
.B2(n_311),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_329),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_330),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_309),
.Y(n_331)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_331),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_314),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_321),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_333),
.A2(n_338),
.B(n_328),
.Y(n_339)
);

NOR2x1_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_7),
.Y(n_341)
);

AOI322xp5_ASAP7_75t_L g342 ( 
.A1(n_339),
.A2(n_340),
.A3(n_341),
.B1(n_336),
.B2(n_337),
.C1(n_12),
.C2(n_13),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_334),
.Y(n_340)
);

OAI311xp33_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_9),
.A3(n_10),
.B1(n_14),
.C1(n_15),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_14),
.B(n_15),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_344),
.B(n_14),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_16),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_16),
.C(n_23),
.Y(n_347)
);


endmodule