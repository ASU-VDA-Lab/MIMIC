module real_aes_7322_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
INVx1_ASAP7_75t_L g512 ( .A(n_1), .Y(n_512) );
INVx1_ASAP7_75t_L g164 ( .A(n_2), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_3), .A2(n_37), .B1(n_189), .B2(n_468), .Y(n_497) );
AOI21xp33_ASAP7_75t_L g208 ( .A1(n_4), .A2(n_180), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_5), .B(n_178), .Y(n_523) );
AND2x6_ASAP7_75t_L g157 ( .A(n_6), .B(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_7), .A2(n_262), .B(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_8), .B(n_38), .Y(n_126) );
INVx1_ASAP7_75t_L g214 ( .A(n_9), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_10), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g149 ( .A(n_11), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_12), .B(n_170), .Y(n_476) );
INVx1_ASAP7_75t_L g268 ( .A(n_13), .Y(n_268) );
INVx1_ASAP7_75t_L g506 ( .A(n_14), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_15), .B(n_145), .Y(n_528) );
AO32x2_ASAP7_75t_L g495 ( .A1(n_16), .A2(n_144), .A3(n_178), .B1(n_470), .B2(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_17), .B(n_189), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_18), .B(n_185), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_19), .B(n_145), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_20), .A2(n_30), .B1(n_744), .B2(n_745), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_20), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_21), .A2(n_49), .B1(n_189), .B2(n_468), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_22), .B(n_180), .Y(n_225) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_23), .A2(n_77), .B1(n_170), .B2(n_189), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_24), .B(n_189), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_25), .B(n_192), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_26), .A2(n_266), .B(n_267), .C(n_269), .Y(n_265) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_27), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_28), .B(n_175), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_29), .B(n_168), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_30), .Y(n_745) );
INVx1_ASAP7_75t_L g203 ( .A(n_31), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_32), .B(n_175), .Y(n_493) );
INVx2_ASAP7_75t_L g155 ( .A(n_33), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_34), .B(n_189), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_35), .B(n_175), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_36), .A2(n_157), .B(n_160), .C(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_38), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g201 ( .A(n_39), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_40), .B(n_168), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_41), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_42), .B(n_189), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_43), .A2(n_87), .B1(n_232), .B2(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_44), .B(n_189), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_45), .B(n_189), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g204 ( .A(n_46), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_47), .B(n_511), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_48), .B(n_180), .Y(n_245) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_50), .A2(n_60), .B1(n_170), .B2(n_189), .Y(n_532) );
AOI222xp33_ASAP7_75t_SL g128 ( .A1(n_51), .A2(n_129), .B1(n_132), .B2(n_732), .C1(n_733), .C2(n_735), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_52), .A2(n_160), .B1(n_170), .B2(n_199), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_53), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_54), .B(n_189), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g151 ( .A(n_55), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_56), .B(n_189), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_57), .A2(n_188), .B(n_212), .C(n_213), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_58), .Y(n_259) );
INVx1_ASAP7_75t_L g210 ( .A(n_59), .Y(n_210) );
INVx1_ASAP7_75t_L g158 ( .A(n_61), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_62), .A2(n_102), .B1(n_115), .B2(n_747), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_63), .B(n_189), .Y(n_513) );
INVx1_ASAP7_75t_L g148 ( .A(n_64), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_65), .Y(n_119) );
AO32x2_ASAP7_75t_L g465 ( .A1(n_66), .A2(n_178), .A3(n_237), .B1(n_466), .B2(n_470), .Y(n_465) );
INVx1_ASAP7_75t_L g545 ( .A(n_67), .Y(n_545) );
INVx1_ASAP7_75t_L g488 ( .A(n_68), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_69), .A2(n_76), .B1(n_130), .B2(n_131), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_69), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_SL g184 ( .A1(n_70), .A2(n_185), .B(n_186), .C(n_188), .Y(n_184) );
INVxp67_ASAP7_75t_L g187 ( .A(n_71), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_72), .B(n_170), .Y(n_489) );
INVx1_ASAP7_75t_L g114 ( .A(n_73), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_74), .Y(n_206) );
INVx1_ASAP7_75t_L g252 ( .A(n_75), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_76), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_78), .A2(n_157), .B(n_160), .C(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_79), .B(n_468), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_80), .B(n_170), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_81), .B(n_165), .Y(n_228) );
INVx2_ASAP7_75t_L g146 ( .A(n_82), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_83), .B(n_185), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_84), .B(n_170), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g159 ( .A1(n_85), .A2(n_157), .B(n_160), .C(n_163), .Y(n_159) );
INVx2_ASAP7_75t_L g111 ( .A(n_86), .Y(n_111) );
OR2x2_ASAP7_75t_L g123 ( .A(n_86), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g135 ( .A(n_86), .B(n_125), .Y(n_135) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_88), .A2(n_100), .B1(n_170), .B2(n_171), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_89), .B(n_175), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_90), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_91), .A2(n_157), .B(n_160), .C(n_240), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_92), .Y(n_247) );
INVx1_ASAP7_75t_L g183 ( .A(n_93), .Y(n_183) );
CKINVDCx16_ASAP7_75t_R g264 ( .A(n_94), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_95), .B(n_165), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_96), .B(n_170), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_97), .B(n_178), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_98), .B(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_99), .A2(n_180), .B(n_181), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g749 ( .A(n_104), .Y(n_749) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .C(n_112), .Y(n_109) );
AND2x2_ASAP7_75t_L g125 ( .A(n_110), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g456 ( .A(n_111), .B(n_125), .Y(n_456) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_111), .B(n_124), .Y(n_737) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AOI22x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_128), .B1(n_738), .B2(n_740), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_120), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g739 ( .A(n_119), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_120), .A2(n_741), .B(n_746), .Y(n_740) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_127), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_123), .Y(n_746) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g732 ( .A(n_129), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_136), .B1(n_454), .B2(n_457), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_133), .A2(n_137), .B1(n_458), .B2(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g741 ( .A1(n_136), .A2(n_137), .B1(n_742), .B2(n_743), .Y(n_741) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR4x1_ASAP7_75t_L g137 ( .A(n_138), .B(n_343), .C(n_403), .D(n_430), .Y(n_137) );
NAND4xp25_ASAP7_75t_SL g138 ( .A(n_139), .B(n_291), .C(n_322), .D(n_339), .Y(n_138) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_216), .B(n_218), .C(n_271), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_194), .Y(n_140) );
INVx1_ASAP7_75t_L g333 ( .A(n_141), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_141), .A2(n_374), .B1(n_422), .B2(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_176), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_142), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g284 ( .A(n_142), .B(n_196), .Y(n_284) );
AND2x2_ASAP7_75t_L g326 ( .A(n_142), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_142), .B(n_217), .Y(n_338) );
INVx1_ASAP7_75t_L g378 ( .A(n_142), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_142), .B(n_432), .Y(n_431) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g306 ( .A(n_143), .B(n_196), .Y(n_306) );
INVx3_ASAP7_75t_L g310 ( .A(n_143), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_143), .B(n_368), .Y(n_367) );
AO21x2_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_150), .B(n_172), .Y(n_143) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_144), .A2(n_197), .B(n_205), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_144), .B(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g233 ( .A(n_144), .Y(n_233) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_145), .Y(n_178) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_146), .B(n_147), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
OAI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_159), .Y(n_150) );
OAI22xp33_ASAP7_75t_L g197 ( .A1(n_152), .A2(n_190), .B1(n_198), .B2(n_204), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_152), .A2(n_252), .B(n_253), .Y(n_251) );
NAND2x1p5_ASAP7_75t_L g152 ( .A(n_153), .B(n_157), .Y(n_152) );
AND2x4_ASAP7_75t_L g180 ( .A(n_153), .B(n_157), .Y(n_180) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_156), .Y(n_153) );
INVx1_ASAP7_75t_L g511 ( .A(n_154), .Y(n_511) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
INVx1_ASAP7_75t_L g171 ( .A(n_155), .Y(n_171) );
INVx1_ASAP7_75t_L g162 ( .A(n_156), .Y(n_162) );
INVx3_ASAP7_75t_L g166 ( .A(n_156), .Y(n_166) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_156), .Y(n_168) );
INVx1_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_156), .Y(n_200) );
INVx4_ASAP7_75t_SL g190 ( .A(n_157), .Y(n_190) );
BUFx3_ASAP7_75t_L g470 ( .A(n_157), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_157), .A2(n_474), .B(n_478), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_157), .A2(n_487), .B(n_490), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_157), .A2(n_505), .B(n_509), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_157), .A2(n_517), .B(n_520), .Y(n_516) );
INVx5_ASAP7_75t_L g182 ( .A(n_160), .Y(n_182) );
AND2x6_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_161), .Y(n_189) );
BUFx3_ASAP7_75t_L g232 ( .A(n_161), .Y(n_232) );
INVx1_ASAP7_75t_L g468 ( .A(n_161), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_167), .C(n_169), .Y(n_163) );
O2A1O1Ixp5_ASAP7_75t_SL g487 ( .A1(n_165), .A2(n_188), .B(n_488), .C(n_489), .Y(n_487) );
INVx2_ASAP7_75t_L g498 ( .A(n_165), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_165), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_165), .A2(n_542), .B(n_543), .Y(n_541) );
INVx5_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_166), .B(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_166), .B(n_214), .Y(n_213) );
OAI22xp5_ASAP7_75t_SL g466 ( .A1(n_166), .A2(n_168), .B1(n_467), .B2(n_469), .Y(n_466) );
INVx2_ASAP7_75t_L g212 ( .A(n_168), .Y(n_212) );
INVx4_ASAP7_75t_L g243 ( .A(n_168), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_168), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_168), .A2(n_498), .B1(n_531), .B2(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_169), .A2(n_506), .B(n_507), .C(n_508), .Y(n_505) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_174), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_174), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g237 ( .A(n_175), .Y(n_237) );
OA21x2_ASAP7_75t_L g260 ( .A1(n_175), .A2(n_261), .B(n_270), .Y(n_260) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_175), .A2(n_473), .B(n_481), .Y(n_472) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_175), .A2(n_486), .B(n_493), .Y(n_485) );
AND2x2_ASAP7_75t_L g397 ( .A(n_176), .B(n_207), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_176), .B(n_310), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_176), .B(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g217 ( .A(n_177), .B(n_196), .Y(n_217) );
INVx1_ASAP7_75t_L g279 ( .A(n_177), .Y(n_279) );
BUFx2_ASAP7_75t_L g283 ( .A(n_177), .Y(n_283) );
AND2x2_ASAP7_75t_L g327 ( .A(n_177), .B(n_195), .Y(n_327) );
OR2x2_ASAP7_75t_L g366 ( .A(n_177), .B(n_195), .Y(n_366) );
AND2x2_ASAP7_75t_L g391 ( .A(n_177), .B(n_207), .Y(n_391) );
AND2x2_ASAP7_75t_L g450 ( .A(n_177), .B(n_280), .Y(n_450) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_191), .Y(n_177) );
INVx4_ASAP7_75t_L g193 ( .A(n_178), .Y(n_193) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_178), .A2(n_516), .B(n_523), .Y(n_515) );
BUFx2_ASAP7_75t_L g262 ( .A(n_180), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_184), .C(n_190), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_182), .A2(n_190), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_182), .A2(n_190), .B(n_264), .C(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g477 ( .A(n_185), .Y(n_477) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_189), .Y(n_244) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_192), .A2(n_208), .B(n_215), .Y(n_207) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_SL g234 ( .A(n_193), .B(n_235), .Y(n_234) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_193), .B(n_470), .C(n_530), .Y(n_529) );
AO21x1_ASAP7_75t_L g576 ( .A1(n_193), .A2(n_530), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g425 ( .A(n_194), .Y(n_425) );
OR2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_207), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_195), .B(n_207), .Y(n_311) );
AND2x2_ASAP7_75t_L g321 ( .A(n_195), .B(n_310), .Y(n_321) );
BUFx2_ASAP7_75t_L g332 ( .A(n_195), .Y(n_332) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g354 ( .A(n_196), .B(n_207), .Y(n_354) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_196), .Y(n_409) );
OAI22xp5_ASAP7_75t_SL g199 ( .A1(n_200), .A2(n_201), .B1(n_202), .B2(n_203), .Y(n_199) );
INVx2_ASAP7_75t_L g202 ( .A(n_200), .Y(n_202) );
INVx4_ASAP7_75t_L g266 ( .A(n_200), .Y(n_266) );
AND2x2_ASAP7_75t_SL g216 ( .A(n_207), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_SL g280 ( .A(n_207), .Y(n_280) );
BUFx2_ASAP7_75t_L g305 ( .A(n_207), .Y(n_305) );
INVx2_ASAP7_75t_L g324 ( .A(n_207), .Y(n_324) );
AND2x2_ASAP7_75t_L g386 ( .A(n_207), .B(n_310), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_212), .A2(n_479), .B(n_480), .Y(n_478) );
O2A1O1Ixp5_ASAP7_75t_L g544 ( .A1(n_212), .A2(n_510), .B(n_545), .C(n_546), .Y(n_544) );
AOI321xp33_ASAP7_75t_L g405 ( .A1(n_216), .A2(n_406), .A3(n_407), .B1(n_408), .B2(n_410), .C(n_411), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_217), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_217), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g399 ( .A(n_217), .B(n_378), .Y(n_399) );
AND2x2_ASAP7_75t_L g432 ( .A(n_217), .B(n_324), .Y(n_432) );
INVx1_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_248), .Y(n_219) );
OR2x2_ASAP7_75t_L g334 ( .A(n_220), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_236), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx3_ASAP7_75t_L g286 ( .A(n_223), .Y(n_286) );
AND2x2_ASAP7_75t_L g296 ( .A(n_223), .B(n_250), .Y(n_296) );
AND2x2_ASAP7_75t_L g301 ( .A(n_223), .B(n_276), .Y(n_301) );
INVx1_ASAP7_75t_L g318 ( .A(n_223), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_223), .B(n_299), .Y(n_337) );
AND2x2_ASAP7_75t_L g342 ( .A(n_223), .B(n_275), .Y(n_342) );
OR2x2_ASAP7_75t_L g374 ( .A(n_223), .B(n_363), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_223), .B(n_287), .Y(n_413) );
AND2x2_ASAP7_75t_L g447 ( .A(n_223), .B(n_273), .Y(n_447) );
OR2x6_ASAP7_75t_L g223 ( .A(n_224), .B(n_234), .Y(n_223) );
AOI21xp5_ASAP7_75t_SL g224 ( .A1(n_225), .A2(n_226), .B(n_233), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_230), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_230), .A2(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g269 ( .A(n_232), .Y(n_269) );
INVx1_ASAP7_75t_L g257 ( .A(n_233), .Y(n_257) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_233), .A2(n_504), .B(n_514), .Y(n_503) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_233), .A2(n_540), .B(n_547), .Y(n_539) );
INVx1_ASAP7_75t_L g274 ( .A(n_236), .Y(n_274) );
INVx2_ASAP7_75t_L g289 ( .A(n_236), .Y(n_289) );
AND2x2_ASAP7_75t_L g329 ( .A(n_236), .B(n_300), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_236), .B(n_276), .Y(n_351) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_246), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_245), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_244), .Y(n_240) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g435 ( .A(n_249), .B(n_286), .Y(n_435) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_260), .Y(n_249) );
INVx2_ASAP7_75t_L g276 ( .A(n_250), .Y(n_276) );
AND2x2_ASAP7_75t_L g429 ( .A(n_250), .B(n_289), .Y(n_429) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_257), .B(n_258), .Y(n_250) );
AND2x2_ASAP7_75t_L g275 ( .A(n_260), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g290 ( .A(n_260), .Y(n_290) );
INVx1_ASAP7_75t_L g300 ( .A(n_260), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_266), .B(n_268), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_266), .A2(n_491), .B(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g508 ( .A(n_266), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_277), .B1(n_281), .B2(n_285), .Y(n_271) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_272), .A2(n_390), .B1(n_427), .B2(n_428), .Y(n_426) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g341 ( .A(n_274), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_275), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g336 ( .A(n_276), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_276), .B(n_289), .Y(n_363) );
INVx1_ASAP7_75t_L g379 ( .A(n_276), .Y(n_379) );
AND2x2_ASAP7_75t_L g320 ( .A(n_278), .B(n_321), .Y(n_320) );
INVx3_ASAP7_75t_SL g359 ( .A(n_278), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_278), .B(n_284), .Y(n_436) );
AND2x4_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g445 ( .A(n_281), .Y(n_445) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_282), .B(n_378), .Y(n_420) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx3_ASAP7_75t_SL g325 ( .A(n_284), .Y(n_325) );
NAND2x1_ASAP7_75t_SL g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x2_ASAP7_75t_L g346 ( .A(n_286), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g353 ( .A(n_286), .B(n_290), .Y(n_353) );
AND2x2_ASAP7_75t_L g358 ( .A(n_286), .B(n_299), .Y(n_358) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_286), .Y(n_407) );
OAI311xp33_ASAP7_75t_L g430 ( .A1(n_287), .A2(n_431), .A3(n_433), .B1(n_434), .C1(n_444), .Y(n_430) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g443 ( .A(n_288), .B(n_316), .Y(n_443) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AND2x2_ASAP7_75t_L g299 ( .A(n_289), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g347 ( .A(n_289), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g402 ( .A(n_289), .Y(n_402) );
INVx1_ASAP7_75t_L g295 ( .A(n_290), .Y(n_295) );
INVx1_ASAP7_75t_L g315 ( .A(n_290), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_290), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g348 ( .A(n_290), .Y(n_348) );
AOI221xp5_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_294), .B1(n_302), .B2(n_307), .C(n_312), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_297), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx4_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
AND2x2_ASAP7_75t_L g410 ( .A(n_296), .B(n_329), .Y(n_410) );
AND2x2_ASAP7_75t_L g417 ( .A(n_296), .B(n_299), .Y(n_417) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_299), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g328 ( .A(n_301), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_304), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g453 ( .A(n_306), .B(n_397), .Y(n_453) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g438 ( .A(n_310), .B(n_366), .Y(n_438) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_311), .A2(n_404), .B(n_405), .C(n_418), .Y(n_403) );
AOI21xp33_ASAP7_75t_SL g312 ( .A1(n_313), .A2(n_317), .B(n_319), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NOR2xp67_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g382 ( .A(n_316), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_317), .A2(n_412), .B1(n_413), .B2(n_414), .C(n_415), .Y(n_411) );
AND2x2_ASAP7_75t_L g388 ( .A(n_318), .B(n_329), .Y(n_388) );
AND2x2_ASAP7_75t_L g441 ( .A(n_318), .B(n_336), .Y(n_441) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_321), .B(n_359), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_326), .B(n_328), .C(n_330), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g369 ( .A(n_324), .B(n_327), .Y(n_369) );
OR2x2_ASAP7_75t_L g412 ( .A(n_324), .B(n_366), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_325), .B(n_391), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_325), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g356 ( .A(n_326), .Y(n_356) );
INVx1_ASAP7_75t_L g422 ( .A(n_329), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .B1(n_337), .B2(n_338), .Y(n_330) );
INVx1_ASAP7_75t_L g345 ( .A(n_331), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_332), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g408 ( .A(n_333), .B(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_L g394 ( .A(n_335), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_336), .B(n_422), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g395 ( .A1(n_337), .A2(n_396), .B1(n_398), .B2(n_400), .Y(n_395) );
INVx1_ASAP7_75t_L g404 ( .A(n_340), .Y(n_404) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g446 ( .A(n_341), .B(n_441), .Y(n_446) );
AOI222xp33_ASAP7_75t_L g375 ( .A1(n_342), .A2(n_376), .B1(n_379), .B2(n_380), .C1(n_383), .C2(n_384), .Y(n_375) );
NAND4xp25_ASAP7_75t_SL g343 ( .A(n_344), .B(n_364), .C(n_375), .D(n_387), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B1(n_349), .B2(n_354), .C(n_355), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_347), .B(n_382), .Y(n_381) );
INVxp67_ASAP7_75t_L g373 ( .A(n_348), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_349), .A2(n_419), .B1(n_421), .B2(n_423), .C(n_426), .Y(n_418) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g361 ( .A(n_353), .B(n_362), .Y(n_361) );
OAI21xp33_ASAP7_75t_L g415 ( .A1(n_354), .A2(n_416), .B(n_417), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B1(n_359), .B2(n_360), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B(n_370), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g406 ( .A(n_377), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_378), .B(n_397), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_378), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_382), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g414 ( .A(n_386), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_392), .B2(n_394), .C(n_395), .Y(n_387) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI222xp33_ASAP7_75t_L g434 ( .A1(n_397), .A2(n_435), .B1(n_436), .B2(n_437), .C1(n_439), .C2(n_442), .Y(n_434) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_401), .B(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g433 ( .A(n_407), .Y(n_433) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp33_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_447), .B2(n_448), .C(n_451), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVxp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g734 ( .A(n_455), .Y(n_734) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND3x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_652), .C(n_700), .Y(n_459) );
NOR4xp25_ASAP7_75t_L g460 ( .A(n_461), .B(n_580), .C(n_625), .D(n_639), .Y(n_460) );
OAI311xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_500), .A3(n_524), .B1(n_533), .C1(n_548), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_471), .Y(n_462) );
OAI21xp33_ASAP7_75t_L g533 ( .A1(n_463), .A2(n_534), .B(n_536), .Y(n_533) );
AND2x2_ASAP7_75t_L g641 ( .A(n_463), .B(n_568), .Y(n_641) );
AND2x2_ASAP7_75t_L g698 ( .A(n_463), .B(n_584), .Y(n_698) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g591 ( .A(n_464), .B(n_494), .Y(n_591) );
AND2x2_ASAP7_75t_L g648 ( .A(n_464), .B(n_596), .Y(n_648) );
INVx1_ASAP7_75t_L g689 ( .A(n_464), .Y(n_689) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_465), .Y(n_557) );
AND2x2_ASAP7_75t_L g598 ( .A(n_465), .B(n_494), .Y(n_598) );
AND2x2_ASAP7_75t_L g602 ( .A(n_465), .B(n_495), .Y(n_602) );
INVx1_ASAP7_75t_L g614 ( .A(n_465), .Y(n_614) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_470), .A2(n_541), .B(n_544), .Y(n_540) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_482), .Y(n_471) );
AND2x2_ASAP7_75t_L g535 ( .A(n_472), .B(n_494), .Y(n_535) );
INVx2_ASAP7_75t_L g569 ( .A(n_472), .Y(n_569) );
AND2x2_ASAP7_75t_L g584 ( .A(n_472), .B(n_495), .Y(n_584) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_472), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_472), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g604 ( .A(n_472), .B(n_567), .Y(n_604) );
INVx1_ASAP7_75t_L g616 ( .A(n_472), .Y(n_616) );
INVx1_ASAP7_75t_L g657 ( .A(n_472), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_472), .B(n_557), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_477), .Y(n_474) );
NOR2xp67_ASAP7_75t_L g482 ( .A(n_483), .B(n_494), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g534 ( .A(n_484), .B(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_484), .Y(n_562) );
AND2x2_ASAP7_75t_SL g615 ( .A(n_484), .B(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g619 ( .A(n_484), .B(n_494), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_484), .B(n_614), .Y(n_677) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g567 ( .A(n_485), .Y(n_567) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_485), .Y(n_583) );
OR2x2_ASAP7_75t_L g656 ( .A(n_485), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g563 ( .A(n_495), .Y(n_563) );
AND2x2_ASAP7_75t_L g568 ( .A(n_495), .B(n_569), .Y(n_568) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_498), .A2(n_510), .B(n_512), .C(n_513), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_498), .A2(n_521), .B(n_522), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_500), .B(n_551), .Y(n_714) );
INVx1_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g684 ( .A(n_501), .B(n_526), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_515), .Y(n_501) );
AND2x2_ASAP7_75t_L g560 ( .A(n_502), .B(n_551), .Y(n_560) );
INVx2_ASAP7_75t_L g572 ( .A(n_502), .Y(n_572) );
AND2x2_ASAP7_75t_L g606 ( .A(n_502), .B(n_554), .Y(n_606) );
AND2x2_ASAP7_75t_L g673 ( .A(n_502), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_503), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g553 ( .A(n_503), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g593 ( .A(n_503), .B(n_515), .Y(n_593) );
AND2x2_ASAP7_75t_L g610 ( .A(n_503), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g536 ( .A(n_515), .B(n_537), .Y(n_536) );
INVx3_ASAP7_75t_L g554 ( .A(n_515), .Y(n_554) );
AND2x2_ASAP7_75t_L g559 ( .A(n_515), .B(n_539), .Y(n_559) );
AND2x2_ASAP7_75t_L g632 ( .A(n_515), .B(n_611), .Y(n_632) );
AND2x2_ASAP7_75t_L g697 ( .A(n_515), .B(n_687), .Y(n_697) );
OAI311xp33_ASAP7_75t_L g580 ( .A1(n_524), .A2(n_581), .A3(n_585), .B1(n_587), .C1(n_607), .Y(n_580) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g592 ( .A(n_525), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g651 ( .A(n_525), .B(n_559), .Y(n_651) );
AND2x2_ASAP7_75t_L g725 ( .A(n_525), .B(n_606), .Y(n_725) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_526), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g660 ( .A(n_526), .Y(n_660) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g551 ( .A(n_527), .Y(n_551) );
NOR2x1_ASAP7_75t_L g623 ( .A(n_527), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g680 ( .A(n_527), .B(n_554), .Y(n_680) );
AND2x4_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g577 ( .A(n_528), .Y(n_577) );
AND2x2_ASAP7_75t_L g555 ( .A(n_535), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g608 ( .A(n_535), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g688 ( .A(n_535), .B(n_689), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_536), .A2(n_568), .B1(n_588), .B2(n_592), .C(n_594), .Y(n_587) );
INVx1_ASAP7_75t_L g712 ( .A(n_537), .Y(n_712) );
OR2x2_ASAP7_75t_L g678 ( .A(n_538), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g573 ( .A(n_539), .B(n_554), .Y(n_573) );
OR2x2_ASAP7_75t_L g575 ( .A(n_539), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g600 ( .A(n_539), .Y(n_600) );
INVx2_ASAP7_75t_L g611 ( .A(n_539), .Y(n_611) );
AND2x2_ASAP7_75t_L g638 ( .A(n_539), .B(n_576), .Y(n_638) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_539), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_555), .B1(n_558), .B2(n_561), .C(n_564), .Y(n_548) );
INVx1_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
AND2x2_ASAP7_75t_L g649 ( .A(n_551), .B(n_559), .Y(n_649) );
AND2x2_ASAP7_75t_L g699 ( .A(n_551), .B(n_553), .Y(n_699) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g586 ( .A(n_553), .B(n_557), .Y(n_586) );
AND2x2_ASAP7_75t_L g665 ( .A(n_553), .B(n_638), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_554), .B(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g624 ( .A(n_554), .Y(n_624) );
OAI21xp33_ASAP7_75t_L g634 ( .A1(n_555), .A2(n_635), .B(n_637), .Y(n_634) );
OR2x2_ASAP7_75t_L g578 ( .A(n_556), .B(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g644 ( .A(n_556), .B(n_604), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_556), .B(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g621 ( .A(n_557), .B(n_590), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_557), .B(n_704), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_558), .B(n_584), .Y(n_694) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g617 ( .A(n_559), .B(n_572), .Y(n_617) );
INVx1_ASAP7_75t_L g633 ( .A(n_560), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_570), .B1(n_574), .B2(n_578), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx2_ASAP7_75t_L g596 ( .A(n_567), .Y(n_596) );
INVx1_ASAP7_75t_L g609 ( .A(n_567), .Y(n_609) );
INVx1_ASAP7_75t_L g579 ( .A(n_568), .Y(n_579) );
AND2x2_ASAP7_75t_L g650 ( .A(n_568), .B(n_596), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_568), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
OR2x2_ASAP7_75t_L g574 ( .A(n_571), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_571), .B(n_687), .Y(n_686) );
NOR2xp67_ASAP7_75t_L g718 ( .A(n_571), .B(n_719), .Y(n_718) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g721 ( .A(n_573), .B(n_673), .Y(n_721) );
INVx1_ASAP7_75t_SL g687 ( .A(n_575), .Y(n_687) );
AND2x2_ASAP7_75t_L g627 ( .A(n_576), .B(n_611), .Y(n_627) );
INVx1_ASAP7_75t_L g674 ( .A(n_576), .Y(n_674) );
OAI222xp33_ASAP7_75t_L g715 ( .A1(n_581), .A2(n_671), .B1(n_716), .B2(n_717), .C1(n_720), .C2(n_722), .Y(n_715) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g636 ( .A(n_583), .Y(n_636) );
AND2x2_ASAP7_75t_L g647 ( .A(n_584), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_584), .B(n_689), .Y(n_716) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_586), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g691 ( .A(n_588), .Y(n_691) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_SL g629 ( .A(n_591), .Y(n_629) );
AND2x2_ASAP7_75t_L g708 ( .A(n_591), .B(n_669), .Y(n_708) );
AND2x2_ASAP7_75t_L g731 ( .A(n_591), .B(n_615), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_593), .B(n_627), .Y(n_626) );
OAI32xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .A3(n_599), .B1(n_601), .B2(n_605), .Y(n_594) );
BUFx2_ASAP7_75t_L g669 ( .A(n_596), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_597), .B(n_615), .Y(n_696) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g635 ( .A(n_598), .B(n_636), .Y(n_635) );
AND2x4_ASAP7_75t_L g703 ( .A(n_598), .B(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g692 ( .A(n_599), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g663 ( .A(n_602), .B(n_636), .Y(n_663) );
INVx2_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
OAI221xp5_ASAP7_75t_SL g625 ( .A1(n_604), .A2(n_626), .B1(n_628), .B2(n_630), .C(n_634), .Y(n_625) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g637 ( .A(n_606), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g643 ( .A(n_606), .B(n_627), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_610), .B1(n_612), .B2(n_617), .C(n_618), .Y(n_607) );
INVx1_ASAP7_75t_L g726 ( .A(n_608), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_609), .B(n_703), .Y(n_702) );
NAND2x1p5_ASAP7_75t_L g622 ( .A(n_610), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_615), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g681 ( .A(n_615), .Y(n_681) );
BUFx3_ASAP7_75t_L g704 ( .A(n_616), .Y(n_704) );
INVx1_ASAP7_75t_SL g645 ( .A(n_617), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_617), .B(n_659), .Y(n_658) );
AOI21xp33_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_620), .B(n_622), .Y(n_618) );
OAI221xp5_ASAP7_75t_L g723 ( .A1(n_619), .A2(n_720), .B1(n_724), .B2(n_726), .C(n_727), .Y(n_723) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g666 ( .A(n_624), .B(n_627), .Y(n_666) );
INVx1_ASAP7_75t_L g730 ( .A(n_624), .Y(n_730) );
INVx2_ASAP7_75t_L g719 ( .A(n_627), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_627), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g672 ( .A(n_632), .B(n_673), .Y(n_672) );
OAI221xp5_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_642), .B1(n_644), .B2(n_645), .C(n_646), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B1(n_650), .B2(n_651), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_648), .A2(n_710), .B1(n_711), .B2(n_713), .Y(n_709) );
OAI21xp5_ASAP7_75t_L g727 ( .A1(n_651), .A2(n_728), .B(n_731), .Y(n_727) );
NOR4xp25_ASAP7_75t_SL g652 ( .A(n_653), .B(n_661), .C(n_670), .D(n_690), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_658), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_664), .B1(n_667), .B2(n_668), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g706 ( .A(n_666), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_675), .B1(n_678), .B2(n_681), .C(n_682), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g693 ( .A(n_673), .Y(n_693) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI21xp5_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_685), .B(n_688), .Y(n_682) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI211xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B(n_694), .C(n_695), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_695) );
CKINVDCx14_ASAP7_75t_R g705 ( .A(n_699), .Y(n_705) );
NOR3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_715), .C(n_723), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_705), .B1(n_706), .B2(n_707), .C(n_709), .Y(n_701) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
CKINVDCx16_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx3_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
endmodule