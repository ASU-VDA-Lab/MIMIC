module real_aes_9020_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_404;
wire n_147;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g183 ( .A1(n_0), .A2(n_184), .B(n_185), .C(n_189), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_1), .B(n_178), .Y(n_191) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_3), .B(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_4), .A2(n_172), .B(n_478), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_5), .A2(n_152), .B(n_169), .C(n_522), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_6), .A2(n_172), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_7), .B(n_178), .Y(n_484) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_8), .A2(n_144), .B(n_266), .Y(n_265) );
AND2x6_ASAP7_75t_L g169 ( .A(n_9), .B(n_170), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_10), .A2(n_152), .B(n_169), .C(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g575 ( .A(n_11), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_12), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_12), .B(n_40), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_13), .B(n_188), .Y(n_524) );
INVx1_ASAP7_75t_L g149 ( .A(n_14), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_15), .B(n_163), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_16), .A2(n_164), .B(n_533), .C(n_535), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_17), .B(n_178), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_18), .B(n_206), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_19), .A2(n_152), .B(n_198), .C(n_205), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_20), .A2(n_187), .B(n_240), .C(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_21), .B(n_188), .Y(n_506) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_22), .A2(n_454), .B1(n_723), .B2(n_724), .C1(n_733), .C2(n_737), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_23), .B(n_188), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g502 ( .A(n_24), .Y(n_502) );
INVx1_ASAP7_75t_L g472 ( .A(n_25), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_26), .A2(n_152), .B(n_205), .C(n_269), .Y(n_268) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_27), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_28), .Y(n_520) );
INVx1_ASAP7_75t_L g496 ( .A(n_29), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_30), .A2(n_172), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_31), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g154 ( .A(n_32), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_33), .A2(n_167), .B(n_221), .C(n_222), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_34), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_35), .A2(n_187), .B(n_481), .C(n_483), .Y(n_480) );
INVxp67_ASAP7_75t_L g497 ( .A(n_36), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_37), .B(n_271), .Y(n_270) );
CKINVDCx14_ASAP7_75t_R g479 ( .A(n_38), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_39), .A2(n_152), .B(n_205), .C(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g114 ( .A(n_40), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_L g572 ( .A1(n_41), .A2(n_189), .B(n_573), .C(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_42), .B(n_196), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_43), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_44), .B(n_163), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_45), .B(n_172), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_46), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_47), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_48), .A2(n_167), .B(n_221), .C(n_249), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_49), .A2(n_105), .B1(n_115), .B2(n_740), .Y(n_104) );
INVx1_ASAP7_75t_L g186 ( .A(n_50), .Y(n_186) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_51), .A2(n_67), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_51), .Y(n_132) );
INVx1_ASAP7_75t_L g250 ( .A(n_52), .Y(n_250) );
INVx1_ASAP7_75t_L g540 ( .A(n_53), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_54), .B(n_172), .Y(n_247) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_55), .A2(n_72), .B1(n_135), .B2(n_136), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_55), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_56), .Y(n_210) );
CKINVDCx14_ASAP7_75t_R g571 ( .A(n_57), .Y(n_571) );
INVx1_ASAP7_75t_L g170 ( .A(n_58), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_59), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_60), .B(n_178), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_61), .A2(n_159), .B(n_204), .C(n_261), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_62), .A2(n_71), .B1(n_730), .B2(n_731), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_62), .Y(n_730) );
INVx1_ASAP7_75t_L g148 ( .A(n_63), .Y(n_148) );
INVx1_ASAP7_75t_SL g482 ( .A(n_64), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_65), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_66), .B(n_163), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_67), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_67), .B(n_178), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_68), .B(n_164), .Y(n_237) );
INVx1_ASAP7_75t_L g505 ( .A(n_69), .Y(n_505) );
CKINVDCx16_ASAP7_75t_R g181 ( .A(n_70), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_71), .Y(n_731) );
INVx1_ASAP7_75t_L g136 ( .A(n_72), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_73), .B(n_200), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_74), .A2(n_152), .B(n_157), .C(n_167), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_75), .Y(n_259) );
INVx1_ASAP7_75t_L g112 ( .A(n_76), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_77), .A2(n_172), .B(n_570), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_78), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_79), .A2(n_172), .B(n_530), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_80), .A2(n_196), .B(n_492), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g469 ( .A(n_81), .Y(n_469) );
INVx1_ASAP7_75t_L g531 ( .A(n_82), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_83), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_83), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_84), .B(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_85), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_86), .A2(n_172), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g534 ( .A(n_87), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_88), .A2(n_725), .B1(n_726), .B2(n_732), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_88), .Y(n_725) );
INVx2_ASAP7_75t_L g146 ( .A(n_89), .Y(n_146) );
INVx1_ASAP7_75t_L g523 ( .A(n_90), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_91), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_92), .B(n_188), .Y(n_238) );
INVx2_ASAP7_75t_L g109 ( .A(n_93), .Y(n_109) );
OR2x2_ASAP7_75t_L g125 ( .A(n_93), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g458 ( .A(n_93), .B(n_127), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_94), .A2(n_152), .B(n_167), .C(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_95), .B(n_172), .Y(n_219) );
INVx1_ASAP7_75t_L g223 ( .A(n_96), .Y(n_223) );
INVxp67_ASAP7_75t_L g262 ( .A(n_97), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_98), .B(n_144), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g158 ( .A(n_100), .Y(n_158) );
INVx1_ASAP7_75t_L g233 ( .A(n_101), .Y(n_233) );
INVx2_ASAP7_75t_L g543 ( .A(n_102), .Y(n_543) );
AND2x2_ASAP7_75t_L g252 ( .A(n_103), .B(n_208), .Y(n_252) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g741 ( .A(n_106), .Y(n_741) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_113), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g127 ( .A(n_108), .B(n_128), .Y(n_127) );
OR2x2_ASAP7_75t_L g722 ( .A(n_109), .B(n_127), .Y(n_722) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_109), .B(n_126), .Y(n_739) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_452), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_117), .B(n_449), .C(n_453), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_129), .B(n_449), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_125), .Y(n_451) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_133), .B1(n_447), .B2(n_448), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_130), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_133), .Y(n_448) );
XNOR2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_137), .Y(n_133) );
INVx1_ASAP7_75t_L g455 ( .A(n_137), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_137), .A2(n_460), .B1(n_734), .B2(n_735), .Y(n_733) );
OR3x1_ASAP7_75t_L g137 ( .A(n_138), .B(n_355), .C(n_404), .Y(n_137) );
NAND5xp2_ASAP7_75t_L g138 ( .A(n_139), .B(n_289), .C(n_318), .D(n_326), .E(n_341), .Y(n_138) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_212), .B(n_228), .C(n_273), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_192), .Y(n_140) );
AND2x2_ASAP7_75t_L g284 ( .A(n_141), .B(n_281), .Y(n_284) );
AND2x2_ASAP7_75t_L g317 ( .A(n_141), .B(n_193), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_141), .B(n_216), .Y(n_410) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_177), .Y(n_141) );
INVx2_ASAP7_75t_L g215 ( .A(n_142), .Y(n_215) );
BUFx2_ASAP7_75t_L g384 ( .A(n_142), .Y(n_384) );
AO21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_150), .B(n_175), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_143), .B(n_176), .Y(n_175) );
INVx3_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_143), .B(n_227), .Y(n_226) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_143), .A2(n_232), .B(n_242), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_143), .B(n_475), .Y(n_474) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_143), .A2(n_501), .B(n_508), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_143), .B(n_526), .Y(n_525) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_144), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_144), .A2(n_267), .B(n_268), .Y(n_266) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g244 ( .A(n_145), .Y(n_244) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
AND2x2_ASAP7_75t_SL g208 ( .A(n_146), .B(n_147), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_171), .Y(n_150) );
INVx5_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_153), .Y(n_166) );
BUFx3_ASAP7_75t_L g190 ( .A(n_153), .Y(n_190) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g174 ( .A(n_154), .Y(n_174) );
INVx1_ASAP7_75t_L g241 ( .A(n_154), .Y(n_241) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_156), .Y(n_161) );
INVx3_ASAP7_75t_L g164 ( .A(n_156), .Y(n_164) );
AND2x2_ASAP7_75t_L g173 ( .A(n_156), .B(n_174), .Y(n_173) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_156), .Y(n_188) );
INVx1_ASAP7_75t_L g271 ( .A(n_156), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_162), .C(n_165), .Y(n_157) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_160), .A2(n_163), .B1(n_496), .B2(n_497), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_160), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_160), .B(n_543), .Y(n_542) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g200 ( .A(n_161), .Y(n_200) );
INVx2_ASAP7_75t_L g184 ( .A(n_163), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_163), .B(n_262), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_163), .A2(n_203), .B(n_472), .C(n_473), .Y(n_471) );
INVx5_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_164), .B(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g483 ( .A(n_166), .Y(n_483) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_SL g180 ( .A1(n_168), .A2(n_181), .B(n_182), .C(n_183), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_168), .A2(n_182), .B(n_259), .C(n_260), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_168), .A2(n_182), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g492 ( .A1(n_168), .A2(n_182), .B(n_493), .C(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_168), .A2(n_182), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_SL g539 ( .A1(n_168), .A2(n_182), .B(n_540), .C(n_541), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_SL g570 ( .A1(n_168), .A2(n_182), .B(n_571), .C(n_572), .Y(n_570) );
INVx4_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
AND2x4_ASAP7_75t_L g172 ( .A(n_169), .B(n_173), .Y(n_172) );
BUFx3_ASAP7_75t_L g205 ( .A(n_169), .Y(n_205) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_169), .B(n_173), .Y(n_234) );
BUFx2_ASAP7_75t_L g196 ( .A(n_172), .Y(n_196) );
INVx1_ASAP7_75t_L g204 ( .A(n_174), .Y(n_204) );
AND2x2_ASAP7_75t_L g192 ( .A(n_177), .B(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g282 ( .A(n_177), .Y(n_282) );
AND2x2_ASAP7_75t_L g368 ( .A(n_177), .B(n_281), .Y(n_368) );
AND2x2_ASAP7_75t_L g423 ( .A(n_177), .B(n_215), .Y(n_423) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_191), .Y(n_177) );
INVx2_ASAP7_75t_L g221 ( .A(n_182), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_187), .B(n_482), .Y(n_481) );
INVx4_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g573 ( .A(n_188), .Y(n_573) );
INVx2_ASAP7_75t_L g507 ( .A(n_189), .Y(n_507) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_190), .Y(n_225) );
INVx1_ASAP7_75t_L g535 ( .A(n_190), .Y(n_535) );
INVx1_ASAP7_75t_L g340 ( .A(n_192), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_192), .B(n_216), .Y(n_387) );
INVx5_ASAP7_75t_L g281 ( .A(n_193), .Y(n_281) );
AND2x4_ASAP7_75t_L g302 ( .A(n_193), .B(n_282), .Y(n_302) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_193), .Y(n_324) );
AND2x2_ASAP7_75t_L g399 ( .A(n_193), .B(n_384), .Y(n_399) );
AND2x2_ASAP7_75t_L g402 ( .A(n_193), .B(n_217), .Y(n_402) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_209), .Y(n_193) );
AOI21xp5_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_197), .B(n_206), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_201), .B(n_203), .Y(n_198) );
INVx2_ASAP7_75t_L g202 ( .A(n_200), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_202), .A2(n_223), .B(n_224), .C(n_225), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_202), .A2(n_225), .B(n_250), .C(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g504 ( .A1(n_202), .A2(n_505), .B(n_506), .C(n_507), .Y(n_504) );
O2A1O1Ixp5_ASAP7_75t_L g522 ( .A1(n_202), .A2(n_507), .B(n_523), .C(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_204), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_207), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g211 ( .A(n_208), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_208), .A2(n_219), .B(n_220), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_208), .A2(n_247), .B(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_208), .A2(n_234), .B(n_469), .C(n_470), .Y(n_468) );
OA21x2_ASAP7_75t_L g568 ( .A1(n_208), .A2(n_569), .B(n_576), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_211), .A2(n_519), .B(n_525), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_212), .B(n_282), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_212), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_216), .Y(n_213) );
AND2x2_ASAP7_75t_L g307 ( .A(n_214), .B(n_282), .Y(n_307) );
AND2x2_ASAP7_75t_L g325 ( .A(n_214), .B(n_217), .Y(n_325) );
INVx1_ASAP7_75t_L g345 ( .A(n_214), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_214), .B(n_281), .Y(n_390) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_214), .Y(n_432) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_215), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_216), .B(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_216), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_216), .A2(n_277), .B(n_338), .C(n_340), .Y(n_337) );
AND2x2_ASAP7_75t_L g344 ( .A(n_216), .B(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g353 ( .A(n_216), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g357 ( .A(n_216), .B(n_281), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_216), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g372 ( .A(n_216), .B(n_282), .Y(n_372) );
AND2x2_ASAP7_75t_L g422 ( .A(n_216), .B(n_423), .Y(n_422) );
INVx5_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g286 ( .A(n_217), .Y(n_286) );
AND2x2_ASAP7_75t_L g327 ( .A(n_217), .B(n_280), .Y(n_327) );
AND2x2_ASAP7_75t_L g339 ( .A(n_217), .B(n_314), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_217), .B(n_368), .Y(n_386) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_226), .Y(n_217) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_253), .Y(n_228) );
INVx1_ASAP7_75t_L g275 ( .A(n_229), .Y(n_275) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_245), .Y(n_229) );
OR2x2_ASAP7_75t_L g277 ( .A(n_230), .B(n_245), .Y(n_277) );
NAND3xp33_ASAP7_75t_L g283 ( .A(n_230), .B(n_284), .C(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_230), .B(n_255), .Y(n_294) );
OR2x2_ASAP7_75t_L g309 ( .A(n_230), .B(n_297), .Y(n_309) );
AND2x2_ASAP7_75t_L g315 ( .A(n_230), .B(n_264), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_230), .B(n_446), .Y(n_445) );
INVx5_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_231), .B(n_255), .Y(n_312) );
AND2x2_ASAP7_75t_L g351 ( .A(n_231), .B(n_265), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_231), .B(n_264), .Y(n_379) );
OR2x2_ASAP7_75t_L g382 ( .A(n_231), .B(n_264), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_235), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_234), .A2(n_502), .B(n_503), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_234), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_239), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_239), .A2(n_270), .B(n_272), .Y(n_269) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx2_ASAP7_75t_L g490 ( .A(n_244), .Y(n_490) );
INVx5_ASAP7_75t_SL g297 ( .A(n_245), .Y(n_297) );
OR2x2_ASAP7_75t_L g303 ( .A(n_245), .B(n_254), .Y(n_303) );
AND2x2_ASAP7_75t_L g319 ( .A(n_245), .B(n_320), .Y(n_319) );
AOI321xp33_ASAP7_75t_L g326 ( .A1(n_245), .A2(n_327), .A3(n_328), .B1(n_329), .B2(n_335), .C(n_337), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_245), .B(n_253), .Y(n_336) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_245), .Y(n_349) );
OR2x2_ASAP7_75t_L g396 ( .A(n_245), .B(n_294), .Y(n_396) );
AND2x2_ASAP7_75t_L g418 ( .A(n_245), .B(n_315), .Y(n_418) );
AND2x2_ASAP7_75t_L g437 ( .A(n_245), .B(n_255), .Y(n_437) );
OR2x6_ASAP7_75t_L g245 ( .A(n_246), .B(n_252), .Y(n_245) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_264), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_255), .B(n_264), .Y(n_278) );
AND2x2_ASAP7_75t_L g287 ( .A(n_255), .B(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g314 ( .A(n_255), .Y(n_314) );
AND2x2_ASAP7_75t_L g320 ( .A(n_255), .B(n_315), .Y(n_320) );
INVxp67_ASAP7_75t_L g350 ( .A(n_255), .Y(n_350) );
OR2x2_ASAP7_75t_L g392 ( .A(n_255), .B(n_297), .Y(n_392) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B(n_263), .Y(n_255) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_256), .A2(n_477), .B(n_484), .Y(n_476) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_256), .A2(n_529), .B(n_536), .Y(n_528) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_256), .A2(n_538), .B(n_544), .Y(n_537) );
OR2x2_ASAP7_75t_L g274 ( .A(n_264), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_SL g288 ( .A(n_264), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_264), .B(n_277), .Y(n_321) );
AND2x2_ASAP7_75t_L g370 ( .A(n_264), .B(n_314), .Y(n_370) );
AND2x2_ASAP7_75t_L g408 ( .A(n_264), .B(n_297), .Y(n_408) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_265), .B(n_297), .Y(n_296) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_276), .B(n_279), .C(n_283), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_274), .A2(n_276), .B1(n_401), .B2(n_403), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_276), .A2(n_299), .B1(n_354), .B2(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_SL g428 ( .A(n_277), .Y(n_428) );
INVx1_ASAP7_75t_SL g328 ( .A(n_278), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_280), .B(n_300), .Y(n_330) );
AOI222xp33_ASAP7_75t_L g341 ( .A1(n_280), .A2(n_321), .B1(n_328), .B2(n_342), .C1(n_346), .C2(n_352), .Y(n_341) );
AND2x2_ASAP7_75t_L g431 ( .A(n_280), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx2_ASAP7_75t_L g306 ( .A(n_281), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_281), .B(n_301), .Y(n_376) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_281), .Y(n_413) );
AND2x2_ASAP7_75t_L g416 ( .A(n_281), .B(n_325), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_281), .B(n_432), .Y(n_442) );
INVx1_ASAP7_75t_L g333 ( .A(n_282), .Y(n_333) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_282), .Y(n_361) );
O2A1O1Ixp33_ASAP7_75t_L g424 ( .A1(n_284), .A2(n_425), .B(n_426), .C(n_429), .Y(n_424) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NAND3xp33_ASAP7_75t_L g347 ( .A(n_286), .B(n_348), .C(n_351), .Y(n_347) );
OR2x2_ASAP7_75t_L g375 ( .A(n_286), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_286), .B(n_302), .Y(n_403) );
OR2x2_ASAP7_75t_L g308 ( .A(n_288), .B(n_309), .Y(n_308) );
AOI211xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_292), .B(n_298), .C(n_310), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_291), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g397 ( .A(n_292), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_293), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g311 ( .A(n_296), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_297), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g365 ( .A(n_297), .B(n_315), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_297), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_297), .B(n_314), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_303), .B1(n_304), .B2(n_308), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_300), .B(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_302), .B(n_344), .Y(n_343) );
OAI221xp5_ASAP7_75t_SL g366 ( .A1(n_303), .A2(n_367), .B1(n_369), .B2(n_371), .C(n_373), .Y(n_366) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x2_ASAP7_75t_L g421 ( .A(n_306), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g434 ( .A(n_306), .B(n_423), .Y(n_434) );
INVx1_ASAP7_75t_L g354 ( .A(n_307), .Y(n_354) );
INVx1_ASAP7_75t_L g425 ( .A(n_308), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_309), .A2(n_392), .B(n_415), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_313), .B(n_316), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI21xp5_ASAP7_75t_SL g318 ( .A1(n_319), .A2(n_321), .B(n_322), .Y(n_318) );
INVx1_ASAP7_75t_L g358 ( .A(n_319), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_320), .A2(n_406), .B1(n_409), .B2(n_411), .C(n_414), .Y(n_405) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_328), .A2(n_418), .B1(n_419), .B2(n_421), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g394 ( .A(n_330), .Y(n_394) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR2xp67_ASAP7_75t_SL g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g398 ( .A(n_334), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g363 ( .A(n_339), .Y(n_363) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_344), .B(n_368), .Y(n_420) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_350), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g436 ( .A(n_351), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g443 ( .A(n_351), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI211xp5_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_358), .B(n_359), .C(n_393), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI211xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B(n_366), .C(n_385), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g446 ( .A(n_370), .Y(n_446) );
AND2x2_ASAP7_75t_L g383 ( .A(n_372), .B(n_384), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .B1(n_381), .B2(n_383), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
OR2x2_ASAP7_75t_L g391 ( .A(n_379), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g444 ( .A(n_380), .Y(n_444) );
INVxp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI31xp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .A3(n_388), .B(n_391), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI211xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B(n_397), .C(n_400), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
CKINVDCx16_ASAP7_75t_R g401 ( .A(n_402), .Y(n_401) );
NAND5xp2_ASAP7_75t_L g404 ( .A(n_405), .B(n_417), .C(n_424), .D(n_438), .E(n_441), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_416), .A2(n_442), .B1(n_443), .B2(n_445), .Y(n_441) );
INVx1_ASAP7_75t_SL g440 ( .A(n_418), .Y(n_440) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI21xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_433), .B(n_435), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OAI22xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_456), .B1(n_459), .B2(n_722), .Y(n_454) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g734 ( .A(n_457), .Y(n_734) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR3x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_633), .C(n_680), .Y(n_460) );
NAND3xp33_ASAP7_75t_SL g461 ( .A(n_462), .B(n_579), .C(n_604), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_517), .B1(n_545), .B2(n_548), .C(n_556), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_485), .B(n_510), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_465), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_465), .B(n_561), .Y(n_677) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_476), .Y(n_465) );
AND2x2_ASAP7_75t_L g547 ( .A(n_466), .B(n_516), .Y(n_547) );
AND2x2_ASAP7_75t_L g597 ( .A(n_466), .B(n_515), .Y(n_597) );
AND2x2_ASAP7_75t_L g618 ( .A(n_466), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g623 ( .A(n_466), .B(n_590), .Y(n_623) );
OR2x2_ASAP7_75t_L g631 ( .A(n_466), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g703 ( .A(n_466), .B(n_499), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_466), .B(n_652), .Y(n_717) );
INVx3_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g562 ( .A(n_467), .B(n_476), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_467), .B(n_499), .Y(n_563) );
AND2x4_ASAP7_75t_L g585 ( .A(n_467), .B(n_516), .Y(n_585) );
AND2x2_ASAP7_75t_L g615 ( .A(n_467), .B(n_487), .Y(n_615) );
AND2x2_ASAP7_75t_L g624 ( .A(n_467), .B(n_614), .Y(n_624) );
AND2x2_ASAP7_75t_L g640 ( .A(n_467), .B(n_500), .Y(n_640) );
OR2x2_ASAP7_75t_L g649 ( .A(n_467), .B(n_632), .Y(n_649) );
AND2x2_ASAP7_75t_L g655 ( .A(n_467), .B(n_590), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_467), .B(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g669 ( .A(n_467), .B(n_512), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_467), .B(n_558), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_467), .B(n_619), .Y(n_708) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_474), .Y(n_467) );
INVx2_ASAP7_75t_L g516 ( .A(n_476), .Y(n_516) );
AND2x2_ASAP7_75t_L g614 ( .A(n_476), .B(n_499), .Y(n_614) );
AND2x2_ASAP7_75t_L g619 ( .A(n_476), .B(n_500), .Y(n_619) );
INVx1_ASAP7_75t_L g675 ( .A(n_476), .Y(n_675) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g584 ( .A(n_486), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_499), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_487), .B(n_547), .Y(n_546) );
BUFx3_ASAP7_75t_L g561 ( .A(n_487), .Y(n_561) );
OR2x2_ASAP7_75t_L g632 ( .A(n_487), .B(n_499), .Y(n_632) );
OR2x2_ASAP7_75t_L g693 ( .A(n_487), .B(n_600), .Y(n_693) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_491), .B(n_498), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_489), .A2(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g513 ( .A(n_491), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_498), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_499), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g652 ( .A(n_499), .B(n_512), .Y(n_652) );
INVx2_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g591 ( .A(n_500), .Y(n_591) );
INVx1_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_511), .A2(n_697), .B1(n_701), .B2(n_704), .C(n_705), .Y(n_696) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_515), .Y(n_511) );
INVx1_ASAP7_75t_SL g559 ( .A(n_512), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_512), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g691 ( .A(n_512), .B(n_547), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_515), .B(n_561), .Y(n_683) );
AND2x2_ASAP7_75t_L g590 ( .A(n_516), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_SL g594 ( .A(n_517), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_517), .B(n_600), .Y(n_630) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_527), .Y(n_517) );
AND2x2_ASAP7_75t_L g555 ( .A(n_518), .B(n_528), .Y(n_555) );
INVx4_ASAP7_75t_L g567 ( .A(n_518), .Y(n_567) );
BUFx3_ASAP7_75t_L g610 ( .A(n_518), .Y(n_610) );
AND3x2_ASAP7_75t_L g625 ( .A(n_518), .B(n_626), .C(n_627), .Y(n_625) );
AND2x2_ASAP7_75t_L g707 ( .A(n_527), .B(n_621), .Y(n_707) );
AND2x2_ASAP7_75t_L g715 ( .A(n_527), .B(n_600), .Y(n_715) );
INVx1_ASAP7_75t_SL g720 ( .A(n_527), .Y(n_720) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_537), .Y(n_527) );
INVx1_ASAP7_75t_SL g578 ( .A(n_528), .Y(n_578) );
AND2x2_ASAP7_75t_L g601 ( .A(n_528), .B(n_567), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_528), .B(n_551), .Y(n_603) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_528), .Y(n_643) );
OR2x2_ASAP7_75t_L g648 ( .A(n_528), .B(n_567), .Y(n_648) );
INVx2_ASAP7_75t_L g553 ( .A(n_537), .Y(n_553) );
AND2x2_ASAP7_75t_L g588 ( .A(n_537), .B(n_568), .Y(n_588) );
OR2x2_ASAP7_75t_L g608 ( .A(n_537), .B(n_568), .Y(n_608) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_537), .Y(n_628) );
INVx1_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
AOI21xp33_ASAP7_75t_L g678 ( .A1(n_546), .A2(n_587), .B(n_679), .Y(n_678) );
AOI322xp5_ASAP7_75t_L g714 ( .A1(n_548), .A2(n_558), .A3(n_585), .B1(n_715), .B2(n_716), .C1(n_718), .C2(n_721), .Y(n_714) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_550), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_551), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g577 ( .A(n_552), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g645 ( .A(n_553), .B(n_567), .Y(n_645) );
AND2x2_ASAP7_75t_L g712 ( .A(n_553), .B(n_568), .Y(n_712) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g653 ( .A(n_555), .B(n_607), .Y(n_653) );
AOI31xp33_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_560), .A3(n_563), .B(n_564), .Y(n_556) );
AND2x2_ASAP7_75t_L g612 ( .A(n_558), .B(n_590), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_558), .B(n_582), .Y(n_694) );
AND2x2_ASAP7_75t_L g713 ( .A(n_558), .B(n_618), .Y(n_713) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_561), .B(n_590), .Y(n_602) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_561), .B(n_619), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_561), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_561), .B(n_703), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_562), .B(n_619), .Y(n_651) );
INVx1_ASAP7_75t_L g695 ( .A(n_562), .Y(n_695) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_577), .Y(n_565) );
INVxp67_ASAP7_75t_L g647 ( .A(n_566), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_567), .B(n_578), .Y(n_583) );
INVx1_ASAP7_75t_L g689 ( .A(n_567), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_567), .B(n_666), .Y(n_700) );
BUFx3_ASAP7_75t_L g600 ( .A(n_568), .Y(n_600) );
AND2x2_ASAP7_75t_L g626 ( .A(n_568), .B(n_578), .Y(n_626) );
INVx2_ASAP7_75t_L g666 ( .A(n_568), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_577), .B(n_699), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_584), .B(n_586), .C(n_595), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI21xp33_ASAP7_75t_L g629 ( .A1(n_581), .A2(n_630), .B(n_631), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_582), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_582), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g662 ( .A(n_583), .B(n_608), .Y(n_662) );
INVx3_ASAP7_75t_L g593 ( .A(n_585), .Y(n_593) );
OAI22xp5_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_589), .B1(n_592), .B2(n_594), .Y(n_586) );
OAI21xp5_ASAP7_75t_SL g611 ( .A1(n_588), .A2(n_612), .B(n_613), .Y(n_611) );
AND2x2_ASAP7_75t_L g637 ( .A(n_588), .B(n_601), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_588), .B(n_689), .Y(n_688) );
INVxp67_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g592 ( .A(n_591), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g661 ( .A(n_591), .Y(n_661) );
OAI21xp5_ASAP7_75t_SL g605 ( .A1(n_592), .A2(n_606), .B(n_611), .Y(n_605) );
OAI22xp33_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_598), .B1(n_602), .B2(n_603), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_597), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g621 ( .A(n_600), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_600), .B(n_643), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_616), .C(n_629), .Y(n_604) );
OAI22xp5_ASAP7_75t_SL g671 ( .A1(n_606), .A2(n_672), .B1(n_676), .B2(n_677), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g676 ( .A(n_608), .B(n_609), .Y(n_676) );
AND2x2_ASAP7_75t_L g684 ( .A(n_609), .B(n_665), .Y(n_684) );
CKINVDCx16_ASAP7_75t_R g609 ( .A(n_610), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_SL g692 ( .A1(n_610), .A2(n_693), .B(n_694), .C(n_695), .Y(n_692) );
OR2x2_ASAP7_75t_L g719 ( .A(n_610), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
OAI21xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_620), .B(n_622), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_618), .A2(n_655), .B(n_656), .C(n_659), .Y(n_654) );
OAI21xp33_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_624), .B(n_625), .Y(n_622) );
AND2x2_ASAP7_75t_L g687 ( .A(n_626), .B(n_645), .Y(n_687) );
INVxp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g665 ( .A(n_628), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g670 ( .A(n_630), .Y(n_670) );
NAND3xp33_ASAP7_75t_SL g633 ( .A(n_634), .B(n_654), .C(n_667), .Y(n_633) );
AOI211xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .B(n_638), .C(n_646), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
INVx1_ASAP7_75t_L g704 ( .A(n_641), .Y(n_704) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g664 ( .A(n_643), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_643), .B(n_712), .Y(n_711) );
INVxp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B(n_649), .C(n_650), .Y(n_646) );
INVx2_ASAP7_75t_SL g658 ( .A(n_648), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_649), .A2(n_660), .B1(n_662), .B2(n_663), .Y(n_659) );
OAI21xp33_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_652), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
AOI211xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .B(n_671), .C(n_678), .Y(n_667) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVxp33_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g721 ( .A(n_675), .Y(n_721) );
NAND4xp25_ASAP7_75t_L g680 ( .A(n_681), .B(n_696), .C(n_709), .D(n_714), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B(n_685), .C(n_692), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B(n_690), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g705 ( .A1(n_686), .A2(n_706), .B(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_693), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_713), .Y(n_709) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g736 ( .A(n_722), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_724), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g732 ( .A(n_726), .Y(n_732) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx3_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
endmodule