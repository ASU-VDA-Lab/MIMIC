module fake_jpeg_15747_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_66),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_68),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_69),
.A2(n_51),
.B1(n_42),
.B2(n_53),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_60),
.B1(n_56),
.B2(n_50),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_75),
.B1(n_79),
.B2(n_82),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_56),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_76),
.B(n_83),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_60),
.B1(n_48),
.B2(n_55),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_45),
.B1(n_58),
.B2(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_2),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_88),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_57),
.B1(n_4),
.B2(n_3),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_88)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_90),
.Y(n_96)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_99),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_86),
.B1(n_87),
.B2(n_91),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_94),
.B1(n_83),
.B2(n_95),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_97),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_104),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_98),
.B1(n_94),
.B2(n_100),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_106),
.B(n_77),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_107),
.A2(n_108),
.B1(n_78),
.B2(n_15),
.Y(n_109)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

NOR2xp67_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_14),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_111),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_78),
.C(n_29),
.Y(n_113)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g115 ( 
.A(n_114),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_25),
.B(n_30),
.Y(n_116)
);

OAI221xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.C(n_38),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_39),
.Y(n_118)
);


endmodule