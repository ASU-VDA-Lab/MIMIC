module fake_ariane_2644_n_207 (n_8, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_207);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_207;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_195;
wire n_110;
wire n_153;
wire n_197;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_205;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_174;
wire n_100;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_204;
wire n_200;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_84;
wire n_199;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_82;
wire n_178;
wire n_57;
wire n_131;
wire n_201;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_144;
wire n_130;
wire n_94;
wire n_101;
wire n_134;
wire n_188;
wire n_185;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_198;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_81;
wire n_87;
wire n_206;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_192;
wire n_80;
wire n_146;
wire n_194;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_78;
wire n_193;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_54;

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

INVxp67_ASAP7_75t_SL g64 ( 
.A(n_1),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_26),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g70 ( 
.A(n_8),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_16),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_29),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

OAI21x1_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_24),
.B(n_46),
.Y(n_86)
);

OA21x2_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_0),
.B(n_2),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

OA21x2_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_2),
.B(n_3),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_25),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_70),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_84),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_95),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_54),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_101),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

AND2x4_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_52),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

AO22x1_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_98),
.B1(n_100),
.B2(n_99),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_108),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_119),
.B(n_65),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_55),
.B1(n_83),
.B2(n_82),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_72),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_98),
.Y(n_137)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_63),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_80),
.Y(n_140)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_114),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_117),
.B(n_77),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_117),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_141),
.B(n_117),
.Y(n_149)
);

BUFx2_ASAP7_75t_SL g150 ( 
.A(n_123),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_3),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_4),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_138),
.B1(n_129),
.B2(n_134),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_74),
.B(n_79),
.C(n_78),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_76),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_81),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_81),
.B(n_5),
.Y(n_162)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_145),
.B(n_148),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_137),
.B(n_131),
.Y(n_164)
);

OAI21x1_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_143),
.B(n_139),
.Y(n_165)
);

AOI32xp33_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_136),
.A3(n_130),
.B1(n_122),
.B2(n_140),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

INVx4_ASAP7_75t_SL g168 ( 
.A(n_152),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_81),
.B1(n_10),
.B2(n_11),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

NOR2xp67_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_49),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_170),
.A2(n_155),
.B1(n_154),
.B2(n_146),
.Y(n_174)
);

INVx4_ASAP7_75t_SL g175 ( 
.A(n_167),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_160),
.B1(n_150),
.B2(n_159),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_157),
.B(n_147),
.C(n_161),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_15),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_165),
.B(n_164),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

AND2x4_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_171),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_169),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_173),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_163),
.Y(n_187)
);

INVx5_ASAP7_75t_SL g188 ( 
.A(n_182),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_28),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

OR2x6_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_32),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_33),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_190),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_192),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_198),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_191),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_194),
.B1(n_36),
.B2(n_37),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_42),
.B(n_43),
.Y(n_207)
);


endmodule