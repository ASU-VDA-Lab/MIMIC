module fake_jpeg_12386_n_615 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_615);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_615;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_483;
wire n_236;
wire n_291;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_312;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_63),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_64),
.Y(n_152)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_66),
.Y(n_164)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_67),
.Y(n_171)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_68),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_37),
.B(n_11),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_69),
.B(n_94),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_7),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_70),
.B(n_83),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_71),
.Y(n_162)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_72),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_73),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_50),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_74),
.B(n_115),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_77),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_81),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_82),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_20),
.B(n_7),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_88),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_89),
.Y(n_205)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_92),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_41),
.B(n_12),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_97),
.Y(n_186)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_98),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_41),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_105),
.Y(n_134)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_100),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_20),
.B(n_12),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_111),
.Y(n_141)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_26),
.B(n_12),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_107),
.Y(n_215)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_109),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_30),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_120),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_23),
.B(n_18),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_40),
.Y(n_112)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_113),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_23),
.B(n_6),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_114),
.B(n_117),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_31),
.B(n_6),
.Y(n_115)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_29),
.B(n_6),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_34),
.B(n_13),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_29),
.B(n_13),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_122),
.B(n_36),
.Y(n_211)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_31),
.Y(n_123)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_124),
.Y(n_210)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_38),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_127),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_38),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_128),
.Y(n_146)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_38),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_46),
.B1(n_42),
.B2(n_40),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_139),
.A2(n_148),
.B1(n_189),
.B2(n_212),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_77),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_140),
.B(n_142),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_45),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_42),
.B1(n_40),
.B2(n_34),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_45),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_150),
.B(n_154),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_116),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_80),
.B(n_51),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_158),
.B(n_179),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_53),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_159),
.B(n_168),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_112),
.A2(n_36),
.B1(n_46),
.B2(n_53),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_161),
.A2(n_177),
.B1(n_200),
.B2(n_160),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_119),
.A2(n_59),
.B(n_52),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g269 ( 
.A(n_167),
.B(n_3),
.CI(n_4),
.CON(n_269),
.SN(n_269)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_96),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_104),
.A2(n_52),
.B(n_32),
.C(n_44),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_170),
.A2(n_5),
.B(n_3),
.C(n_4),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_72),
.A2(n_100),
.B1(n_102),
.B2(n_90),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_106),
.B(n_51),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_107),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_183),
.B(n_188),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_126),
.B(n_55),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_91),
.A2(n_46),
.B1(n_42),
.B2(n_59),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_128),
.B(n_55),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_190),
.B(n_197),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_97),
.B(n_24),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_192),
.B(n_194),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_127),
.B(n_24),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_60),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_62),
.B(n_49),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_199),
.B(n_207),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_75),
.A2(n_47),
.B1(n_35),
.B2(n_50),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_64),
.A2(n_49),
.B1(n_47),
.B2(n_44),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_33),
.B1(n_88),
.B2(n_87),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_128),
.B(n_50),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_76),
.B(n_50),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_211),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_71),
.A2(n_47),
.B1(n_33),
.B2(n_32),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_203),
.A2(n_200),
.B1(n_170),
.B2(n_198),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_216),
.A2(n_231),
.B1(n_277),
.B2(n_160),
.Y(n_317)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_167),
.A2(n_109),
.B1(n_103),
.B2(n_93),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_219),
.A2(n_225),
.B1(n_230),
.B2(n_243),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_133),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_220),
.Y(n_334)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_221),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_222),
.A2(n_261),
.B1(n_289),
.B2(n_232),
.Y(n_305)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_223),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_224),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_212),
.A2(n_89),
.B1(n_82),
.B2(n_79),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_175),
.Y(n_226)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_226),
.Y(n_316)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_227),
.Y(n_322)
);

AO22x1_ASAP7_75t_SL g228 ( 
.A1(n_164),
.A2(n_78),
.B1(n_73),
.B2(n_30),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_228),
.B(n_272),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_166),
.Y(n_229)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_189),
.A2(n_30),
.B1(n_13),
.B2(n_14),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_30),
.B1(n_14),
.B2(n_15),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_182),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_233),
.B(n_246),
.Y(n_292)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_234),
.Y(n_291)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_235),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_146),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_236),
.B(n_266),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_238),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_0),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_239),
.B(n_252),
.C(n_259),
.Y(n_326)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_242),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_139),
.A2(n_30),
.B1(n_18),
.B2(n_17),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_143),
.A2(n_18),
.B1(n_16),
.B2(n_15),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_244),
.A2(n_245),
.B1(n_254),
.B2(n_262),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_143),
.A2(n_16),
.B1(n_15),
.B2(n_2),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_135),
.Y(n_246)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_248),
.Y(n_308)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_166),
.Y(n_249)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_249),
.Y(n_320)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_180),
.Y(n_250)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_250),
.Y(n_323)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_251),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_0),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_186),
.Y(n_253)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_253),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_143),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_147),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_255),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_130),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_256),
.A2(n_263),
.B1(n_205),
.B2(n_204),
.Y(n_333)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_163),
.Y(n_257)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_257),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_163),
.Y(n_258)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_258),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_164),
.B(n_0),
.Y(n_259)
);

NOR2x1_ASAP7_75t_L g347 ( 
.A(n_260),
.B(n_269),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_138),
.A2(n_141),
.B1(n_134),
.B2(n_169),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_178),
.A2(n_184),
.B1(n_156),
.B2(n_187),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_130),
.A2(n_201),
.B1(n_181),
.B2(n_178),
.Y(n_263)
);

BUFx4f_ASAP7_75t_SL g264 ( 
.A(n_196),
.Y(n_264)
);

INVx13_ASAP7_75t_L g329 ( 
.A(n_264),
.Y(n_329)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_132),
.Y(n_265)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_265),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_165),
.Y(n_266)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_132),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_274),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_269),
.A2(n_174),
.B(n_209),
.Y(n_310)
);

BUFx4f_ASAP7_75t_L g270 ( 
.A(n_187),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_270),
.Y(n_300)
);

AO22x1_ASAP7_75t_SL g272 ( 
.A1(n_169),
.A2(n_4),
.B1(n_5),
.B2(n_172),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_186),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_147),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_275),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_165),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_278),
.Y(n_302)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_191),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_145),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_280),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_145),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_129),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_281),
.B(n_136),
.Y(n_327)
);

BUFx12f_ASAP7_75t_L g282 ( 
.A(n_196),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_285),
.Y(n_314)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_153),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_283),
.Y(n_340)
);

BUFx2_ASAP7_75t_SL g284 ( 
.A(n_153),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_284),
.Y(n_341)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_157),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_172),
.B(n_4),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_287),
.B(n_131),
.C(n_152),
.Y(n_338)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_191),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_155),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_247),
.A2(n_214),
.B1(n_151),
.B2(n_193),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_296),
.A2(n_299),
.B1(n_313),
.B2(n_330),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_247),
.A2(n_214),
.B1(n_151),
.B2(n_193),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_305),
.A2(n_317),
.B1(n_240),
.B2(n_286),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_232),
.B(n_144),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_309),
.B(n_346),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_310),
.A2(n_311),
.B(n_347),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_260),
.A2(n_157),
.B(n_155),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_289),
.A2(n_202),
.B1(n_162),
.B2(n_137),
.Y(n_313)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_319),
.Y(n_351)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_327),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_288),
.A2(n_219),
.B1(n_218),
.B2(n_222),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_219),
.A2(n_202),
.B1(n_162),
.B2(n_137),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_331),
.A2(n_348),
.B1(n_227),
.B2(n_237),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_261),
.B(n_185),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_343),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_218),
.A2(n_185),
.B1(n_136),
.B2(n_195),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_337),
.A2(n_282),
.B1(n_280),
.B2(n_266),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_252),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_259),
.B(n_195),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_239),
.B(n_131),
.C(n_152),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_345),
.B(n_331),
.C(n_348),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_273),
.B(n_149),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_219),
.A2(n_149),
.B1(n_205),
.B2(n_204),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_361),
.Y(n_395)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_329),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_352),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_317),
.A2(n_304),
.B1(n_305),
.B2(n_315),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_353),
.A2(n_354),
.B1(n_368),
.B2(n_385),
.Y(n_413)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_324),
.Y(n_357)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_357),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_269),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_359),
.B(n_364),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_330),
.A2(n_252),
.B1(n_239),
.B2(n_287),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_360),
.A2(n_378),
.B(n_339),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_362),
.A2(n_370),
.B1(n_371),
.B2(n_388),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_311),
.B(n_259),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_309),
.B(n_271),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_365),
.B(n_372),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_339),
.Y(n_366)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_366),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_295),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_367),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_304),
.A2(n_228),
.B1(n_272),
.B2(n_267),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_308),
.Y(n_369)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_296),
.A2(n_228),
.B1(n_287),
.B2(n_272),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_299),
.A2(n_281),
.B1(n_238),
.B2(n_221),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_310),
.B(n_241),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

INVx6_ASAP7_75t_L g425 ( 
.A(n_373),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_290),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_380),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_326),
.B(n_265),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_376),
.B(n_377),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_326),
.B(n_250),
.C(n_274),
.Y(n_377)
);

MAJx2_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_253),
.C(n_278),
.Y(n_378)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_294),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_379),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_268),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_292),
.B(n_307),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_390),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_382),
.A2(n_341),
.B(n_300),
.Y(n_406)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_324),
.Y(n_383)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_383),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_347),
.B(n_327),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_393),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_347),
.A2(n_248),
.B1(n_224),
.B2(n_257),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_308),
.Y(n_386)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_293),
.A2(n_279),
.B1(n_258),
.B2(n_285),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_387),
.A2(n_392),
.B1(n_341),
.B2(n_300),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_313),
.A2(n_249),
.B1(n_234),
.B2(n_270),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_323),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_389),
.Y(n_422)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_294),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_307),
.B(n_283),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_340),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_293),
.A2(n_282),
.B1(n_229),
.B2(n_270),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_302),
.B(n_264),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_355),
.A2(n_361),
.B1(n_370),
.B2(n_364),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_400),
.A2(n_408),
.B1(n_416),
.B2(n_427),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_401),
.B(n_380),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_359),
.A2(n_314),
.B(n_303),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_339),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_405),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_406),
.B(n_306),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_393),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_407),
.B(n_409),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_355),
.A2(n_316),
.B1(n_321),
.B2(n_325),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_352),
.Y(n_412)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_412),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_356),
.B(n_350),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_424),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_358),
.A2(n_316),
.B1(n_321),
.B2(n_325),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_374),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_423),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_420),
.A2(n_362),
.B1(n_388),
.B2(n_375),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_369),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_356),
.B(n_318),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_384),
.A2(n_340),
.B(n_318),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_426),
.A2(n_430),
.B(n_329),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_358),
.A2(n_328),
.B1(n_322),
.B2(n_298),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_363),
.B(n_298),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_428),
.B(n_335),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_353),
.A2(n_329),
.B(n_332),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_395),
.B(n_376),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_432),
.B(n_442),
.C(n_448),
.Y(n_493)
);

OAI32xp33_ASAP7_75t_L g433 ( 
.A1(n_403),
.A2(n_350),
.A3(n_368),
.B1(n_351),
.B2(n_385),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_433),
.B(n_401),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_395),
.B(n_349),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_435),
.B(n_445),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_424),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_443),
.Y(n_472)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_394),
.Y(n_439)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_439),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_441),
.A2(n_451),
.B1(n_408),
.B2(n_405),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_395),
.B(n_377),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_409),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_SL g447 ( 
.A(n_396),
.B(n_403),
.C(n_428),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_447),
.A2(n_455),
.B(n_461),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_360),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_400),
.A2(n_375),
.B1(n_392),
.B2(n_351),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_449),
.A2(n_430),
.B1(n_410),
.B2(n_420),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_419),
.B(n_378),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_450),
.B(n_431),
.C(n_421),
.Y(n_496)
);

OAI22x1_ASAP7_75t_SL g451 ( 
.A1(n_413),
.A2(n_371),
.B1(n_383),
.B2(n_357),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_394),
.Y(n_452)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_452),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_419),
.B(n_328),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_453),
.B(n_402),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_416),
.A2(n_373),
.B1(n_306),
.B2(n_320),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_411),
.Y(n_456)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_456),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_457),
.A2(n_397),
.B(n_421),
.Y(n_495)
);

AO22x1_ASAP7_75t_SL g458 ( 
.A1(n_426),
.A2(n_344),
.B1(n_332),
.B2(n_389),
.Y(n_458)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_458),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_398),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_459),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_398),
.Y(n_460)
);

INVxp33_ASAP7_75t_SL g467 ( 
.A(n_460),
.Y(n_467)
);

A2O1A1O1Ixp25_ASAP7_75t_L g461 ( 
.A1(n_396),
.A2(n_344),
.B(n_342),
.C(n_334),
.D(n_264),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_415),
.B(n_386),
.Y(n_462)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_463),
.A2(n_405),
.B(n_420),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_417),
.B(n_301),
.Y(n_464)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_464),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_465),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_404),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_466),
.B(n_486),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_457),
.B(n_410),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_468),
.A2(n_481),
.B(n_495),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_444),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_469),
.B(n_431),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_440),
.A2(n_413),
.B1(n_430),
.B2(n_407),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_471),
.A2(n_478),
.B1(n_483),
.B2(n_434),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_474),
.B(n_487),
.Y(n_512)
);

OAI22x1_ASAP7_75t_L g481 ( 
.A1(n_449),
.A2(n_427),
.B1(n_406),
.B2(n_399),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_482),
.A2(n_463),
.B(n_446),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_440),
.A2(n_402),
.B1(n_414),
.B2(n_399),
.Y(n_483)
);

OAI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_484),
.A2(n_461),
.B1(n_438),
.B2(n_412),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_439),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_436),
.B(n_411),
.Y(n_488)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_488),
.Y(n_499)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_464),
.Y(n_491)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_491),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_451),
.A2(n_405),
.B1(n_423),
.B2(n_425),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_492),
.A2(n_455),
.B1(n_458),
.B2(n_456),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_436),
.B(n_397),
.Y(n_494)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_494),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_448),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_454),
.Y(n_497)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_497),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_498),
.A2(n_484),
.B1(n_492),
.B2(n_485),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_500),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_468),
.A2(n_434),
.B(n_446),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_501),
.B(n_507),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_466),
.B(n_432),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_502),
.B(n_510),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_475),
.C(n_435),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_505),
.B(n_509),
.C(n_521),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_472),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_450),
.C(n_453),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_496),
.B(n_445),
.Y(n_510)
);

XOR2x1_ASAP7_75t_L g511 ( 
.A(n_474),
.B(n_447),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_511),
.B(n_513),
.Y(n_524)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_494),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_514),
.B(n_518),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_486),
.B(n_462),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_471),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_475),
.B(n_483),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_516),
.B(n_522),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_517),
.A2(n_478),
.B1(n_479),
.B2(n_468),
.Y(n_528)
);

CKINVDCx14_ASAP7_75t_R g519 ( 
.A(n_488),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_519),
.A2(n_523),
.B1(n_479),
.B2(n_489),
.Y(n_530)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_470),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_520),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_458),
.C(n_463),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_489),
.B(n_433),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_526),
.B(n_531),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_528),
.A2(n_530),
.B1(n_541),
.B2(n_498),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_502),
.B(n_473),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_505),
.B(n_510),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_536),
.B(n_540),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_537),
.A2(n_412),
.B1(n_425),
.B2(n_418),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_516),
.B(n_481),
.C(n_467),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_538),
.B(n_539),
.C(n_543),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_513),
.B(n_509),
.C(n_508),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_508),
.B(n_482),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_522),
.A2(n_490),
.B1(n_499),
.B2(n_517),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_511),
.B(n_491),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_542),
.B(n_504),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_515),
.B(n_485),
.C(n_480),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_501),
.B(n_512),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_544),
.B(n_504),
.Y(n_559)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_529),
.Y(n_546)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_546),
.Y(n_571)
);

XNOR2x1_ASAP7_75t_L g574 ( 
.A(n_548),
.B(n_557),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_532),
.A2(n_497),
.B1(n_490),
.B2(n_512),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_549),
.B(n_550),
.Y(n_566)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_545),
.Y(n_550)
);

OAI221xp5_ASAP7_75t_L g551 ( 
.A1(n_525),
.A2(n_499),
.B1(n_514),
.B2(n_506),
.C(n_503),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_551),
.B(n_555),
.Y(n_570)
);

FAx1_ASAP7_75t_SL g554 ( 
.A(n_542),
.B(n_521),
.CI(n_506),
.CON(n_554),
.SN(n_554)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_554),
.B(n_560),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_528),
.A2(n_503),
.B1(n_480),
.B2(n_520),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_538),
.A2(n_487),
.B1(n_470),
.B2(n_477),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_556),
.B(n_558),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_535),
.A2(n_477),
.B1(n_476),
.B2(n_500),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_559),
.B(n_562),
.Y(n_575)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_543),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_533),
.B(n_438),
.C(n_476),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_561),
.B(n_563),
.C(n_533),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_527),
.B(n_342),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_562),
.A2(n_535),
.B(n_527),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_564),
.B(n_576),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_565),
.B(n_553),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_561),
.B(n_534),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_568),
.B(n_573),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_559),
.A2(n_534),
.B(n_524),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_569),
.A2(n_572),
.B1(n_547),
.B2(n_418),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_557),
.A2(n_540),
.B(n_539),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_563),
.B(n_536),
.C(n_320),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_551),
.A2(n_554),
.B(n_560),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_554),
.A2(n_418),
.B(n_422),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_578),
.B(n_546),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_579),
.B(n_580),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_566),
.A2(n_552),
.B1(n_550),
.B2(n_553),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_582),
.B(n_583),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_577),
.B(n_552),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_567),
.B(n_429),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_584),
.B(n_585),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_564),
.B(n_547),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_570),
.B(n_425),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_588),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_587),
.B(n_574),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_565),
.B(n_422),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_573),
.B(n_322),
.C(n_291),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_590),
.B(n_575),
.C(n_571),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_589),
.A2(n_576),
.B(n_578),
.Y(n_592)
);

AOI21xp33_ASAP7_75t_L g605 ( 
.A1(n_592),
.A2(n_594),
.B(n_312),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_589),
.A2(n_572),
.B(n_569),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_596),
.B(n_597),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g599 ( 
.A1(n_580),
.A2(n_574),
.B(n_575),
.Y(n_599)
);

AOI21x1_ASAP7_75t_L g602 ( 
.A1(n_599),
.A2(n_590),
.B(n_291),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_SL g600 ( 
.A1(n_593),
.A2(n_581),
.B(n_582),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_600),
.B(n_312),
.Y(n_609)
);

BUFx24_ASAP7_75t_SL g601 ( 
.A(n_595),
.Y(n_601)
);

AOI31xp33_ASAP7_75t_L g607 ( 
.A1(n_601),
.A2(n_604),
.A3(n_605),
.B(n_596),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_602),
.A2(n_591),
.B1(n_598),
.B2(n_297),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_598),
.B(n_422),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_606),
.Y(n_610)
);

INVxp33_ASAP7_75t_L g611 ( 
.A(n_607),
.Y(n_611)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_603),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_L g612 ( 
.A(n_611),
.B(n_609),
.C(n_608),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_612),
.B(n_610),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_613),
.A2(n_312),
.B1(n_322),
.B2(n_297),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_614),
.A2(n_323),
.B(n_335),
.Y(n_615)
);


endmodule