module fake_jpeg_13510_n_237 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx2_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_56),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_57),
.Y(n_73)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_28),
.Y(n_95)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_59),
.B(n_63),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_61),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_37),
.Y(n_91)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_0),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_33),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_19),
.C(n_20),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_6),
.C(n_7),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_62),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_20),
.B1(n_22),
.B2(n_34),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_80),
.A2(n_94),
.B1(n_12),
.B2(n_13),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_22),
.B1(n_35),
.B2(n_34),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_59),
.B1(n_41),
.B2(n_54),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_57),
.B(n_29),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_92),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_91),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_27),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_50),
.A2(n_35),
.B1(n_28),
.B2(n_37),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_63),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_42),
.B(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_97),
.B(n_102),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_52),
.B1(n_40),
.B2(n_45),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_98),
.A2(n_112),
.B1(n_77),
.B2(n_65),
.Y(n_140)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_10),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_105),
.B(n_111),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_114),
.B(n_117),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_43),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_1),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_67),
.B(n_14),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_13),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_118),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_54),
.B(n_3),
.C(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_1),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_125),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_66),
.A2(n_7),
.B(n_8),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_10),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_8),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_122),
.C(n_87),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_74),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_88),
.B1(n_75),
.B2(n_78),
.Y(n_143)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_80),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_135),
.Y(n_153)
);

AND2x4_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_74),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_117),
.B(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_90),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_137),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_66),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_142),
.B1(n_122),
.B2(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_141),
.B(n_143),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_75),
.B1(n_65),
.B2(n_78),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_72),
.B1(n_88),
.B2(n_89),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_145),
.A2(n_71),
.B1(n_110),
.B2(n_106),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_71),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_119),
.B1(n_125),
.B2(n_121),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_103),
.C(n_99),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_164),
.C(n_167),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_114),
.B(n_134),
.C(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_161),
.B1(n_162),
.B2(n_166),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_101),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_159),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_170),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_101),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_112),
.B1(n_96),
.B2(n_106),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_71),
.B1(n_100),
.B2(n_143),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_163),
.B(n_127),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_136),
.C(n_130),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_145),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_142),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_130),
.B1(n_147),
.B2(n_134),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_128),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_126),
.C(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_168),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_173),
.B(n_175),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_176),
.B(n_167),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_127),
.C(n_133),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_178),
.C(n_152),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_133),
.C(n_128),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_183),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_126),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_160),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_184),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_190),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_171),
.A2(n_150),
.B1(n_165),
.B2(n_160),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_192),
.B(n_174),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_193),
.B(n_176),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_179),
.B(n_177),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_197),
.Y(n_203)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_199),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_162),
.B1(n_155),
.B2(n_161),
.Y(n_200)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_181),
.B(n_182),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_185),
.B1(n_210),
.B2(n_202),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_182),
.B(n_174),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_192),
.C(n_201),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_201),
.C(n_190),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_209),
.A2(n_187),
.B(n_188),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_193),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_213),
.B(n_214),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_188),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_217),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_200),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_180),
.C(n_185),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_195),
.B1(n_207),
.B2(n_209),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_222),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_225),
.A2(n_216),
.B(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_229),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_223),
.B(n_224),
.Y(n_228)
);

AOI21x1_ASAP7_75t_L g232 ( 
.A1(n_228),
.A2(n_191),
.B(n_158),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_170),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_212),
.C(n_211),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_230),
.A2(n_220),
.B(n_180),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_231),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_233),
.C(n_226),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_230),
.B(n_156),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_235),
.Y(n_237)
);


endmodule