module real_aes_6970_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_314;
wire n_252;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g274 ( .A1(n_0), .A2(n_275), .B(n_276), .C(n_279), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_1), .B(n_263), .Y(n_280) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_3), .B(n_191), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_4), .A2(n_152), .B(n_155), .C(n_535), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_5), .A2(n_147), .B(n_559), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_6), .A2(n_147), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_7), .B(n_263), .Y(n_565) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_8), .A2(n_182), .B(n_219), .Y(n_218) );
AND2x6_ASAP7_75t_L g152 ( .A(n_9), .B(n_153), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_10), .A2(n_152), .B(n_155), .C(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g503 ( .A(n_11), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_12), .B(n_116), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_12), .B(n_40), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_13), .B(n_239), .Y(n_537) );
INVx1_ASAP7_75t_L g173 ( .A(n_14), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_15), .B(n_191), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_16), .A2(n_192), .B(n_521), .C(n_523), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_17), .B(n_263), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_18), .B(n_167), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_19), .A2(n_155), .B(n_158), .C(n_166), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_20), .A2(n_227), .B(n_278), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_21), .B(n_239), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_22), .A2(n_54), .B1(n_758), .B2(n_759), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_22), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_23), .B(n_239), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g550 ( .A(n_24), .Y(n_550) );
INVx1_ASAP7_75t_L g475 ( .A(n_25), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_26), .A2(n_155), .B(n_166), .C(n_222), .Y(n_221) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_27), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_28), .Y(n_533) );
INVx1_ASAP7_75t_L g491 ( .A(n_29), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_30), .A2(n_147), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g150 ( .A(n_31), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_32), .A2(n_195), .B(n_204), .C(n_206), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_33), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_34), .A2(n_278), .B(n_562), .C(n_564), .Y(n_561) );
INVxp67_ASAP7_75t_L g492 ( .A(n_35), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_36), .B(n_224), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_37), .A2(n_155), .B(n_166), .C(n_474), .Y(n_473) );
CKINVDCx14_ASAP7_75t_R g560 ( .A(n_38), .Y(n_560) );
AOI222xp33_ASAP7_75t_SL g129 ( .A1(n_39), .A2(n_130), .B1(n_136), .B2(n_742), .C1(n_743), .C2(n_747), .Y(n_129) );
INVx1_ASAP7_75t_L g116 ( .A(n_40), .Y(n_116) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_41), .A2(n_279), .B(n_501), .C(n_502), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_42), .B(n_146), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_43), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_44), .B(n_191), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_45), .B(n_147), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_46), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_47), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_48), .A2(n_195), .B(n_204), .C(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g277 ( .A(n_49), .Y(n_277) );
OAI22xp5_ASAP7_75t_SL g755 ( .A1(n_50), .A2(n_756), .B1(n_757), .B2(n_760), .Y(n_755) );
CKINVDCx16_ASAP7_75t_R g760 ( .A(n_50), .Y(n_760) );
INVx1_ASAP7_75t_L g249 ( .A(n_51), .Y(n_249) );
INVx1_ASAP7_75t_L g509 ( .A(n_52), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_53), .B(n_147), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_54), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_55), .Y(n_175) );
CKINVDCx14_ASAP7_75t_R g499 ( .A(n_56), .Y(n_499) );
INVx1_ASAP7_75t_L g153 ( .A(n_57), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_58), .B(n_147), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_59), .B(n_263), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_60), .A2(n_165), .B(n_188), .C(n_260), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_61), .Y(n_128) );
INVx1_ASAP7_75t_L g172 ( .A(n_62), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_63), .A2(n_102), .B1(n_132), .B2(n_133), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_63), .Y(n_133) );
INVx1_ASAP7_75t_SL g563 ( .A(n_64), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_65), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_66), .B(n_191), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_67), .B(n_263), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_68), .B(n_192), .Y(n_237) );
INVx1_ASAP7_75t_L g553 ( .A(n_69), .Y(n_553) );
CKINVDCx16_ASAP7_75t_R g273 ( .A(n_70), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_71), .B(n_160), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_72), .A2(n_155), .B(n_186), .C(n_195), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_73), .Y(n_258) );
INVx1_ASAP7_75t_L g113 ( .A(n_74), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_75), .A2(n_147), .B(n_498), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_76), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_77), .A2(n_147), .B(n_518), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_78), .A2(n_146), .B(n_487), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g472 ( .A(n_79), .Y(n_472) );
INVx1_ASAP7_75t_L g519 ( .A(n_80), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_81), .B(n_163), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_82), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_83), .A2(n_147), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g522 ( .A(n_84), .Y(n_522) );
INVx2_ASAP7_75t_L g170 ( .A(n_85), .Y(n_170) );
INVx1_ASAP7_75t_L g536 ( .A(n_86), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_87), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_88), .B(n_239), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_89), .A2(n_104), .B1(n_117), .B2(n_762), .Y(n_103) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_90), .B(n_110), .C(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g124 ( .A(n_90), .B(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g464 ( .A(n_90), .B(n_126), .Y(n_464) );
INVx2_ASAP7_75t_L g741 ( .A(n_90), .Y(n_741) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_91), .A2(n_131), .B1(n_134), .B2(n_135), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_91), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_92), .A2(n_155), .B(n_195), .C(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_93), .B(n_147), .Y(n_202) );
INVx1_ASAP7_75t_L g207 ( .A(n_94), .Y(n_207) );
INVxp67_ASAP7_75t_L g261 ( .A(n_95), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_96), .B(n_182), .Y(n_504) );
INVx2_ASAP7_75t_L g512 ( .A(n_97), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_98), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g187 ( .A(n_99), .Y(n_187) );
INVx1_ASAP7_75t_L g233 ( .A(n_100), .Y(n_233) );
AND2x2_ASAP7_75t_L g251 ( .A(n_101), .B(n_169), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_102), .Y(n_132) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_SL g763 ( .A(n_107), .Y(n_763) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_114), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g126 ( .A(n_110), .B(n_127), .Y(n_126) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI22x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_129), .B1(n_750), .B2(n_752), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_122), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g751 ( .A(n_121), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_122), .A2(n_753), .B(n_761), .Y(n_752) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_128), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx2_ASAP7_75t_L g761 ( .A(n_124), .Y(n_761) );
NOR2x2_ASAP7_75t_L g749 ( .A(n_125), .B(n_741), .Y(n_749) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g740 ( .A(n_126), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_130), .Y(n_742) );
INVx1_ASAP7_75t_L g134 ( .A(n_131), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_462), .B1(n_465), .B2(n_738), .Y(n_136) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_137), .A2(n_745), .B1(n_754), .B2(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx2_ASAP7_75t_L g745 ( .A(n_138), .Y(n_745) );
AND3x1_ASAP7_75t_L g138 ( .A(n_139), .B(n_366), .C(n_423), .Y(n_138) );
NOR3xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_311), .C(n_347), .Y(n_139) );
OAI211xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_213), .B(n_265), .C(n_298), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_177), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g268 ( .A(n_143), .B(n_269), .Y(n_268) );
INVx5_ASAP7_75t_L g297 ( .A(n_143), .Y(n_297) );
AND2x2_ASAP7_75t_L g370 ( .A(n_143), .B(n_286), .Y(n_370) );
AND2x2_ASAP7_75t_L g408 ( .A(n_143), .B(n_314), .Y(n_408) );
AND2x2_ASAP7_75t_L g428 ( .A(n_143), .B(n_270), .Y(n_428) );
OR2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_174), .Y(n_143) );
AOI21xp5_ASAP7_75t_SL g144 ( .A1(n_145), .A2(n_154), .B(n_167), .Y(n_144) );
BUFx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_148), .B(n_152), .Y(n_234) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx1_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
INVx1_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_151), .Y(n_161) );
INVx3_ASAP7_75t_L g192 ( .A(n_151), .Y(n_192) );
INVx1_ASAP7_75t_L g224 ( .A(n_151), .Y(n_224) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_151), .Y(n_239) );
BUFx3_ASAP7_75t_L g166 ( .A(n_152), .Y(n_166) );
INVx4_ASAP7_75t_SL g196 ( .A(n_152), .Y(n_196) );
INVx5_ASAP7_75t_L g205 ( .A(n_155), .Y(n_205) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_156), .Y(n_194) );
BUFx3_ASAP7_75t_L g210 ( .A(n_156), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_162), .B(n_164), .Y(n_158) );
INVx2_ASAP7_75t_L g163 ( .A(n_160), .Y(n_163) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx4_ASAP7_75t_L g189 ( .A(n_161), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_163), .A2(n_207), .B(n_208), .C(n_209), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_163), .A2(n_209), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp5_ASAP7_75t_L g535 ( .A1(n_163), .A2(n_536), .B(n_537), .C(n_538), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g552 ( .A1(n_163), .A2(n_538), .B(n_553), .C(n_554), .Y(n_552) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_164), .A2(n_191), .B(n_475), .C(n_476), .Y(n_474) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_165), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_168), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g176 ( .A(n_169), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_169), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_169), .A2(n_246), .B(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_169), .A2(n_234), .B(n_472), .C(n_473), .Y(n_471) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_169), .A2(n_497), .B(n_504), .Y(n_496) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_170), .B(n_171), .Y(n_169) );
AND2x2_ASAP7_75t_L g183 ( .A(n_170), .B(n_171), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_176), .A2(n_532), .B(n_539), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_177), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_200), .Y(n_177) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_178), .Y(n_309) );
AND2x2_ASAP7_75t_L g323 ( .A(n_178), .B(n_269), .Y(n_323) );
INVx1_ASAP7_75t_L g346 ( .A(n_178), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_178), .B(n_297), .Y(n_385) );
OR2x2_ASAP7_75t_L g422 ( .A(n_178), .B(n_267), .Y(n_422) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_179), .Y(n_358) );
AND2x2_ASAP7_75t_L g365 ( .A(n_179), .B(n_270), .Y(n_365) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g286 ( .A(n_180), .B(n_270), .Y(n_286) );
BUFx2_ASAP7_75t_L g314 ( .A(n_180), .Y(n_314) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_184), .B(n_198), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_181), .B(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_181), .B(n_212), .Y(n_211) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_181), .A2(n_232), .B(n_240), .Y(n_231) );
INVx3_ASAP7_75t_L g263 ( .A(n_181), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_181), .B(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_181), .B(n_540), .Y(n_539) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_181), .A2(n_549), .B(n_555), .Y(n_548) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_182), .A2(n_220), .B(n_221), .Y(n_219) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_182), .Y(n_255) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g242 ( .A(n_183), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_185), .B(n_197), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_190), .C(n_193), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g490 ( .A1(n_189), .A2(n_191), .B1(n_491), .B2(n_492), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_189), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_189), .B(n_522), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_191), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g275 ( .A(n_191), .Y(n_275) );
INVx5_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_192), .B(n_503), .Y(n_502) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g564 ( .A(n_194), .Y(n_564) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_196), .A2(n_205), .B(n_258), .C(n_259), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_SL g272 ( .A1(n_196), .A2(n_205), .B(n_273), .C(n_274), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_SL g487 ( .A1(n_196), .A2(n_205), .B(n_488), .C(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_SL g498 ( .A1(n_196), .A2(n_205), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_SL g508 ( .A1(n_196), .A2(n_205), .B(n_509), .C(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_196), .A2(n_205), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_196), .A2(n_205), .B(n_560), .C(n_561), .Y(n_559) );
INVx5_ASAP7_75t_L g267 ( .A(n_200), .Y(n_267) );
BUFx2_ASAP7_75t_L g290 ( .A(n_200), .Y(n_290) );
AND2x2_ASAP7_75t_L g447 ( .A(n_200), .B(n_301), .Y(n_447) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g279 ( .A(n_210), .Y(n_279) );
INVx1_ASAP7_75t_L g523 ( .A(n_210), .Y(n_523) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp33_ASAP7_75t_L g214 ( .A(n_215), .B(n_252), .Y(n_214) );
OAI221xp5_ASAP7_75t_L g347 ( .A1(n_215), .A2(n_348), .B1(n_355), .B2(n_356), .C(n_359), .Y(n_347) );
OR2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_229), .Y(n_215) );
AND2x2_ASAP7_75t_L g253 ( .A(n_216), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_216), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g282 ( .A(n_217), .B(n_230), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_217), .B(n_231), .Y(n_292) );
OR2x2_ASAP7_75t_L g303 ( .A(n_217), .B(n_254), .Y(n_303) );
AND2x2_ASAP7_75t_L g306 ( .A(n_217), .B(n_294), .Y(n_306) );
AND2x2_ASAP7_75t_L g322 ( .A(n_217), .B(n_243), .Y(n_322) );
OR2x2_ASAP7_75t_L g338 ( .A(n_217), .B(n_231), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_217), .B(n_254), .Y(n_400) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_218), .B(n_243), .Y(n_392) );
AND2x2_ASAP7_75t_L g395 ( .A(n_218), .B(n_231), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_225), .B(n_226), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_226), .A2(n_237), .B(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g316 ( .A(n_229), .B(n_303), .Y(n_316) );
INVx2_ASAP7_75t_L g342 ( .A(n_229), .Y(n_342) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_243), .Y(n_229) );
AND2x2_ASAP7_75t_L g264 ( .A(n_230), .B(n_244), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_230), .B(n_254), .Y(n_321) );
OR2x2_ASAP7_75t_L g332 ( .A(n_230), .B(n_244), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_230), .B(n_294), .Y(n_391) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_230), .A2(n_425), .B1(n_427), .B2(n_429), .C(n_432), .Y(n_424) );
INVx5_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_231), .B(n_254), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_235), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_234), .A2(n_533), .B(n_534), .Y(n_532) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_234), .A2(n_550), .B(n_551), .Y(n_549) );
INVx4_ASAP7_75t_L g278 ( .A(n_239), .Y(n_278) );
INVx2_ASAP7_75t_L g501 ( .A(n_239), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g484 ( .A(n_242), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_243), .B(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_243), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g310 ( .A(n_243), .B(n_282), .Y(n_310) );
OR2x2_ASAP7_75t_L g354 ( .A(n_243), .B(n_254), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_243), .B(n_306), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_243), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g419 ( .A(n_243), .B(n_420), .Y(n_419) );
INVx5_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_SL g283 ( .A(n_244), .B(n_253), .Y(n_283) );
O2A1O1Ixp33_ASAP7_75t_SL g287 ( .A1(n_244), .A2(n_288), .B(n_291), .C(n_295), .Y(n_287) );
OR2x2_ASAP7_75t_L g325 ( .A(n_244), .B(n_321), .Y(n_325) );
OR2x2_ASAP7_75t_L g361 ( .A(n_244), .B(n_303), .Y(n_361) );
OAI311xp33_ASAP7_75t_L g367 ( .A1(n_244), .A2(n_306), .A3(n_368), .B1(n_371), .C1(n_378), .Y(n_367) );
AND2x2_ASAP7_75t_L g418 ( .A(n_244), .B(n_254), .Y(n_418) );
AND2x2_ASAP7_75t_L g426 ( .A(n_244), .B(n_281), .Y(n_426) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_244), .Y(n_444) );
AND2x2_ASAP7_75t_L g461 ( .A(n_244), .B(n_282), .Y(n_461) );
OR2x6_ASAP7_75t_L g244 ( .A(n_245), .B(n_251), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_264), .Y(n_252) );
AND2x2_ASAP7_75t_L g289 ( .A(n_253), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g445 ( .A(n_253), .Y(n_445) );
AND2x2_ASAP7_75t_L g281 ( .A(n_254), .B(n_282), .Y(n_281) );
INVx3_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_254), .Y(n_337) );
INVxp67_ASAP7_75t_L g376 ( .A(n_254), .Y(n_376) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_262), .Y(n_254) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_255), .A2(n_507), .B(n_513), .Y(n_506) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_255), .A2(n_517), .B(n_524), .Y(n_516) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_255), .A2(n_558), .B(n_565), .Y(n_557) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_263), .A2(n_271), .B(n_280), .Y(n_270) );
AND2x2_ASAP7_75t_L g454 ( .A(n_264), .B(n_302), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_281), .B1(n_283), .B2(n_284), .C(n_287), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_267), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g307 ( .A(n_267), .B(n_297), .Y(n_307) );
AND2x2_ASAP7_75t_L g315 ( .A(n_267), .B(n_269), .Y(n_315) );
OR2x2_ASAP7_75t_L g327 ( .A(n_267), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g345 ( .A(n_267), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g369 ( .A(n_267), .B(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_267), .Y(n_389) );
AND2x2_ASAP7_75t_L g441 ( .A(n_267), .B(n_365), .Y(n_441) );
OAI31xp33_ASAP7_75t_L g449 ( .A1(n_267), .A2(n_318), .A3(n_417), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_268), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g413 ( .A(n_268), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_268), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g301 ( .A(n_269), .B(n_297), .Y(n_301) );
INVx1_ASAP7_75t_L g388 ( .A(n_269), .Y(n_388) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g438 ( .A(n_270), .B(n_297), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_278), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g538 ( .A(n_279), .Y(n_538) );
INVx1_ASAP7_75t_SL g448 ( .A(n_281), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_282), .B(n_353), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_283), .A2(n_395), .B1(n_433), .B2(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g296 ( .A(n_286), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g355 ( .A(n_286), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_286), .B(n_307), .Y(n_460) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g430 ( .A(n_289), .B(n_431), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_290), .A2(n_349), .B(n_351), .Y(n_348) );
OR2x2_ASAP7_75t_L g356 ( .A(n_290), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g377 ( .A(n_290), .B(n_365), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_290), .B(n_388), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_290), .B(n_428), .Y(n_427) );
OAI221xp5_ASAP7_75t_SL g404 ( .A1(n_291), .A2(n_405), .B1(n_410), .B2(n_413), .C(n_414), .Y(n_404) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
OR2x2_ASAP7_75t_L g381 ( .A(n_292), .B(n_354), .Y(n_381) );
INVx1_ASAP7_75t_L g420 ( .A(n_292), .Y(n_420) );
INVx2_ASAP7_75t_L g396 ( .A(n_293), .Y(n_396) );
INVx1_ASAP7_75t_L g330 ( .A(n_294), .Y(n_330) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g335 ( .A(n_297), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_297), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g364 ( .A(n_297), .B(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g452 ( .A(n_297), .B(n_422), .Y(n_452) );
AOI222xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B1(n_304), .B2(n_307), .C1(n_308), .C2(n_310), .Y(n_298) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g308 ( .A(n_301), .B(n_309), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_301), .A2(n_351), .B1(n_379), .B2(n_380), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_301), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OAI21xp33_ASAP7_75t_SL g339 ( .A1(n_310), .A2(n_340), .B(n_343), .Y(n_339) );
OAI211xp5_ASAP7_75t_SL g311 ( .A1(n_312), .A2(n_316), .B(n_317), .C(n_339), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_315), .A2(n_318), .B1(n_323), .B2(n_324), .C(n_326), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_315), .B(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g409 ( .A(n_315), .Y(n_409) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
AND2x2_ASAP7_75t_L g411 ( .A(n_320), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g328 ( .A(n_323), .Y(n_328) );
AND2x2_ASAP7_75t_L g334 ( .A(n_323), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_329), .B1(n_333), .B2(n_336), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_330), .B(n_342), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_331), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g431 ( .A(n_335), .Y(n_431) );
AND2x2_ASAP7_75t_L g450 ( .A(n_335), .B(n_365), .Y(n_450) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_342), .B(n_399), .Y(n_458) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_345), .B(n_413), .Y(n_456) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g379 ( .A(n_357), .Y(n_379) );
BUFx2_ASAP7_75t_L g403 ( .A(n_358), .Y(n_403) );
OAI21xp5_ASAP7_75t_SL g359 ( .A1(n_360), .A2(n_362), .B(n_364), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NOR3xp33_ASAP7_75t_L g366 ( .A(n_367), .B(n_382), .C(n_404), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_374), .B(n_377), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
A2O1A1Ixp33_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_386), .B(n_390), .C(n_393), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_383), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp67_ASAP7_75t_SL g387 ( .A(n_388), .B(n_389), .Y(n_387) );
OR2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_SL g412 ( .A(n_392), .Y(n_412) );
OAI21xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B(n_401), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
AND2x2_ASAP7_75t_L g417 ( .A(n_395), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_417), .B1(n_419), .B2(n_421), .Y(n_414) );
INVx2_ASAP7_75t_SL g435 ( .A(n_422), .Y(n_435) );
NOR3xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_439), .C(n_451), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_435), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_442), .B1(n_446), .B2(n_448), .C(n_449), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_440), .A2(n_452), .B(n_453), .C(n_455), .Y(n_451) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_459), .B2(n_461), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g744 ( .A(n_463), .Y(n_744) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_SL g746 ( .A(n_465), .Y(n_746) );
OR5x1_ASAP7_75t_L g465 ( .A(n_466), .B(n_632), .C(n_696), .D(n_712), .E(n_727), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_467), .B(n_566), .C(n_593), .D(n_616), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_514), .B(n_525), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_479), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx3_ASAP7_75t_SL g545 ( .A(n_470), .Y(n_545) );
AND2x4_ASAP7_75t_L g579 ( .A(n_470), .B(n_568), .Y(n_579) );
OR2x2_ASAP7_75t_L g589 ( .A(n_470), .B(n_547), .Y(n_589) );
OR2x2_ASAP7_75t_L g635 ( .A(n_470), .B(n_482), .Y(n_635) );
AND2x2_ASAP7_75t_L g649 ( .A(n_470), .B(n_546), .Y(n_649) );
AND2x2_ASAP7_75t_L g692 ( .A(n_470), .B(n_582), .Y(n_692) );
AND2x2_ASAP7_75t_L g699 ( .A(n_470), .B(n_557), .Y(n_699) );
AND2x2_ASAP7_75t_L g718 ( .A(n_470), .B(n_608), .Y(n_718) );
AND2x2_ASAP7_75t_L g736 ( .A(n_470), .B(n_578), .Y(n_736) );
OR2x6_ASAP7_75t_L g470 ( .A(n_471), .B(n_477), .Y(n_470) );
INVx1_ASAP7_75t_L g701 ( .A(n_479), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_495), .Y(n_479) );
AND2x2_ASAP7_75t_L g611 ( .A(n_480), .B(n_546), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_480), .B(n_631), .Y(n_630) );
AOI32xp33_ASAP7_75t_L g644 ( .A1(n_480), .A2(n_645), .A3(n_648), .B1(n_650), .B2(n_654), .Y(n_644) );
AND2x2_ASAP7_75t_L g714 ( .A(n_480), .B(n_608), .Y(n_714) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g578 ( .A(n_482), .B(n_547), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_482), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g620 ( .A(n_482), .B(n_567), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_482), .B(n_699), .Y(n_698) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_485), .B(n_493), .Y(n_482) );
INVx1_ASAP7_75t_L g583 ( .A(n_483), .Y(n_583) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OA21x2_ASAP7_75t_L g582 ( .A1(n_486), .A2(n_494), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g585 ( .A(n_495), .B(n_529), .Y(n_585) );
AND2x2_ASAP7_75t_L g661 ( .A(n_495), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g733 ( .A(n_495), .Y(n_733) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_505), .Y(n_495) );
OR2x2_ASAP7_75t_L g528 ( .A(n_496), .B(n_506), .Y(n_528) );
AND2x2_ASAP7_75t_L g542 ( .A(n_496), .B(n_543), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_496), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g592 ( .A(n_496), .Y(n_592) );
AND2x2_ASAP7_75t_L g619 ( .A(n_496), .B(n_506), .Y(n_619) );
BUFx3_ASAP7_75t_L g622 ( .A(n_496), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_496), .B(n_597), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_496), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g573 ( .A(n_505), .Y(n_573) );
AND2x2_ASAP7_75t_L g591 ( .A(n_505), .B(n_571), .Y(n_591) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g602 ( .A(n_506), .B(n_516), .Y(n_602) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_506), .Y(n_615) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_515), .B(n_622), .Y(n_672) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_SL g543 ( .A(n_516), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g590 ( .A(n_516), .B(n_591), .C(n_592), .Y(n_590) );
OR2x2_ASAP7_75t_L g598 ( .A(n_516), .B(n_571), .Y(n_598) );
AND2x2_ASAP7_75t_L g618 ( .A(n_516), .B(n_571), .Y(n_618) );
AND2x2_ASAP7_75t_L g662 ( .A(n_516), .B(n_531), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_541), .B(n_544), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_527), .B(n_529), .Y(n_526) );
AND2x2_ASAP7_75t_L g737 ( .A(n_527), .B(n_662), .Y(n_737) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_528), .A2(n_635), .B1(n_677), .B2(n_679), .Y(n_676) );
OR2x2_ASAP7_75t_L g683 ( .A(n_528), .B(n_598), .Y(n_683) );
OR2x2_ASAP7_75t_L g707 ( .A(n_528), .B(n_708), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_528), .B(n_627), .Y(n_720) );
AND2x2_ASAP7_75t_L g613 ( .A(n_529), .B(n_614), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_529), .A2(n_686), .B(n_701), .Y(n_700) );
AOI32xp33_ASAP7_75t_L g721 ( .A1(n_529), .A2(n_611), .A3(n_722), .B1(n_724), .B2(n_725), .Y(n_721) );
OR2x2_ASAP7_75t_L g732 ( .A(n_529), .B(n_733), .Y(n_732) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g600 ( .A(n_530), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_530), .B(n_614), .Y(n_679) );
BUFx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx4_ASAP7_75t_L g571 ( .A(n_531), .Y(n_571) );
AND2x2_ASAP7_75t_L g637 ( .A(n_531), .B(n_602), .Y(n_637) );
AND3x2_ASAP7_75t_L g646 ( .A(n_531), .B(n_542), .C(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g572 ( .A(n_543), .B(n_573), .Y(n_572) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_543), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_543), .B(n_571), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
AND2x2_ASAP7_75t_L g567 ( .A(n_545), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g607 ( .A(n_545), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g625 ( .A(n_545), .B(n_557), .Y(n_625) );
AND2x2_ASAP7_75t_L g643 ( .A(n_545), .B(n_547), .Y(n_643) );
OR2x2_ASAP7_75t_L g657 ( .A(n_545), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g703 ( .A(n_545), .B(n_631), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_546), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_557), .Y(n_546) );
AND2x2_ASAP7_75t_L g604 ( .A(n_547), .B(n_582), .Y(n_604) );
OR2x2_ASAP7_75t_L g658 ( .A(n_547), .B(n_582), .Y(n_658) );
AND2x2_ASAP7_75t_L g711 ( .A(n_547), .B(n_568), .Y(n_711) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
BUFx2_ASAP7_75t_L g609 ( .A(n_548), .Y(n_609) );
AND2x2_ASAP7_75t_L g631 ( .A(n_548), .B(n_557), .Y(n_631) );
INVx2_ASAP7_75t_L g568 ( .A(n_557), .Y(n_568) );
INVx1_ASAP7_75t_L g588 ( .A(n_557), .Y(n_588) );
AOI211xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_569), .B(n_574), .C(n_586), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_567), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g730 ( .A(n_567), .Y(n_730) );
AND2x2_ASAP7_75t_L g608 ( .A(n_568), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_571), .B(n_572), .Y(n_580) );
INVx1_ASAP7_75t_L g665 ( .A(n_571), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_571), .B(n_592), .Y(n_689) );
AND2x2_ASAP7_75t_L g705 ( .A(n_571), .B(n_619), .Y(n_705) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_572), .B(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g596 ( .A(n_573), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_580), .B1(n_581), .B2(n_584), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_577), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_578), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g603 ( .A(n_579), .B(n_604), .Y(n_603) );
AOI221xp5_ASAP7_75t_SL g668 ( .A1(n_579), .A2(n_621), .B1(n_669), .B2(n_674), .C(n_676), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_579), .B(n_642), .Y(n_675) );
INVx1_ASAP7_75t_L g735 ( .A(n_581), .Y(n_735) );
BUFx3_ASAP7_75t_L g642 ( .A(n_582), .Y(n_642) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI21xp33_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_589), .B(n_590), .Y(n_586) );
INVx1_ASAP7_75t_L g651 ( .A(n_588), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_588), .B(n_642), .Y(n_695) );
INVx1_ASAP7_75t_L g652 ( .A(n_589), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_589), .B(n_642), .Y(n_653) );
INVxp67_ASAP7_75t_L g673 ( .A(n_591), .Y(n_673) );
AND2x2_ASAP7_75t_L g614 ( .A(n_592), .B(n_615), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_599), .B(n_603), .C(n_605), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_SL g628 ( .A(n_596), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_597), .B(n_628), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_597), .B(n_619), .Y(n_670) );
INVx2_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_600), .A2(n_606), .B1(n_610), .B2(n_612), .Y(n_605) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g621 ( .A(n_602), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g666 ( .A(n_602), .B(n_667), .Y(n_666) );
OAI21xp33_ASAP7_75t_L g669 ( .A1(n_604), .A2(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_608), .A2(n_617), .B1(n_620), .B2(n_621), .C(n_623), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_608), .B(n_642), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_608), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g724 ( .A(n_614), .Y(n_724) );
INVxp67_ASAP7_75t_L g647 ( .A(n_615), .Y(n_647) );
INVx1_ASAP7_75t_L g654 ( .A(n_617), .Y(n_654) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AND2x2_ASAP7_75t_L g693 ( .A(n_618), .B(n_622), .Y(n_693) );
INVx1_ASAP7_75t_L g667 ( .A(n_622), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_622), .B(n_637), .Y(n_697) );
OAI32xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .A3(n_628), .B1(n_629), .B2(n_630), .Y(n_623) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_SL g636 ( .A(n_631), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_631), .B(n_663), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_631), .B(n_692), .Y(n_723) );
NAND2x1p5_ASAP7_75t_L g731 ( .A(n_631), .B(n_642), .Y(n_731) );
NAND5xp2_ASAP7_75t_L g632 ( .A(n_633), .B(n_655), .C(n_668), .D(n_680), .E(n_681), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_637), .B1(n_638), .B2(n_640), .C(n_644), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp33_ASAP7_75t_SL g659 ( .A(n_639), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_642), .B(n_711), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_643), .A2(n_656), .B1(n_659), .B2(n_663), .Y(n_655) );
INVx2_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
OAI211xp5_ASAP7_75t_SL g650 ( .A1(n_646), .A2(n_651), .B(n_652), .C(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g678 ( .A(n_658), .Y(n_678) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_667), .B(n_716), .Y(n_726) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B1(n_686), .B2(n_690), .C1(n_693), .C2(n_694), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI221xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B1(n_700), .B2(n_702), .C(n_704), .Y(n_696) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
OAI21xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B(n_709), .Y(n_704) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g716 ( .A(n_708), .Y(n_716) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B1(n_717), .B2(n_719), .C(n_721), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_731), .B(n_732), .C(n_734), .Y(n_727) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI21xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B(n_737), .Y(n_734) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_740), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
BUFx4f_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
endmodule