module fake_jpeg_18506_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_43),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_56),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_25),
.B1(n_20),
.B2(n_21),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_37),
.B1(n_38),
.B2(n_36),
.Y(n_78)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_37),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_26),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_68),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_77),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_81),
.Y(n_111)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_37),
.B1(n_25),
.B2(n_21),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_78),
.B1(n_91),
.B2(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_42),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_37),
.B(n_41),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_37),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_22),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_59),
.B(n_22),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_88),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_35),
.C(n_38),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_39),
.C(n_38),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_25),
.B1(n_20),
.B2(n_30),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_93),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_95),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_41),
.B1(n_20),
.B2(n_35),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_45),
.B1(n_41),
.B2(n_64),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_75),
.B1(n_71),
.B2(n_81),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_35),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_107),
.C(n_39),
.Y(n_133)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_44),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_38),
.C(n_39),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_69),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_109),
.B(n_114),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

XNOR2x1_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_40),
.Y(n_113)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_113),
.B(n_79),
.CI(n_40),
.CON(n_127),
.SN(n_127)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_63),
.B(n_73),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_124),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_69),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_109),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_30),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_105),
.B1(n_106),
.B2(n_117),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_127),
.A2(n_136),
.B(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_66),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_132),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_87),
.B(n_91),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_151),
.B(n_105),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_83),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_88),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_137),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_74),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_95),
.B1(n_96),
.B2(n_84),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_135),
.A2(n_139),
.B1(n_140),
.B2(n_98),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_44),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_40),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_148),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_70),
.B1(n_41),
.B2(n_82),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_70),
.B1(n_41),
.B2(n_67),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_65),
.B1(n_45),
.B2(n_64),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_144),
.B1(n_149),
.B2(n_150),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_44),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_76),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_147),
.B(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_40),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_119),
.A2(n_76),
.B1(n_40),
.B2(n_80),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_119),
.A2(n_40),
.B1(n_80),
.B2(n_44),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_112),
.A2(n_33),
.B(n_16),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_44),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_89),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_107),
.C(n_104),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_185),
.C(n_127),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_158),
.A2(n_176),
.B(n_180),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_170),
.B1(n_182),
.B2(n_186),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_103),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_166),
.B(n_173),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_116),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_189),
.Y(n_208)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_118),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_184),
.Y(n_190)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_106),
.B(n_116),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_117),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_177),
.B(n_178),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_138),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_143),
.B1(n_136),
.B2(n_126),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_181),
.B1(n_32),
.B2(n_34),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_97),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_124),
.B1(n_97),
.B2(n_98),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_135),
.A2(n_121),
.B1(n_110),
.B2(n_122),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_121),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_123),
.C(n_69),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_129),
.A2(n_110),
.B1(n_122),
.B2(n_16),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_132),
.B(n_80),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_152),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_197),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_210),
.C(n_185),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_156),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_127),
.B1(n_144),
.B2(n_150),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_200),
.A2(n_209),
.B1(n_215),
.B2(n_198),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_165),
.A2(n_151),
.B1(n_155),
.B2(n_33),
.Y(n_201)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_159),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_202),
.B(n_206),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_164),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_26),
.Y(n_207)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_182),
.B1(n_188),
.B2(n_165),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_108),
.C(n_155),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_160),
.B1(n_179),
.B2(n_157),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_18),
.Y(n_213)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_32),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_189),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_180),
.A2(n_10),
.B1(n_14),
.B2(n_12),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_175),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_18),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_162),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_219),
.A2(n_162),
.B(n_181),
.Y(n_222)
);

OA21x2_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_158),
.B(n_176),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_222),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_168),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_228),
.A2(n_233),
.B1(n_238),
.B2(n_215),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_236),
.C(n_237),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_197),
.B(n_10),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_204),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_198),
.B1(n_213),
.B2(n_218),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_160),
.B1(n_1),
.B2(n_2),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_31),
.C(n_24),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_31),
.C(n_24),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_195),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_31),
.C(n_24),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_200),
.C(n_194),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_209),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_241),
.B(n_192),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_205),
.A2(n_32),
.B(n_28),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_244),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_224),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_247),
.Y(n_267)
);

XOR2x2_ASAP7_75t_SL g247 ( 
.A(n_228),
.B(n_205),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_243),
.Y(n_248)
);

BUFx2_ASAP7_75t_SL g277 ( 
.A(n_248),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_251),
.C(n_260),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_214),
.C(n_216),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_190),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_261),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_238),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_255),
.A2(n_23),
.B1(n_18),
.B2(n_34),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_240),
.B1(n_220),
.B2(n_227),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_219),
.B1(n_190),
.B2(n_193),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_220),
.B1(n_242),
.B2(n_233),
.Y(n_266)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_207),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_216),
.C(n_193),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_237),
.C(n_234),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_226),
.A2(n_199),
.B1(n_217),
.B2(n_191),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_240),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_270),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_268),
.A2(n_261),
.B1(n_262),
.B2(n_23),
.Y(n_285)
);

OAI322xp33_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_239),
.A3(n_191),
.B1(n_227),
.B2(n_199),
.C1(n_32),
.C2(n_28),
.Y(n_271)
);

AOI21xp33_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_277),
.B(n_272),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_249),
.A2(n_7),
.B(n_11),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_9),
.B(n_8),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_252),
.B(n_7),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_278),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_254),
.Y(n_279)
);

NAND4xp25_ASAP7_75t_SL g293 ( 
.A(n_279),
.B(n_9),
.C(n_8),
.D(n_7),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_23),
.C(n_6),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_251),
.C(n_245),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_260),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_289),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_244),
.B1(n_250),
.B2(n_246),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_285),
.B1(n_276),
.B2(n_278),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_291),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_262),
.C(n_11),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_294),
.C(n_272),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_11),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_280),
.C(n_273),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_0),
.B(n_3),
.Y(n_304)
);

OA21x2_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_0),
.B(n_1),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_3),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_8),
.C(n_2),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_268),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_297),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_302),
.C(n_304),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_287),
.B(n_264),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_299),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_264),
.C(n_274),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_300),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_289),
.C(n_291),
.Y(n_309)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_309),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_298),
.A2(n_294),
.B1(n_286),
.B2(n_288),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_310),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_281),
.C(n_292),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_291),
.C(n_293),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_317),
.B(n_308),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_295),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_300),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_3),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_320),
.C(n_321),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_SL g321 ( 
.A1(n_316),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_314),
.B(n_4),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_323),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_4),
.B(n_5),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_5),
.Y(n_326)
);


endmodule