module real_jpeg_15448_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_465),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_0),
.B(n_466),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_1),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_1),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_1),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_1),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_1),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_1),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_1),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_1),
.B(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_2),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_2),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_3),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_3),
.Y(n_339)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_4),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_5),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_5),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_5),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_5),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_5),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_5),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_5),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_5),
.B(n_87),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_6),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_6),
.B(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_6),
.A2(n_11),
.B1(n_118),
.B2(n_121),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_6),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_6),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_6),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_6),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_7),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_7),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_7),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_7),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_7),
.B(n_360),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_7),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_7),
.B(n_412),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_8),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_8),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_8),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_8),
.B(n_146),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_8),
.B(n_120),
.Y(n_179)
);

NAND2x1p5_ASAP7_75t_L g191 ( 
.A(n_8),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_8),
.B(n_262),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_8),
.B(n_104),
.Y(n_295)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_9),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_9),
.Y(n_142)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_10),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_10),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_10),
.Y(n_224)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_10),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_11),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_11),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_11),
.B(n_100),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_11),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_11),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_11),
.B(n_442),
.Y(n_441)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_12),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_13),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_13),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_13),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_13),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_13),
.B(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_13),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_14),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_15),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_15),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_15),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_15),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_15),
.B(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_15),
.B(n_64),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_15),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_15),
.B(n_398),
.Y(n_416)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_16),
.Y(n_110)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_17),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g448 ( 
.A(n_17),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_R g19 ( 
.A1(n_20),
.A2(n_428),
.B1(n_463),
.B2(n_464),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_21),
.Y(n_463)
);

NAND2x1_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_319),
.Y(n_21)
);

A2O1A1O1Ixp25_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_232),
.B(n_281),
.C(n_282),
.D(n_318),
.Y(n_22)
);

OAI21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_203),
.B(n_231),
.Y(n_23)
);

NOR2x1_ASAP7_75t_L g320 ( 
.A(n_24),
.B(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_155),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_25),
.B(n_155),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_101),
.C(n_126),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_26),
.B(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_66),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_44),
.Y(n_27)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_28),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_40),
.B2(n_41),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_31),
.B(n_39),
.C(n_40),
.Y(n_181)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_33),
.Y(n_169)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_33),
.Y(n_457)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_37),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_40),
.A2(n_41),
.B1(n_314),
.B2(n_317),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_41),
.B(n_311),
.C(n_317),
.Y(n_459)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_44),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_55),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_46),
.A2(n_50),
.B(n_55),
.C(n_200),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_48),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_48),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_48),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_48),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_49),
.B(n_54),
.Y(n_200)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.C(n_63),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_56),
.A2(n_63),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_56),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_56),
.A2(n_99),
.B1(n_129),
.B2(n_215),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_59),
.B(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_61),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_63),
.B(n_270),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_66),
.B(n_157),
.C(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_82),
.C(n_92),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_67),
.B(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_74),
.C(n_78),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_76),
.Y(n_396)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_77),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_77),
.Y(n_342)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_77),
.Y(n_368)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_82),
.A2(n_83),
.B1(n_92),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_178),
.Y(n_216)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_88),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_89),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_89),
.Y(n_178)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_92),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.C(n_99),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_93),
.A2(n_99),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_93),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_95),
.B(n_213),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_98),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_99),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_99),
.A2(n_145),
.B1(n_215),
.B2(n_266),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_99),
.B(n_266),
.C(n_303),
.Y(n_460)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_100),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_100),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_101),
.B(n_126),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_114),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_102),
.B(n_116),
.C(n_125),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_103),
.B(n_107),
.C(n_111),
.Y(n_197)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_111),
.B2(n_113),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_109),
.Y(n_415)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_111),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_113),
.B(n_145),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_125),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_132),
.B(n_138),
.Y(n_131)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.C(n_143),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_127),
.B(n_131),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_130),
.B(n_271),
.C(n_278),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_133),
.B(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_133),
.B(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_143),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_151),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_144),
.B(n_332),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_145),
.A2(n_179),
.B1(n_180),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_145),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_145),
.B(n_180),
.C(n_261),
.Y(n_296)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_332)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_156),
.B(n_184),
.C(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_184),
.B2(n_185),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_161),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_173),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_162),
.B(n_181),
.C(n_182),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_163),
.B(n_168),
.C(n_170),
.Y(n_256)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_170),
.A2(n_439),
.B1(n_440),
.B2(n_441),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_170),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_172),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_173)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_175),
.B(n_178),
.C(n_180),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_179),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_179),
.B(n_341),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_180),
.B(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_197),
.B2(n_198),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_190)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_191),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_193),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_194),
.B(n_196),
.C(n_198),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_197),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_229),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_204),
.B(n_229),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.C(n_211),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_205),
.B(n_325),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_211),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.C(n_217),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_212),
.B(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_216),
.B(n_217),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.C(n_225),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_218),
.B(n_225),
.Y(n_375)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_222),
.B(n_375),
.Y(n_374)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND4xp25_ASAP7_75t_SL g319 ( 
.A(n_232),
.B(n_282),
.C(n_320),
.D(n_322),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_235),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_236),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.C(n_239),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_259),
.B1(n_279),
.B2(n_280),
.Y(n_240)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_258),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_242),
.B(n_245),
.C(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_257),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_247),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_256),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_252),
.C(n_256),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_253),
.B(n_298),
.C(n_451),
.Y(n_450)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_279),
.C(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_268),
.C(n_269),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_265),
.Y(n_260)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_278),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_285),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_286),
.B(n_288),
.C(n_300),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_300),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_299),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_289),
.B(n_292),
.C(n_293),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_291),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

AO22x1_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_293)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_294),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_295),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_296),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_308),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_301),
.B(n_309),
.C(n_310),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_304),
.B(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

OAI21x1_ASAP7_75t_SL g322 ( 
.A1(n_323),
.A2(n_343),
.B(n_427),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_324),
.B(n_327),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_331),
.C(n_333),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_328),
.A2(n_329),
.B1(n_424),
.B2(n_425),
.Y(n_423)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_331),
.B(n_333),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.C(n_340),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_334),
.A2(n_335),
.B1(n_336),
.B2(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_340),
.B(n_377),
.Y(n_376)
);

AOI21x1_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_421),
.B(n_426),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_379),
.B(n_420),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_371),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_346),
.B(n_371),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_362),
.C(n_369),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_347),
.A2(n_348),
.B1(n_387),
.B2(n_389),
.Y(n_386)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_358),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_355),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_355),
.C(n_358),
.Y(n_373)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_362),
.A2(n_369),
.B1(n_370),
.B2(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_362),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_363),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.Y(n_382)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_376),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_373),
.B(n_374),
.C(n_376),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_390),
.B(n_419),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_386),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_381),
.B(n_386),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.C(n_385),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_402),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_383),
.A2(n_384),
.B1(n_385),
.B2(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_385),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_387),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_391),
.A2(n_404),
.B(n_418),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_401),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_392),
.B(n_401),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_397),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_397),
.Y(n_409)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_410),
.B(n_417),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_406),
.B(n_409),
.Y(n_417)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_416),
.Y(n_410)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_422),
.B(n_423),
.Y(n_426)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_428),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_462),
.Y(n_428)
);

OR2x6_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_461),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_430),
.B(n_461),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_452),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_450),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_438),
.B1(n_445),
.B2(n_449),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_445),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_447),
.Y(n_446)
);

INVx8_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_458),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

INVx6_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);


endmodule