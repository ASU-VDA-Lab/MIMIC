module fake_jpeg_28035_n_250 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_16),
.B1(n_30),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_49),
.B1(n_50),
.B2(n_57),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_16),
.B1(n_30),
.B2(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_16),
.B1(n_30),
.B2(n_37),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_18),
.B(n_33),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_29),
.C(n_39),
.Y(n_67)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_56),
.B(n_15),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_29),
.B1(n_32),
.B2(n_31),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_64),
.B(n_66),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_22),
.Y(n_66)
);

HB1xp67_ASAP7_75t_SL g89 ( 
.A(n_67),
.Y(n_89)
);

OR2x4_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_43),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_75),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_81),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_71),
.B(n_73),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_24),
.A3(n_31),
.B1(n_21),
.B2(n_17),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_59),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_24),
.A3(n_31),
.B1(n_21),
.B2(n_17),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_26),
.B1(n_28),
.B2(n_51),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_17),
.B1(n_21),
.B2(n_24),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_79),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_23),
.B1(n_39),
.B2(n_33),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_48),
.B1(n_46),
.B2(n_51),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_13),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_23),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_27),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_73),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_96),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_58),
.B1(n_46),
.B2(n_48),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_101),
.B1(n_80),
.B2(n_81),
.Y(n_115)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_95),
.A2(n_93),
.B1(n_110),
.B2(n_97),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_40),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_40),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_59),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_74),
.B1(n_72),
.B2(n_65),
.Y(n_135)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_107),
.Y(n_126)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_69),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_51),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_118),
.B1(n_135),
.B2(n_112),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_68),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_109),
.Y(n_160)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_112),
.A2(n_83),
.B1(n_69),
.B2(n_74),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_28),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_127),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_124),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_62),
.C(n_40),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_131),
.C(n_62),
.Y(n_158)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_28),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_128),
.B(n_130),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_62),
.C(n_40),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_99),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_28),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_95),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_146),
.A2(n_148),
.B1(n_161),
.B2(n_42),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_105),
.B(n_89),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_147),
.A2(n_150),
.B(n_151),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_138),
.A2(n_92),
.B1(n_110),
.B2(n_93),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_132),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_154),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_102),
.B(n_106),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_109),
.B(n_102),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_124),
.B1(n_128),
.B2(n_130),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_123),
.B(n_119),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_1),
.B(n_2),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_156),
.A2(n_159),
.B1(n_33),
.B2(n_38),
.Y(n_173)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_115),
.A2(n_72),
.B1(n_65),
.B2(n_42),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_171),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_114),
.C(n_122),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_170),
.C(n_2),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_143),
.B(n_133),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_168),
.B(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_135),
.C(n_85),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_1),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_174),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_1),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_175),
.A2(n_176),
.B(n_181),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_38),
.Y(n_176)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_183),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_161),
.B1(n_148),
.B2(n_144),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_42),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_162),
.Y(n_183)
);

INVxp33_ASAP7_75t_SL g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_184),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_186),
.A2(n_194),
.B1(n_197),
.B2(n_190),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_144),
.B(n_140),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_189),
.A2(n_202),
.B(n_176),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_163),
.Y(n_193)
);

AO21x1_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_4),
.B(n_7),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_147),
.B1(n_145),
.B2(n_139),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_166),
.B(n_151),
.Y(n_195)
);

A2O1A1O1Ixp25_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_175),
.B(n_182),
.C(n_167),
.D(n_179),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_201),
.C(n_10),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_11),
.C(n_6),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_4),
.B(n_7),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_199),
.B1(n_186),
.B2(n_190),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_195),
.A2(n_178),
.B1(n_181),
.B2(n_170),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_213),
.B1(n_209),
.B2(n_215),
.Y(n_223)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_198),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_215),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_200),
.A2(n_171),
.B(n_164),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_210),
.B(n_187),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_165),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_201),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_189),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_176),
.B1(n_7),
.B2(n_8),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_209),
.A2(n_197),
.B1(n_194),
.B2(n_202),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_198),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_222),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_221),
.Y(n_227)
);

INVx11_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_225),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_208),
.C(n_207),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_226),
.A2(n_217),
.B(n_203),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_230),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_225),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_227),
.A2(n_224),
.B1(n_204),
.B2(n_206),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_237),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_220),
.B1(n_211),
.B2(n_221),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_222),
.C(n_188),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_232),
.C(n_228),
.Y(n_241)
);

NAND5xp2_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_185),
.C(n_188),
.D(n_212),
.E(n_187),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_234),
.B(n_237),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_238),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_239),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_245),
.B(n_246),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_229),
.B(n_192),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_240),
.B(n_213),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_11),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_11),
.Y(n_250)
);


endmodule