module fake_jpeg_16764_n_116 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_116);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_0),
.C(n_1),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_2),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_41),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_24),
.B1(n_25),
.B2(n_19),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_22),
.B1(n_20),
.B2(n_17),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_24),
.B1(n_19),
.B2(n_17),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_12),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_51),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_58),
.B1(n_61),
.B2(n_36),
.Y(n_72)
);

BUFx2_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_15),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_18),
.B(n_20),
.C(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_14),
.B(n_18),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_23),
.B(n_21),
.C(n_7),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_43),
.Y(n_64)
);

XNOR2x2_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_49),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_46),
.B1(n_37),
.B2(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_47),
.B1(n_21),
.B2(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_36),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_46),
.B1(n_37),
.B2(n_9),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_5),
.Y(n_83)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_80),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_62),
.C(n_61),
.Y(n_79)
);

A2O1A1O1Ixp25_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_74),
.B(n_67),
.C(n_60),
.D(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_82),
.B(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_84),
.B(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_64),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_66),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_71),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_76),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_81),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_70),
.B(n_67),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_93),
.B(n_89),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_55),
.B(n_48),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_88),
.B1(n_91),
.B2(n_83),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_6),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_98),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_99),
.B1(n_5),
.B2(n_6),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_45),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_104),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_96),
.B(n_10),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_100),
.A2(n_65),
.B1(n_56),
.B2(n_10),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_65),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_107),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_28),
.B(n_30),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_105),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_111),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_103),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_28),
.B(n_30),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_113),
.A2(n_110),
.B1(n_28),
.B2(n_30),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_114),
.Y(n_116)
);


endmodule