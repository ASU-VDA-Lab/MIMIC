module fake_aes_4408_n_1075 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1075);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1075;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_801;
wire n_988;
wire n_1059;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_1030;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_599;
wire n_724;
wire n_857;
wire n_786;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_624;
wire n_426;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_1018;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_459;
wire n_863;
wire n_322;
wire n_907;
wire n_708;
wire n_1062;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_935;
wire n_460;
wire n_1046;
wire n_478;
wire n_482;
wire n_415;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_501;
wire n_871;
wire n_803;
wire n_338;
wire n_519;
wire n_699;
wire n_805;
wire n_729;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_881;
wire n_806;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_591;
wire n_933;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_654;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_947;
wire n_912;
wire n_924;
wire n_1043;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_504;
wire n_581;
wire n_458;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_991;
wire n_515;
wire n_670;
wire n_843;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_695;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_606;
wire n_934;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_405;
wire n_772;
wire n_987;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
INVx1_ASAP7_75t_L g319 ( .A(n_145), .Y(n_319) );
INVx1_ASAP7_75t_SL g320 ( .A(n_125), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_202), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_108), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_120), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_243), .Y(n_324) );
CKINVDCx14_ASAP7_75t_R g325 ( .A(n_123), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_151), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_298), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_237), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_62), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_127), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_316), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_293), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_317), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_134), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_5), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_302), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_126), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_98), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_18), .Y(n_339) );
CKINVDCx14_ASAP7_75t_R g340 ( .A(n_2), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_30), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_205), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_306), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_130), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_112), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_20), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_187), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_95), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_111), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_242), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_56), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_158), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_285), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_305), .Y(n_354) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_157), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_147), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_281), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_8), .Y(n_358) );
BUFx10_ASAP7_75t_L g359 ( .A(n_60), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_303), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_297), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_165), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_32), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_194), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_96), .Y(n_365) );
NOR2xp67_ASAP7_75t_L g366 ( .A(n_160), .B(n_232), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_100), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_217), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_136), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_313), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_284), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_209), .Y(n_372) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_296), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_311), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_69), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_230), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_135), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_40), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_138), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_203), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_171), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_274), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_207), .Y(n_383) );
INVx1_ASAP7_75t_SL g384 ( .A(n_299), .Y(n_384) );
CKINVDCx16_ASAP7_75t_R g385 ( .A(n_201), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_291), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_211), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_39), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_124), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_220), .Y(n_390) );
BUFx8_ASAP7_75t_SL g391 ( .A(n_99), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_55), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_118), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_301), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_140), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_215), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_270), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_236), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_94), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_110), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_294), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_104), .Y(n_402) );
CKINVDCx14_ASAP7_75t_R g403 ( .A(n_79), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_290), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_44), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_77), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_188), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_5), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_88), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_252), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_141), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_65), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_300), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_286), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_97), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_289), .Y(n_416) );
INVx2_ASAP7_75t_SL g417 ( .A(n_318), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_164), .Y(n_418) );
BUFx10_ASAP7_75t_L g419 ( .A(n_307), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_73), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_304), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_15), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_206), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_287), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_101), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_27), .Y(n_426) );
BUFx10_ASAP7_75t_L g427 ( .A(n_10), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_156), .Y(n_428) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_189), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_260), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_161), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_10), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_224), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_128), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_49), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_292), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_310), .Y(n_437) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_288), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_42), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_131), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_76), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_295), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_66), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_137), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_20), .B(n_227), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_247), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_282), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_277), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_417), .Y(n_449) );
BUFx12f_ASAP7_75t_L g450 ( .A(n_427), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_337), .Y(n_451) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_344), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_345), .B(n_0), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_391), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_369), .Y(n_455) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_344), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_340), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_335), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_427), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_364), .B(n_0), .Y(n_460) );
INVx3_ASAP7_75t_L g461 ( .A(n_359), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_444), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_346), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_339), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_353), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_359), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_380), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_344), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_373), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_358), .Y(n_470) );
NOR2xp33_ASAP7_75t_R g471 ( .A(n_454), .B(n_325), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_465), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_457), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_450), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_457), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_463), .Y(n_476) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_453), .A2(n_323), .B(n_319), .Y(n_477) );
INVxp33_ASAP7_75t_SL g478 ( .A(n_458), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_463), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_470), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_470), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_459), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_449), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_458), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_459), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_466), .Y(n_486) );
NOR2xp67_ASAP7_75t_L g487 ( .A(n_461), .B(n_448), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_453), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_462), .A2(n_355), .B1(n_385), .B2(n_363), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_461), .Y(n_490) );
NOR2xp33_ASAP7_75t_SL g491 ( .A(n_478), .B(n_396), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_477), .B(n_460), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_484), .B(n_460), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_476), .B(n_408), .C(n_426), .Y(n_494) );
NOR2xp33_ASAP7_75t_SL g495 ( .A(n_479), .B(n_398), .Y(n_495) );
OAI21xp33_ASAP7_75t_L g496 ( .A1(n_483), .A2(n_455), .B(n_451), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_485), .B(n_321), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_482), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_482), .Y(n_499) );
NAND2xp33_ASAP7_75t_L g500 ( .A(n_471), .B(n_322), .Y(n_500) );
NAND2xp33_ASAP7_75t_SL g501 ( .A(n_488), .B(n_413), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_477), .Y(n_502) );
AND2x6_ASAP7_75t_L g503 ( .A(n_489), .B(n_327), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_480), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_486), .B(n_464), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_487), .B(n_481), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_490), .B(n_467), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_490), .B(n_419), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_474), .B(n_324), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_473), .B(n_419), .Y(n_510) );
INVxp33_ASAP7_75t_L g511 ( .A(n_475), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_472), .Y(n_512) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_482), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_483), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_477), .B(n_403), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_477), .B(n_328), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_489), .B(n_432), .C(n_341), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_502), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_514), .B(n_428), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_513), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_493), .A2(n_445), .B1(n_332), .B2(n_350), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_504), .Y(n_522) );
INVx5_ASAP7_75t_L g523 ( .A(n_513), .Y(n_523) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_513), .Y(n_524) );
INVxp67_ASAP7_75t_L g525 ( .A(n_491), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_496), .Y(n_526) );
OR2x2_ASAP7_75t_SL g527 ( .A(n_491), .B(n_422), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_501), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_492), .B(n_326), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_505), .B(n_330), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_499), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_506), .B(n_331), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_498), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_507), .B(n_333), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_516), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_516), .Y(n_536) );
INVx8_ASAP7_75t_L g537 ( .A(n_503), .Y(n_537) );
OAI22xp5_ASAP7_75t_SL g538 ( .A1(n_511), .A2(n_336), .B1(n_338), .B2(n_334), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_515), .Y(n_539) );
NAND2x1p5_ASAP7_75t_L g540 ( .A(n_512), .B(n_320), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_517), .B(n_342), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_495), .B(n_343), .Y(n_542) );
INVx5_ASAP7_75t_L g543 ( .A(n_503), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_508), .A2(n_354), .B1(n_356), .B2(n_329), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_510), .B(n_1), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_503), .B(n_347), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_497), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_535), .B(n_503), .Y(n_548) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_544), .A2(n_494), .B(n_500), .C(n_495), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_536), .A2(n_509), .B(n_362), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_522), .A2(n_370), .B1(n_371), .B2(n_361), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_518), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_529), .A2(n_378), .B(n_372), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_518), .A2(n_527), .B1(n_519), .B2(n_539), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_523), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_534), .A2(n_526), .B(n_531), .Y(n_556) );
CKINVDCx16_ASAP7_75t_R g557 ( .A(n_538), .Y(n_557) );
OAI22xp5_ASAP7_75t_SL g558 ( .A1(n_540), .A2(n_349), .B1(n_351), .B2(n_348), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_533), .A2(n_387), .B(n_386), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_521), .B(n_389), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_547), .B(n_393), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_543), .B(n_397), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_524), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_530), .A2(n_401), .B(n_399), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_541), .Y(n_565) );
CKINVDCx8_ASAP7_75t_R g566 ( .A(n_537), .Y(n_566) );
INVx3_ASAP7_75t_L g567 ( .A(n_523), .Y(n_567) );
O2A1O1Ixp5_ASAP7_75t_L g568 ( .A1(n_542), .A2(n_382), .B(n_394), .C(n_381), .Y(n_568) );
NAND2x1p5_ASAP7_75t_L g569 ( .A(n_523), .B(n_384), .Y(n_569) );
AOI22x1_ASAP7_75t_L g570 ( .A1(n_539), .A2(n_469), .B1(n_424), .B2(n_416), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_545), .A2(n_410), .B(n_412), .C(n_407), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_539), .A2(n_415), .B1(n_357), .B2(n_360), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_532), .A2(n_423), .B(n_414), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_520), .A2(n_439), .B(n_437), .Y(n_574) );
OAI22xp5_ASAP7_75t_SL g575 ( .A1(n_528), .A2(n_367), .B1(n_368), .B2(n_352), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_520), .A2(n_442), .B(n_441), .Y(n_576) );
NOR3xp33_ASAP7_75t_SL g577 ( .A(n_546), .B(n_375), .C(n_374), .Y(n_577) );
O2A1O1Ixp33_ASAP7_75t_L g578 ( .A1(n_525), .A2(n_447), .B(n_404), .C(n_365), .Y(n_578) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_543), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_543), .B(n_376), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_524), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_524), .A2(n_366), .B(n_379), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_537), .B(n_383), .Y(n_583) );
AOI22x1_ASAP7_75t_L g584 ( .A1(n_553), .A2(n_456), .B1(n_468), .B2(n_452), .Y(n_584) );
AOI21x1_ASAP7_75t_L g585 ( .A1(n_554), .A2(n_469), .B(n_456), .Y(n_585) );
NAND2x1p5_ASAP7_75t_L g586 ( .A(n_567), .B(n_373), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_552), .Y(n_587) );
BUFx3_ASAP7_75t_L g588 ( .A(n_567), .Y(n_588) );
AO21x2_ASAP7_75t_L g589 ( .A1(n_556), .A2(n_469), .B(n_456), .Y(n_589) );
AO21x2_ASAP7_75t_L g590 ( .A1(n_582), .A2(n_469), .B(n_468), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_565), .B(n_1), .Y(n_591) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_570), .A2(n_377), .B(n_373), .Y(n_592) );
BUFx3_ASAP7_75t_L g593 ( .A(n_566), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g594 ( .A1(n_564), .A2(n_390), .B(n_388), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_569), .Y(n_595) );
INVxp67_ASAP7_75t_SL g596 ( .A(n_581), .Y(n_596) );
INVx4_ASAP7_75t_L g597 ( .A(n_569), .Y(n_597) );
OAI21x1_ASAP7_75t_L g598 ( .A1(n_563), .A2(n_395), .B(n_377), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_548), .Y(n_599) );
BUFx6f_ASAP7_75t_SL g600 ( .A(n_557), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_561), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_562), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_571), .B(n_2), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_555), .Y(n_604) );
OAI21x1_ASAP7_75t_L g605 ( .A1(n_582), .A2(n_395), .B(n_377), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_579), .Y(n_606) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_580), .Y(n_607) );
AO21x2_ASAP7_75t_L g608 ( .A1(n_559), .A2(n_468), .B(n_452), .Y(n_608) );
OAI21x1_ASAP7_75t_L g609 ( .A1(n_568), .A2(n_429), .B(n_395), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_560), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_551), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_550), .Y(n_612) );
OAI21x1_ASAP7_75t_L g613 ( .A1(n_574), .A2(n_436), .B(n_429), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_549), .Y(n_614) );
BUFx2_ASAP7_75t_SL g615 ( .A(n_572), .Y(n_615) );
OAI21x1_ASAP7_75t_L g616 ( .A1(n_576), .A2(n_436), .B(n_429), .Y(n_616) );
BUFx4_ASAP7_75t_SL g617 ( .A(n_558), .Y(n_617) );
AO21x2_ASAP7_75t_L g618 ( .A1(n_578), .A2(n_452), .B(n_438), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_577), .B(n_3), .Y(n_619) );
OAI21x1_ASAP7_75t_L g620 ( .A1(n_573), .A2(n_438), .B(n_436), .Y(n_620) );
OAI21x1_ASAP7_75t_L g621 ( .A1(n_583), .A2(n_438), .B(n_34), .Y(n_621) );
AOI22x1_ASAP7_75t_L g622 ( .A1(n_575), .A2(n_400), .B1(n_402), .B2(n_392), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_552), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_567), .B(n_3), .Y(n_624) );
NAND2x1_ASAP7_75t_L g625 ( .A(n_552), .B(n_33), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_565), .A2(n_406), .B1(n_409), .B2(n_405), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_552), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_556), .A2(n_418), .B(n_411), .Y(n_628) );
INVxp67_ASAP7_75t_SL g629 ( .A(n_552), .Y(n_629) );
BUFx2_ASAP7_75t_L g630 ( .A(n_569), .Y(n_630) );
BUFx3_ASAP7_75t_L g631 ( .A(n_567), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_557), .B(n_4), .Y(n_632) );
AO21x2_ASAP7_75t_L g633 ( .A1(n_556), .A2(n_36), .B(n_35), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_552), .Y(n_634) );
AOI22x1_ASAP7_75t_L g635 ( .A1(n_553), .A2(n_421), .B1(n_425), .B2(n_420), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_552), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_636), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_623), .Y(n_638) );
AOI21x1_ASAP7_75t_L g639 ( .A1(n_585), .A2(n_431), .B(n_430), .Y(n_639) );
BUFx2_ASAP7_75t_R g640 ( .A(n_593), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_634), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_587), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_587), .Y(n_643) );
AOI21x1_ASAP7_75t_L g644 ( .A1(n_614), .A2(n_434), .B(n_433), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_629), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_623), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_611), .A2(n_440), .B1(n_443), .B2(n_435), .Y(n_647) );
BUFx8_ASAP7_75t_SL g648 ( .A(n_600), .Y(n_648) );
BUFx4f_ASAP7_75t_L g649 ( .A(n_624), .Y(n_649) );
AO21x2_ASAP7_75t_L g650 ( .A1(n_589), .A2(n_4), .B(n_6), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_591), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_627), .A2(n_446), .B1(n_8), .B2(n_6), .Y(n_652) );
AO21x1_ASAP7_75t_L g653 ( .A1(n_624), .A2(n_7), .B(n_9), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_630), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_627), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_597), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_629), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_610), .A2(n_11), .B1(n_7), .B2(n_9), .Y(n_658) );
NOR2x1_ASAP7_75t_SL g659 ( .A(n_597), .B(n_11), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_601), .A2(n_14), .B1(n_12), .B2(n_13), .Y(n_660) );
CKINVDCx11_ASAP7_75t_R g661 ( .A(n_606), .Y(n_661) );
INVx4_ASAP7_75t_SL g662 ( .A(n_600), .Y(n_662) );
CKINVDCx11_ASAP7_75t_R g663 ( .A(n_606), .Y(n_663) );
INVx4_ASAP7_75t_L g664 ( .A(n_588), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_586), .Y(n_665) );
BUFx4f_ASAP7_75t_SL g666 ( .A(n_631), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_586), .Y(n_667) );
INVx6_ASAP7_75t_L g668 ( .A(n_588), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_603), .A2(n_14), .B1(n_12), .B2(n_13), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_591), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_599), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_607), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_632), .A2(n_17), .B1(n_15), .B2(n_16), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_595), .B(n_16), .Y(n_674) );
BUFx4_ASAP7_75t_SL g675 ( .A(n_604), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_617), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_607), .Y(n_677) );
AO21x2_ASAP7_75t_L g678 ( .A1(n_589), .A2(n_17), .B(n_18), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_607), .Y(n_679) );
BUFx2_ASAP7_75t_L g680 ( .A(n_596), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_603), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_602), .A2(n_22), .B1(n_19), .B2(n_21), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g683 ( .A1(n_612), .A2(n_19), .B(n_21), .Y(n_683) );
BUFx10_ASAP7_75t_L g684 ( .A(n_619), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_615), .A2(n_24), .B1(n_22), .B2(n_23), .Y(n_685) );
INVx2_ASAP7_75t_SL g686 ( .A(n_617), .Y(n_686) );
BUFx3_ASAP7_75t_L g687 ( .A(n_619), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_607), .Y(n_688) );
INVx4_ASAP7_75t_L g689 ( .A(n_618), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_596), .B(n_23), .Y(n_690) );
OAI21x1_ASAP7_75t_L g691 ( .A1(n_598), .A2(n_38), .B(n_37), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_590), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_621), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_626), .B(n_24), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_590), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_605), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_609), .A2(n_43), .B(n_41), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_608), .Y(n_698) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_608), .Y(n_699) );
INVxp67_ASAP7_75t_L g700 ( .A(n_622), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_633), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_594), .A2(n_27), .B1(n_25), .B2(n_26), .Y(n_702) );
NAND2x1p5_ASAP7_75t_L g703 ( .A(n_625), .B(n_25), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_594), .A2(n_29), .B1(n_26), .B2(n_28), .Y(n_704) );
AOI22xp33_ASAP7_75t_SL g705 ( .A1(n_618), .A2(n_30), .B1(n_28), .B2(n_29), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_620), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_626), .B(n_31), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_633), .Y(n_708) );
INVx11_ASAP7_75t_L g709 ( .A(n_635), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_613), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_616), .Y(n_711) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_592), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_584), .Y(n_713) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_628), .Y(n_714) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_628), .A2(n_31), .B1(n_32), .B2(n_45), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_610), .B(n_315), .Y(n_716) );
BUFx2_ASAP7_75t_SL g717 ( .A(n_593), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_634), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_611), .A2(n_48), .B1(n_46), .B2(n_47), .Y(n_719) );
INVx2_ASAP7_75t_SL g720 ( .A(n_593), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_629), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_611), .A2(n_52), .B1(n_50), .B2(n_51), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_637), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g724 ( .A(n_686), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_638), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_645), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_646), .B(n_53), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_680), .Y(n_728) );
OAI21x1_ASAP7_75t_L g729 ( .A1(n_696), .A2(n_54), .B(n_57), .Y(n_729) );
NAND2xp33_ASAP7_75t_R g730 ( .A(n_676), .B(n_58), .Y(n_730) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_656), .Y(n_731) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_645), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_641), .Y(n_733) );
NAND2xp33_ASAP7_75t_SL g734 ( .A(n_664), .B(n_59), .Y(n_734) );
NOR2xp33_ASAP7_75t_R g735 ( .A(n_661), .B(n_61), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_649), .A2(n_63), .B1(n_64), .B2(n_67), .Y(n_736) );
NOR2xp33_ASAP7_75t_R g737 ( .A(n_663), .B(n_68), .Y(n_737) );
OAI21xp33_ASAP7_75t_L g738 ( .A1(n_687), .A2(n_70), .B(n_71), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_721), .Y(n_739) );
NOR2xp33_ASAP7_75t_R g740 ( .A(n_649), .B(n_72), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_721), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_666), .Y(n_742) );
AND2x4_ASAP7_75t_L g743 ( .A(n_664), .B(n_74), .Y(n_743) );
INVxp33_ASAP7_75t_L g744 ( .A(n_648), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_718), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_657), .Y(n_746) );
BUFx2_ASAP7_75t_L g747 ( .A(n_668), .Y(n_747) );
NAND2xp33_ASAP7_75t_R g748 ( .A(n_674), .B(n_75), .Y(n_748) );
NAND2xp33_ASAP7_75t_R g749 ( .A(n_674), .B(n_694), .Y(n_749) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_675), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_654), .B(n_314), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_690), .B(n_78), .Y(n_752) );
BUFx3_ASAP7_75t_L g753 ( .A(n_720), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_671), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_707), .B(n_80), .Y(n_755) );
INVxp33_ASAP7_75t_SL g756 ( .A(n_717), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_684), .B(n_640), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_671), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_642), .Y(n_759) );
INVx4_ASAP7_75t_L g760 ( .A(n_662), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_702), .A2(n_704), .B1(n_685), .B2(n_658), .Y(n_761) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_643), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_655), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_672), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_659), .B(n_81), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_684), .B(n_82), .Y(n_766) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_668), .Y(n_767) );
CKINVDCx16_ASAP7_75t_R g768 ( .A(n_662), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_651), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_677), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_682), .B(n_83), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_673), .A2(n_84), .B1(n_85), .B2(n_86), .Y(n_772) );
NAND2xp33_ASAP7_75t_R g773 ( .A(n_665), .B(n_87), .Y(n_773) );
NAND2x1p5_ASAP7_75t_L g774 ( .A(n_667), .B(n_89), .Y(n_774) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_709), .Y(n_775) );
CKINVDCx11_ASAP7_75t_R g776 ( .A(n_679), .Y(n_776) );
NAND3xp33_ASAP7_75t_SL g777 ( .A(n_653), .B(n_90), .C(n_91), .Y(n_777) );
AND2x2_ASAP7_75t_SL g778 ( .A(n_660), .B(n_92), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_670), .B(n_312), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_688), .Y(n_780) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_650), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_652), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_700), .B(n_93), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_681), .B(n_102), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_669), .B(n_103), .Y(n_785) );
NOR2xp33_ASAP7_75t_R g786 ( .A(n_644), .B(n_105), .Y(n_786) );
NOR3xp33_ASAP7_75t_SL g787 ( .A(n_715), .B(n_106), .C(n_107), .Y(n_787) );
OR2x6_ASAP7_75t_L g788 ( .A(n_703), .B(n_109), .Y(n_788) );
AO31x2_ASAP7_75t_L g789 ( .A1(n_701), .A2(n_113), .A3(n_114), .B(n_115), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_716), .B(n_116), .Y(n_790) );
NOR2x1_ASAP7_75t_L g791 ( .A(n_650), .B(n_117), .Y(n_791) );
CKINVDCx16_ASAP7_75t_R g792 ( .A(n_714), .Y(n_792) );
BUFx4f_ASAP7_75t_SL g793 ( .A(n_714), .Y(n_793) );
INVxp67_ASAP7_75t_L g794 ( .A(n_714), .Y(n_794) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_689), .Y(n_795) );
OA21x2_ASAP7_75t_L g796 ( .A1(n_701), .A2(n_119), .B(n_121), .Y(n_796) );
BUFx6f_ASAP7_75t_L g797 ( .A(n_689), .Y(n_797) );
OR2x6_ASAP7_75t_L g798 ( .A(n_691), .B(n_122), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_678), .Y(n_799) );
NOR3xp33_ASAP7_75t_SL g800 ( .A(n_683), .B(n_129), .C(n_132), .Y(n_800) );
AND2x4_ASAP7_75t_L g801 ( .A(n_678), .B(n_133), .Y(n_801) );
AND3x2_ASAP7_75t_L g802 ( .A(n_699), .B(n_139), .C(n_142), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_705), .B(n_647), .Y(n_803) );
BUFx6f_ASAP7_75t_L g804 ( .A(n_698), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_693), .Y(n_805) );
NOR2xp33_ASAP7_75t_R g806 ( .A(n_639), .B(n_143), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_692), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_708), .A2(n_144), .B1(n_146), .B2(n_148), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_692), .B(n_149), .Y(n_809) );
INVxp67_ASAP7_75t_R g810 ( .A(n_713), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_719), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_695), .Y(n_812) );
NAND2x1p5_ASAP7_75t_L g813 ( .A(n_710), .B(n_150), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_710), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_711), .Y(n_815) );
NAND2xp5_ASAP7_75t_SL g816 ( .A(n_722), .B(n_152), .Y(n_816) );
AOI21x1_ASAP7_75t_L g817 ( .A1(n_711), .A2(n_153), .B(n_154), .Y(n_817) );
NOR3xp33_ASAP7_75t_SL g818 ( .A(n_697), .B(n_155), .C(n_159), .Y(n_818) );
NAND2xp33_ASAP7_75t_R g819 ( .A(n_706), .B(n_162), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_712), .B(n_163), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_712), .Y(n_821) );
A2O1A1Ixp33_ASAP7_75t_L g822 ( .A1(n_712), .A2(n_166), .B(n_167), .C(n_168), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_637), .B(n_169), .Y(n_823) );
NOR3xp33_ASAP7_75t_SL g824 ( .A(n_676), .B(n_170), .C(n_172), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_637), .B(n_309), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_637), .B(n_173), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_637), .Y(n_827) );
AND2x4_ASAP7_75t_L g828 ( .A(n_664), .B(n_174), .Y(n_828) );
BUFx3_ASAP7_75t_L g829 ( .A(n_666), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_731), .B(n_175), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_728), .B(n_723), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_827), .B(n_176), .Y(n_832) );
AND2x4_ASAP7_75t_SL g833 ( .A(n_743), .B(n_177), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_725), .B(n_754), .Y(n_834) );
INVx11_ASAP7_75t_L g835 ( .A(n_756), .Y(n_835) );
OR2x2_ASAP7_75t_L g836 ( .A(n_732), .B(n_178), .Y(n_836) );
OR2x2_ASAP7_75t_L g837 ( .A(n_758), .B(n_179), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_726), .Y(n_838) );
INVx3_ASAP7_75t_L g839 ( .A(n_795), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_769), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_733), .B(n_180), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_745), .B(n_181), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_782), .B(n_182), .Y(n_843) );
NOR2xp67_ASAP7_75t_SL g844 ( .A(n_768), .B(n_183), .Y(n_844) );
BUFx3_ASAP7_75t_L g845 ( .A(n_747), .Y(n_845) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_762), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_739), .B(n_184), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_741), .Y(n_848) );
NOR2x1_ASAP7_75t_SL g849 ( .A(n_788), .B(n_185), .Y(n_849) );
OR2x2_ASAP7_75t_L g850 ( .A(n_746), .B(n_186), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_759), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_763), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_807), .B(n_190), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_805), .Y(n_854) );
BUFx3_ASAP7_75t_L g855 ( .A(n_776), .Y(n_855) );
BUFx2_ASAP7_75t_L g856 ( .A(n_767), .Y(n_856) );
BUFx2_ASAP7_75t_L g857 ( .A(n_743), .Y(n_857) );
AND2x4_ASAP7_75t_L g858 ( .A(n_760), .B(n_794), .Y(n_858) );
OAI21x1_ASAP7_75t_L g859 ( .A1(n_791), .A2(n_191), .B(n_192), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_814), .B(n_193), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_815), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_764), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_753), .B(n_195), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_770), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_780), .B(n_196), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_812), .Y(n_866) );
INVxp67_ASAP7_75t_SL g867 ( .A(n_804), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_799), .B(n_197), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_781), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_809), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_804), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_810), .B(n_198), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_792), .B(n_199), .Y(n_873) );
OR2x2_ASAP7_75t_L g874 ( .A(n_724), .B(n_200), .Y(n_874) );
BUFx2_ASAP7_75t_L g875 ( .A(n_828), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_804), .Y(n_876) );
AO21x2_ASAP7_75t_L g877 ( .A1(n_777), .A2(n_204), .B(n_208), .Y(n_877) );
AND2x4_ASAP7_75t_L g878 ( .A(n_795), .B(n_210), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_727), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_828), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_795), .Y(n_881) );
OR2x2_ASAP7_75t_L g882 ( .A(n_751), .B(n_212), .Y(n_882) );
INVx2_ASAP7_75t_L g883 ( .A(n_797), .Y(n_883) );
INVxp67_ASAP7_75t_L g884 ( .A(n_749), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_752), .B(n_213), .Y(n_885) );
OR2x2_ASAP7_75t_L g886 ( .A(n_742), .B(n_214), .Y(n_886) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_797), .Y(n_887) );
INVx2_ASAP7_75t_L g888 ( .A(n_797), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_761), .B(n_216), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_823), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_784), .B(n_218), .Y(n_891) );
BUFx2_ASAP7_75t_L g892 ( .A(n_740), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_811), .B(n_219), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_778), .A2(n_221), .B1(n_222), .B2(n_223), .Y(n_894) );
INVx2_ASAP7_75t_SL g895 ( .A(n_829), .Y(n_895) );
BUFx3_ASAP7_75t_L g896 ( .A(n_793), .Y(n_896) );
AND2x4_ASAP7_75t_L g897 ( .A(n_788), .B(n_225), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_821), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_820), .Y(n_899) );
AND2x4_ASAP7_75t_L g900 ( .A(n_757), .B(n_226), .Y(n_900) );
INVx3_ASAP7_75t_L g901 ( .A(n_813), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_801), .Y(n_902) );
NOR2xp33_ASAP7_75t_L g903 ( .A(n_803), .B(n_228), .Y(n_903) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_789), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_825), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_755), .B(n_229), .Y(n_906) );
BUFx3_ASAP7_75t_L g907 ( .A(n_750), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_826), .Y(n_908) );
INVx1_ASAP7_75t_SL g909 ( .A(n_734), .Y(n_909) );
OR2x2_ASAP7_75t_L g910 ( .A(n_846), .B(n_744), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_831), .B(n_801), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_846), .B(n_789), .Y(n_912) );
OAI21xp5_ASAP7_75t_SL g913 ( .A1(n_892), .A2(n_802), .B(n_737), .Y(n_913) );
AND2x2_ASAP7_75t_L g914 ( .A(n_856), .B(n_765), .Y(n_914) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_845), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_884), .B(n_766), .Y(n_916) );
OAI221xp5_ASAP7_75t_SL g917 ( .A1(n_884), .A2(n_738), .B1(n_771), .B2(n_785), .C(n_748), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_840), .B(n_789), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_861), .B(n_787), .Y(n_919) );
OR2x2_ASAP7_75t_L g920 ( .A(n_848), .B(n_779), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_854), .B(n_800), .Y(n_921) );
BUFx3_ASAP7_75t_L g922 ( .A(n_855), .Y(n_922) );
AND2x4_ASAP7_75t_L g923 ( .A(n_887), .B(n_798), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g924 ( .A(n_855), .B(n_775), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_834), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_851), .B(n_796), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_845), .B(n_735), .Y(n_927) );
NAND4xp25_ASAP7_75t_L g928 ( .A(n_903), .B(n_730), .C(n_773), .D(n_819), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_852), .B(n_796), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_857), .B(n_798), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_866), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_875), .B(n_783), .Y(n_932) );
AND2x2_ASAP7_75t_L g933 ( .A(n_887), .B(n_774), .Y(n_933) );
OAI21xp33_ASAP7_75t_L g934 ( .A1(n_889), .A2(n_786), .B(n_824), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_838), .B(n_729), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_862), .Y(n_936) );
NAND3xp33_ASAP7_75t_L g937 ( .A(n_869), .B(n_772), .C(n_818), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_864), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_880), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_899), .B(n_808), .Y(n_940) );
HB1xp67_ASAP7_75t_SL g941 ( .A(n_907), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_902), .B(n_806), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_898), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_868), .Y(n_944) );
HB1xp67_ASAP7_75t_L g945 ( .A(n_839), .Y(n_945) );
NOR2x1_ASAP7_75t_SL g946 ( .A(n_896), .B(n_817), .Y(n_946) );
INVx2_ASAP7_75t_L g947 ( .A(n_839), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_881), .Y(n_948) );
OR2x2_ASAP7_75t_L g949 ( .A(n_883), .B(n_822), .Y(n_949) );
INVx2_ASAP7_75t_L g950 ( .A(n_888), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_868), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_904), .B(n_790), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_853), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_853), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_904), .B(n_816), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_870), .B(n_736), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_858), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_871), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_943), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_911), .B(n_867), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_915), .B(n_867), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_957), .B(n_876), .Y(n_962) );
AND2x4_ASAP7_75t_SL g963 ( .A(n_923), .B(n_858), .Y(n_963) );
NOR2xp33_ASAP7_75t_L g964 ( .A(n_910), .B(n_889), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_931), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_925), .B(n_879), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_936), .Y(n_967) );
NAND2x1p5_ASAP7_75t_L g968 ( .A(n_923), .B(n_897), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_939), .B(n_890), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_930), .B(n_895), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_938), .B(n_905), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_948), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_945), .Y(n_973) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_950), .Y(n_974) );
AND2x4_ASAP7_75t_L g975 ( .A(n_958), .B(n_896), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_952), .B(n_908), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_914), .B(n_907), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_918), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_952), .B(n_909), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_918), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_916), .B(n_909), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_944), .B(n_903), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_951), .Y(n_983) );
AND2x4_ASAP7_75t_L g984 ( .A(n_947), .B(n_901), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_926), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_926), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_932), .B(n_830), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_953), .B(n_901), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_927), .B(n_900), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_976), .B(n_954), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_968), .A2(n_941), .B1(n_913), .B2(n_917), .Y(n_991) );
OAI22xp33_ASAP7_75t_SL g992 ( .A1(n_968), .A2(n_922), .B1(n_874), .B2(n_942), .Y(n_992) );
NOR2xp33_ASAP7_75t_L g993 ( .A(n_977), .B(n_924), .Y(n_993) );
NAND2x2_ASAP7_75t_L g994 ( .A(n_982), .B(n_835), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_976), .B(n_912), .Y(n_995) );
XNOR2xp5_ASAP7_75t_L g996 ( .A(n_970), .B(n_928), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_981), .B(n_933), .Y(n_997) );
INVx2_ASAP7_75t_L g998 ( .A(n_974), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_964), .A2(n_934), .B1(n_919), .B2(n_942), .Y(n_999) );
NOR2xp67_ASAP7_75t_SL g1000 ( .A(n_989), .B(n_886), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_965), .Y(n_1001) );
OAI322xp33_ASAP7_75t_L g1002 ( .A1(n_964), .A2(n_919), .A3(n_921), .B1(n_912), .B2(n_920), .C1(n_956), .C2(n_893), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_965), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_978), .B(n_921), .Y(n_1004) );
AOI22xp5_ASAP7_75t_L g1005 ( .A1(n_988), .A2(n_897), .B1(n_843), .B2(n_956), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_963), .A2(n_894), .B1(n_833), .B2(n_937), .Y(n_1006) );
OAI322xp33_ASAP7_75t_L g1007 ( .A1(n_966), .A2(n_893), .A3(n_843), .B1(n_955), .B2(n_882), .C1(n_836), .C2(n_949), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_980), .B(n_955), .Y(n_1008) );
OR2x2_ASAP7_75t_L g1009 ( .A(n_972), .B(n_929), .Y(n_1009) );
OR2x2_ASAP7_75t_L g1010 ( .A(n_995), .B(n_986), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1004), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_991), .A2(n_963), .B1(n_975), .B2(n_979), .Y(n_1012) );
A2O1A1Ixp33_ASAP7_75t_L g1013 ( .A1(n_993), .A2(n_975), .B(n_833), .C(n_900), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g1014 ( .A1(n_1006), .A2(n_979), .B1(n_987), .B2(n_960), .Y(n_1014) );
AOI21xp5_ASAP7_75t_L g1015 ( .A1(n_992), .A2(n_975), .B(n_946), .Y(n_1015) );
AND3x2_ASAP7_75t_L g1016 ( .A(n_994), .B(n_872), .C(n_863), .Y(n_1016) );
OAI221xp5_ASAP7_75t_SL g1017 ( .A1(n_999), .A2(n_894), .B1(n_971), .B2(n_961), .C(n_983), .Y(n_1017) );
INVx2_ASAP7_75t_L g1018 ( .A(n_998), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_1005), .A2(n_974), .B1(n_984), .B2(n_973), .Y(n_1019) );
OAI21xp5_ASAP7_75t_L g1020 ( .A1(n_996), .A2(n_984), .B(n_969), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_1008), .B(n_985), .Y(n_1021) );
AND2x4_ASAP7_75t_L g1022 ( .A(n_997), .B(n_984), .Y(n_1022) );
O2A1O1Ixp33_ASAP7_75t_SL g1023 ( .A1(n_1013), .A2(n_1005), .B(n_990), .C(n_1009), .Y(n_1023) );
NOR4xp25_ASAP7_75t_SL g1024 ( .A(n_1017), .B(n_1002), .C(n_967), .D(n_1001), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_1011), .B(n_969), .Y(n_1025) );
INVxp67_ASAP7_75t_SL g1026 ( .A(n_1015), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_1018), .Y(n_1027) );
AOI221xp5_ASAP7_75t_L g1028 ( .A1(n_1012), .A2(n_1007), .B1(n_1003), .B2(n_1000), .C(n_985), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_1014), .B(n_962), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_1020), .B(n_959), .Y(n_1030) );
OAI21xp33_ASAP7_75t_L g1031 ( .A1(n_1019), .A2(n_959), .B(n_940), .Y(n_1031) );
BUFx2_ASAP7_75t_L g1032 ( .A(n_1026), .Y(n_1032) );
OAI21xp5_ASAP7_75t_L g1033 ( .A1(n_1028), .A2(n_1021), .B(n_1022), .Y(n_1033) );
NOR2xp33_ASAP7_75t_L g1034 ( .A(n_1023), .B(n_1016), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1025), .Y(n_1035) );
AOI221xp5_ASAP7_75t_SL g1036 ( .A1(n_1031), .A2(n_1010), .B1(n_873), .B2(n_885), .C(n_906), .Y(n_1036) );
CKINVDCx20_ASAP7_75t_R g1037 ( .A(n_1029), .Y(n_1037) );
INVx1_ASAP7_75t_SL g1038 ( .A(n_1032), .Y(n_1038) );
AOI22xp5_ASAP7_75t_L g1039 ( .A1(n_1037), .A2(n_1030), .B1(n_1027), .B2(n_1024), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_1035), .Y(n_1040) );
OAI21x1_ASAP7_75t_SL g1041 ( .A1(n_1033), .A2(n_849), .B(n_873), .Y(n_1041) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_1034), .A2(n_844), .B1(n_935), .B2(n_891), .Y(n_1042) );
A2O1A1Ixp33_ASAP7_75t_L g1043 ( .A1(n_1039), .A2(n_1036), .B(n_859), .C(n_832), .Y(n_1043) );
AOI22xp5_ASAP7_75t_L g1044 ( .A1(n_1038), .A2(n_877), .B1(n_878), .B2(n_929), .Y(n_1044) );
OA211x2_ASAP7_75t_L g1045 ( .A1(n_1041), .A2(n_847), .B(n_860), .C(n_877), .Y(n_1045) );
O2A1O1Ixp5_ASAP7_75t_L g1046 ( .A1(n_1040), .A2(n_878), .B(n_860), .C(n_847), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1046), .Y(n_1047) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_1043), .A2(n_1042), .B1(n_842), .B2(n_841), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1044), .Y(n_1049) );
NAND2x1p5_ASAP7_75t_L g1050 ( .A(n_1047), .B(n_1045), .Y(n_1050) );
AOI221xp5_ASAP7_75t_L g1051 ( .A1(n_1049), .A2(n_865), .B1(n_837), .B2(n_850), .C(n_235), .Y(n_1051) );
OAI311xp33_ASAP7_75t_L g1052 ( .A1(n_1048), .A2(n_231), .A3(n_233), .B1(n_234), .C1(n_238), .Y(n_1052) );
CKINVDCx5p33_ASAP7_75t_R g1053 ( .A(n_1050), .Y(n_1053) );
XOR2xp5_ASAP7_75t_L g1054 ( .A(n_1052), .B(n_239), .Y(n_1054) );
NOR2x1_ASAP7_75t_L g1055 ( .A(n_1051), .B(n_240), .Y(n_1055) );
AO22x2_ASAP7_75t_L g1056 ( .A1(n_1054), .A2(n_308), .B1(n_244), .B2(n_245), .Y(n_1056) );
NOR2xp33_ASAP7_75t_L g1057 ( .A(n_1053), .B(n_241), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g1058 ( .A1(n_1055), .A2(n_246), .B1(n_248), .B2(n_249), .Y(n_1058) );
AOI31xp33_ASAP7_75t_L g1059 ( .A1(n_1057), .A2(n_250), .A3(n_251), .B(n_253), .Y(n_1059) );
BUFx2_ASAP7_75t_L g1060 ( .A(n_1056), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1058), .Y(n_1061) );
AND2x4_ASAP7_75t_L g1062 ( .A(n_1061), .B(n_254), .Y(n_1062) );
XOR2x1_ASAP7_75t_L g1063 ( .A(n_1060), .B(n_255), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_1059), .A2(n_256), .B1(n_257), .B2(n_258), .Y(n_1064) );
OAI22xp5_ASAP7_75t_SL g1065 ( .A1(n_1062), .A2(n_259), .B1(n_261), .B2(n_262), .Y(n_1065) );
OAI221xp5_ASAP7_75t_L g1066 ( .A1(n_1064), .A2(n_263), .B1(n_264), .B2(n_265), .C(n_266), .Y(n_1066) );
BUFx4f_ASAP7_75t_SL g1067 ( .A(n_1063), .Y(n_1067) );
AOI21xp5_ASAP7_75t_L g1068 ( .A1(n_1065), .A2(n_1066), .B(n_1067), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_1067), .B(n_267), .Y(n_1069) );
AOI21xp5_ASAP7_75t_L g1070 ( .A1(n_1065), .A2(n_268), .B(n_269), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_1069), .A2(n_271), .B1(n_272), .B2(n_273), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_1068), .A2(n_275), .B1(n_276), .B2(n_278), .Y(n_1072) );
OR2x6_ASAP7_75t_L g1073 ( .A(n_1072), .B(n_1070), .Y(n_1073) );
OR2x6_ASAP7_75t_L g1074 ( .A(n_1071), .B(n_279), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_1073), .A2(n_1074), .B1(n_280), .B2(n_283), .Y(n_1075) );
endmodule