module real_aes_6914_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_0), .B(n_107), .C(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g446 ( .A(n_0), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_1), .A2(n_134), .B(n_138), .C(n_233), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_2), .A2(n_170), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g467 ( .A(n_3), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_4), .A2(n_454), .B1(n_734), .B2(n_737), .C1(n_740), .C2(n_741), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_5), .B(n_210), .Y(n_267) );
AOI21xp33_ASAP7_75t_L g494 ( .A1(n_6), .A2(n_170), .B(n_495), .Y(n_494) );
AND2x6_ASAP7_75t_L g134 ( .A(n_7), .B(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g193 ( .A(n_8), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_9), .B(n_40), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_9), .B(n_40), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_10), .A2(n_169), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_11), .B(n_146), .Y(n_237) );
INVx1_ASAP7_75t_L g499 ( .A(n_12), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_13), .B(n_204), .Y(n_522) );
INVx1_ASAP7_75t_L g154 ( .A(n_14), .Y(n_154) );
INVx1_ASAP7_75t_L g544 ( .A(n_15), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_16), .A2(n_144), .B(n_218), .C(n_220), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_17), .B(n_210), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_18), .B(n_478), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_19), .B(n_170), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_20), .B(n_183), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_21), .A2(n_204), .B(n_205), .C(n_207), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_22), .B(n_210), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_23), .B(n_146), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_24), .A2(n_178), .B(n_220), .C(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_25), .B(n_146), .Y(n_145) );
CKINVDCx16_ASAP7_75t_R g250 ( .A(n_26), .Y(n_250) );
INVx1_ASAP7_75t_L g142 ( .A(n_27), .Y(n_142) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_28), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_29), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_30), .B(n_146), .Y(n_468) );
INVx1_ASAP7_75t_L g176 ( .A(n_31), .Y(n_176) );
INVx1_ASAP7_75t_L g489 ( .A(n_32), .Y(n_489) );
INVx2_ASAP7_75t_L g132 ( .A(n_33), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_34), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_35), .A2(n_204), .B(n_263), .C(n_265), .Y(n_262) );
INVxp67_ASAP7_75t_L g177 ( .A(n_36), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g137 ( .A1(n_37), .A2(n_138), .B(n_141), .C(n_149), .Y(n_137) );
CKINVDCx14_ASAP7_75t_R g261 ( .A(n_38), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_39), .A2(n_134), .B(n_138), .C(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g488 ( .A(n_41), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_42), .A2(n_191), .B(n_192), .C(n_194), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_43), .B(n_146), .Y(n_534) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_44), .A2(n_47), .B1(n_120), .B2(n_121), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_44), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_45), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_46), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_47), .Y(n_120) );
INVx1_ASAP7_75t_L g202 ( .A(n_48), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_49), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_50), .B(n_170), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_51), .A2(n_138), .B1(n_207), .B2(n_487), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_52), .Y(n_516) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_53), .Y(n_464) );
CKINVDCx14_ASAP7_75t_R g189 ( .A(n_54), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_55), .A2(n_191), .B(n_265), .C(n_498), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_56), .Y(n_537) );
INVx1_ASAP7_75t_L g496 ( .A(n_57), .Y(n_496) );
INVx1_ASAP7_75t_L g135 ( .A(n_58), .Y(n_135) );
INVx1_ASAP7_75t_L g153 ( .A(n_59), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_60), .A2(n_89), .B1(n_735), .B2(n_736), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_60), .Y(n_735) );
INVx1_ASAP7_75t_SL g264 ( .A(n_61), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_62), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_63), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_64), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g253 ( .A(n_65), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_SL g477 ( .A1(n_66), .A2(n_265), .B(n_478), .C(n_479), .Y(n_477) );
INVxp67_ASAP7_75t_L g480 ( .A(n_67), .Y(n_480) );
INVx1_ASAP7_75t_L g110 ( .A(n_68), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_69), .A2(n_170), .B(n_188), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_70), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_71), .A2(n_170), .B(n_215), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_72), .Y(n_492) );
INVx1_ASAP7_75t_L g531 ( .A(n_73), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_74), .A2(n_169), .B(n_171), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g136 ( .A(n_75), .Y(n_136) );
INVx1_ASAP7_75t_L g216 ( .A(n_76), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_77), .A2(n_134), .B(n_138), .C(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_78), .A2(n_170), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g219 ( .A(n_79), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_80), .B(n_143), .Y(n_513) );
INVx2_ASAP7_75t_L g151 ( .A(n_81), .Y(n_151) );
INVx1_ASAP7_75t_L g234 ( .A(n_82), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_83), .B(n_478), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_84), .A2(n_134), .B(n_138), .C(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g107 ( .A(n_85), .Y(n_107) );
OR2x2_ASAP7_75t_L g443 ( .A(n_85), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g733 ( .A(n_85), .B(n_445), .Y(n_733) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_86), .A2(n_138), .B(n_252), .C(n_255), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_87), .B(n_150), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_88), .Y(n_471) );
CKINVDCx14_ASAP7_75t_R g736 ( .A(n_89), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_90), .A2(n_134), .B(n_138), .C(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_91), .Y(n_526) );
INVx1_ASAP7_75t_L g476 ( .A(n_92), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_93), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_94), .B(n_143), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_95), .B(n_158), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_96), .B(n_158), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_97), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g206 ( .A(n_98), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_99), .A2(n_170), .B(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_100), .A2(n_102), .B1(n_111), .B2(n_744), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g745 ( .A(n_103), .Y(n_745) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
OR2x2_ASAP7_75t_L g731 ( .A(n_107), .B(n_445), .Y(n_731) );
NOR2x2_ASAP7_75t_L g741 ( .A(n_107), .B(n_444), .Y(n_741) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_117), .B(n_452), .Y(n_111) );
BUFx2_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g743 ( .A(n_115), .Y(n_743) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI21xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_440), .B(n_448), .Y(n_117) );
XNOR2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_122), .Y(n_118) );
INVx1_ASAP7_75t_SL g732 ( .A(n_122), .Y(n_732) );
OAI22xp5_ASAP7_75t_SL g737 ( .A1(n_122), .A2(n_456), .B1(n_729), .B2(n_738), .Y(n_737) );
OR5x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_334), .C(n_398), .D(n_414), .E(n_429), .Y(n_122) );
NAND4xp25_ASAP7_75t_L g123 ( .A(n_124), .B(n_268), .C(n_295), .D(n_318), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_211), .B(n_222), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_160), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx3_ASAP7_75t_SL g245 ( .A(n_127), .Y(n_245) );
AND2x4_ASAP7_75t_L g281 ( .A(n_127), .B(n_270), .Y(n_281) );
OR2x2_ASAP7_75t_L g291 ( .A(n_127), .B(n_247), .Y(n_291) );
OR2x2_ASAP7_75t_L g337 ( .A(n_127), .B(n_163), .Y(n_337) );
AND2x2_ASAP7_75t_L g351 ( .A(n_127), .B(n_246), .Y(n_351) );
AND2x2_ASAP7_75t_L g394 ( .A(n_127), .B(n_284), .Y(n_394) );
AND2x2_ASAP7_75t_L g401 ( .A(n_127), .B(n_258), .Y(n_401) );
AND2x2_ASAP7_75t_L g420 ( .A(n_127), .B(n_310), .Y(n_420) );
AND2x2_ASAP7_75t_L g438 ( .A(n_127), .B(n_280), .Y(n_438) );
OR2x6_ASAP7_75t_L g127 ( .A(n_128), .B(n_155), .Y(n_127) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_136), .B(n_137), .C(n_150), .Y(n_128) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_129), .A2(n_231), .B(n_232), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_129), .A2(n_250), .B(n_251), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_129), .A2(n_464), .B(n_465), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g485 ( .A1(n_129), .A2(n_180), .B1(n_486), .B2(n_490), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_129), .A2(n_531), .B(n_532), .Y(n_530) );
NAND2x1p5_ASAP7_75t_L g129 ( .A(n_130), .B(n_134), .Y(n_129) );
AND2x4_ASAP7_75t_L g170 ( .A(n_130), .B(n_134), .Y(n_170) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx1_ASAP7_75t_L g148 ( .A(n_131), .Y(n_148) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g139 ( .A(n_132), .Y(n_139) );
INVx1_ASAP7_75t_L g208 ( .A(n_132), .Y(n_208) );
INVx1_ASAP7_75t_L g140 ( .A(n_133), .Y(n_140) );
INVx3_ASAP7_75t_L g144 ( .A(n_133), .Y(n_144) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_133), .Y(n_146) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_133), .Y(n_179) );
INVx1_ASAP7_75t_L g478 ( .A(n_133), .Y(n_478) );
BUFx3_ASAP7_75t_L g149 ( .A(n_134), .Y(n_149) );
INVx4_ASAP7_75t_SL g180 ( .A(n_134), .Y(n_180) );
INVx5_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
AND2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
BUFx3_ASAP7_75t_L g195 ( .A(n_139), .Y(n_195) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_139), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_145), .C(n_147), .Y(n_141) );
OAI22xp33_ASAP7_75t_L g175 ( .A1(n_143), .A2(n_176), .B1(n_177), .B2(n_178), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_143), .A2(n_467), .B(n_468), .C(n_469), .Y(n_466) );
INVx5_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_144), .B(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_144), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_144), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
INVx4_ASAP7_75t_L g204 ( .A(n_146), .Y(n_204) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_148), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g184 ( .A(n_150), .Y(n_184) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_150), .A2(n_187), .B(n_196), .Y(n_186) );
INVx1_ASAP7_75t_L g229 ( .A(n_150), .Y(n_229) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_150), .A2(n_539), .B(n_545), .Y(n_538) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AND2x2_ASAP7_75t_L g159 ( .A(n_151), .B(n_152), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx3_ASAP7_75t_L g210 ( .A(n_157), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_157), .B(n_240), .Y(n_239) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_157), .A2(n_249), .B(n_256), .Y(n_248) );
NOR2xp33_ASAP7_75t_SL g515 ( .A(n_157), .B(n_516), .Y(n_515) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_158), .Y(n_199) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_158), .A2(n_474), .B(n_481), .Y(n_473) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g166 ( .A(n_159), .Y(n_166) );
INVx1_ASAP7_75t_L g403 ( .A(n_160), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_185), .Y(n_160) );
AND2x2_ASAP7_75t_L g313 ( .A(n_161), .B(n_246), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_161), .B(n_333), .Y(n_332) );
AOI32xp33_ASAP7_75t_L g346 ( .A1(n_161), .A2(n_347), .A3(n_350), .B1(n_352), .B2(n_356), .Y(n_346) );
AND2x2_ASAP7_75t_L g416 ( .A(n_161), .B(n_310), .Y(n_416) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g280 ( .A(n_163), .B(n_247), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_163), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g322 ( .A(n_163), .B(n_269), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_163), .B(n_401), .Y(n_400) );
AO21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_167), .B(n_181), .Y(n_163) );
INVx1_ASAP7_75t_L g285 ( .A(n_164), .Y(n_285) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_164), .A2(n_530), .B(n_536), .Y(n_529) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_SL g509 ( .A1(n_165), .A2(n_510), .B(n_511), .Y(n_509) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_166), .A2(n_463), .B(n_470), .Y(n_462) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_166), .A2(n_485), .B(n_491), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_166), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_168), .A2(n_182), .B(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_SL g171 ( .A1(n_172), .A2(n_173), .B(n_174), .C(n_180), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g188 ( .A1(n_173), .A2(n_180), .B(n_189), .C(n_190), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_SL g201 ( .A1(n_173), .A2(n_180), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_SL g215 ( .A1(n_173), .A2(n_180), .B(n_216), .C(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g260 ( .A1(n_173), .A2(n_180), .B(n_261), .C(n_262), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_173), .A2(n_180), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_173), .A2(n_180), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_173), .A2(n_180), .B(n_541), .C(n_542), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_178), .B(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_178), .B(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_178), .B(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g236 ( .A(n_179), .Y(n_236) );
OAI22xp5_ASAP7_75t_SL g487 ( .A1(n_179), .A2(n_236), .B1(n_488), .B2(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g255 ( .A(n_180), .Y(n_255) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_184), .B(n_257), .Y(n_256) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_184), .A2(n_518), .B(n_525), .Y(n_517) );
AND2x2_ASAP7_75t_L g287 ( .A(n_185), .B(n_226), .Y(n_287) );
AND2x2_ASAP7_75t_L g363 ( .A(n_185), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g435 ( .A(n_185), .Y(n_435) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_197), .Y(n_185) );
OR2x2_ASAP7_75t_L g225 ( .A(n_186), .B(n_198), .Y(n_225) );
AND2x2_ASAP7_75t_L g242 ( .A(n_186), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_186), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g294 ( .A(n_186), .Y(n_294) );
AND2x2_ASAP7_75t_L g321 ( .A(n_186), .B(n_198), .Y(n_321) );
BUFx3_ASAP7_75t_L g324 ( .A(n_186), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_186), .B(n_299), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_186), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g238 ( .A(n_194), .Y(n_238) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g220 ( .A(n_195), .Y(n_220) );
INVx2_ASAP7_75t_L g275 ( .A(n_197), .Y(n_275) );
AND2x2_ASAP7_75t_L g293 ( .A(n_197), .B(n_273), .Y(n_293) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g304 ( .A(n_198), .B(n_213), .Y(n_304) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_198), .Y(n_317) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_209), .Y(n_198) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_199), .A2(n_214), .B(n_221), .Y(n_213) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_199), .A2(n_259), .B(n_267), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_204), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g469 ( .A(n_207), .Y(n_469) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_210), .A2(n_494), .B(n_500), .Y(n_493) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_212), .B(n_324), .Y(n_374) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_SL g243 ( .A(n_213), .Y(n_243) );
NAND3xp33_ASAP7_75t_L g292 ( .A(n_213), .B(n_293), .C(n_294), .Y(n_292) );
OR2x2_ASAP7_75t_L g300 ( .A(n_213), .B(n_273), .Y(n_300) );
AND2x2_ASAP7_75t_L g320 ( .A(n_213), .B(n_273), .Y(n_320) );
AND2x2_ASAP7_75t_L g364 ( .A(n_213), .B(n_228), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_241), .B(n_244), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_224), .B(n_226), .Y(n_223) );
AND2x2_ASAP7_75t_L g439 ( .A(n_224), .B(n_364), .Y(n_439) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_225), .A2(n_337), .B1(n_379), .B2(n_381), .Y(n_378) );
OR2x2_ASAP7_75t_L g385 ( .A(n_225), .B(n_300), .Y(n_385) );
OR2x2_ASAP7_75t_L g409 ( .A(n_225), .B(n_410), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_225), .B(n_329), .Y(n_422) );
AND2x2_ASAP7_75t_L g315 ( .A(n_226), .B(n_316), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_226), .A2(n_388), .B(n_403), .Y(n_402) );
AOI32xp33_ASAP7_75t_L g423 ( .A1(n_226), .A2(n_313), .A3(n_424), .B1(n_426), .B2(n_427), .Y(n_423) );
OR2x2_ASAP7_75t_L g434 ( .A(n_226), .B(n_435), .Y(n_434) );
CKINVDCx16_ASAP7_75t_R g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g302 ( .A(n_227), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_227), .B(n_316), .Y(n_381) );
BUFx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx4_ASAP7_75t_L g273 ( .A(n_228), .Y(n_273) );
AND2x2_ASAP7_75t_L g339 ( .A(n_228), .B(n_304), .Y(n_339) );
AND3x2_ASAP7_75t_L g348 ( .A(n_228), .B(n_242), .C(n_349), .Y(n_348) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_239), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_229), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_229), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_229), .B(n_537), .Y(n_536) );
O2A1O1Ixp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_237), .C(n_238), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_235), .A2(n_238), .B(n_253), .C(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_238), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_238), .A2(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g274 ( .A(n_243), .B(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_243), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_243), .B(n_273), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
AND2x2_ASAP7_75t_L g269 ( .A(n_245), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g309 ( .A(n_245), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g327 ( .A(n_245), .B(n_258), .Y(n_327) );
AND2x2_ASAP7_75t_L g345 ( .A(n_245), .B(n_247), .Y(n_345) );
OR2x2_ASAP7_75t_L g359 ( .A(n_245), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g405 ( .A(n_245), .B(n_333), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_246), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_258), .Y(n_246) );
AND2x2_ASAP7_75t_L g306 ( .A(n_247), .B(n_284), .Y(n_306) );
OR2x2_ASAP7_75t_L g360 ( .A(n_247), .B(n_284), .Y(n_360) );
AND2x2_ASAP7_75t_L g413 ( .A(n_247), .B(n_270), .Y(n_413) );
INVx2_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
BUFx2_ASAP7_75t_L g311 ( .A(n_248), .Y(n_311) );
AND2x2_ASAP7_75t_L g333 ( .A(n_248), .B(n_258), .Y(n_333) );
INVx2_ASAP7_75t_L g270 ( .A(n_258), .Y(n_270) );
INVx1_ASAP7_75t_L g290 ( .A(n_258), .Y(n_290) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_266), .Y(n_523) );
AOI211xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_271), .B(n_276), .C(n_288), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_269), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g432 ( .A(n_269), .Y(n_432) );
AND2x2_ASAP7_75t_L g310 ( .A(n_270), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_273), .B(n_274), .Y(n_282) );
INVx1_ASAP7_75t_L g367 ( .A(n_273), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_273), .B(n_294), .Y(n_391) );
AND2x2_ASAP7_75t_L g407 ( .A(n_273), .B(n_321), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_274), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g298 ( .A(n_275), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_282), .B1(n_283), .B2(n_286), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_279), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_280), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g305 ( .A(n_281), .B(n_306), .Y(n_305) );
AOI221xp5_ASAP7_75t_SL g370 ( .A1(n_281), .A2(n_323), .B1(n_371), .B2(n_376), .C(n_378), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_281), .B(n_344), .Y(n_377) );
INVx1_ASAP7_75t_L g437 ( .A(n_283), .Y(n_437) );
BUFx3_ASAP7_75t_L g344 ( .A(n_284), .Y(n_344) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AOI21xp33_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_291), .B(n_292), .Y(n_288) );
INVx1_ASAP7_75t_L g353 ( .A(n_290), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_290), .B(n_344), .Y(n_397) );
INVx1_ASAP7_75t_L g354 ( .A(n_291), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_291), .B(n_344), .Y(n_355) );
INVxp67_ASAP7_75t_L g375 ( .A(n_293), .Y(n_375) );
AND2x2_ASAP7_75t_L g316 ( .A(n_294), .B(n_317), .Y(n_316) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_301), .B(n_305), .C(n_307), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_SL g330 ( .A(n_298), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_299), .B(n_330), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_299), .B(n_321), .Y(n_372) );
INVx2_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_302), .A2(n_308), .B1(n_312), .B2(n_314), .Y(n_307) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g323 ( .A(n_304), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g368 ( .A(n_304), .B(n_369), .Y(n_368) );
OAI21xp33_ASAP7_75t_L g371 ( .A1(n_306), .A2(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_310), .A2(n_319), .B1(n_322), .B2(n_323), .C(n_325), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_310), .B(n_344), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_310), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g426 ( .A(n_316), .Y(n_426) );
INVxp67_ASAP7_75t_L g349 ( .A(n_317), .Y(n_349) );
INVx1_ASAP7_75t_L g356 ( .A(n_319), .Y(n_356) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g395 ( .A(n_320), .B(n_324), .Y(n_395) );
INVx1_ASAP7_75t_L g369 ( .A(n_324), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_324), .B(n_339), .Y(n_399) );
OAI32xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .A3(n_330), .B1(n_331), .B2(n_332), .Y(n_325) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_SL g338 ( .A(n_333), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_333), .B(n_365), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_333), .B(n_394), .Y(n_425) );
NAND2x1p5_ASAP7_75t_L g433 ( .A(n_333), .B(n_344), .Y(n_433) );
NAND5xp2_ASAP7_75t_L g334 ( .A(n_335), .B(n_357), .C(n_370), .D(n_382), .E(n_383), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_339), .B1(n_340), .B2(n_342), .C(n_346), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp33_ASAP7_75t_SL g361 ( .A(n_341), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_344), .B(n_413), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_345), .A2(n_358), .B1(n_361), .B2(n_365), .Y(n_357) );
INVx2_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
OAI211xp5_ASAP7_75t_SL g352 ( .A1(n_348), .A2(n_353), .B(n_354), .C(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g380 ( .A(n_360), .Y(n_380) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_369), .B(n_418), .Y(n_428) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI222xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .B1(n_388), .B2(n_392), .C1(n_395), .C2(n_396), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_402), .B2(n_404), .C(n_406), .Y(n_398) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
OAI21xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B(n_411), .Y(n_406) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g418 ( .A(n_410), .Y(n_418) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_417), .B1(n_419), .B2(n_421), .C(n_423), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
A2O1A1Ixp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_433), .B(n_434), .C(n_436), .Y(n_429) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI21xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B(n_439), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g451 ( .A(n_443), .Y(n_451) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_448), .B(n_453), .C(n_742), .Y(n_452) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OAI22xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_729), .B1(n_732), .B2(n_733), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR4x1_ASAP7_75t_L g456 ( .A(n_457), .B(n_618), .C(n_678), .D(n_705), .Y(n_456) );
NAND4xp25_ASAP7_75t_SL g457 ( .A(n_458), .B(n_566), .C(n_597), .D(n_614), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_501), .B(n_503), .C(n_546), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_482), .Y(n_459) );
INVx1_ASAP7_75t_L g608 ( .A(n_460), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_460), .A2(n_649), .B1(n_697), .B2(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_472), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_461), .B(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g559 ( .A(n_461), .B(n_484), .Y(n_559) );
AND2x2_ASAP7_75t_L g601 ( .A(n_461), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_461), .B(n_502), .Y(n_613) );
INVx1_ASAP7_75t_L g653 ( .A(n_461), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_461), .B(n_707), .Y(n_706) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g581 ( .A(n_462), .B(n_484), .Y(n_581) );
INVx3_ASAP7_75t_L g585 ( .A(n_462), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_462), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g672 ( .A(n_472), .B(n_493), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_472), .B(n_585), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_472), .B(n_700), .Y(n_699) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g502 ( .A(n_473), .B(n_484), .Y(n_502) );
INVx1_ASAP7_75t_L g554 ( .A(n_473), .Y(n_554) );
BUFx2_ASAP7_75t_L g558 ( .A(n_473), .Y(n_558) );
AND2x2_ASAP7_75t_L g602 ( .A(n_473), .B(n_483), .Y(n_602) );
OR2x2_ASAP7_75t_L g641 ( .A(n_473), .B(n_483), .Y(n_641) );
AND2x2_ASAP7_75t_L g666 ( .A(n_473), .B(n_493), .Y(n_666) );
AND2x2_ASAP7_75t_L g725 ( .A(n_473), .B(n_555), .Y(n_725) );
INVx1_ASAP7_75t_L g700 ( .A(n_482), .Y(n_700) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_493), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_483), .B(n_493), .Y(n_586) );
AND2x2_ASAP7_75t_L g596 ( .A(n_483), .B(n_585), .Y(n_596) );
BUFx2_ASAP7_75t_L g607 ( .A(n_483), .Y(n_607) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g629 ( .A(n_484), .B(n_493), .Y(n_629) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_484), .Y(n_684) );
AND2x2_ASAP7_75t_SL g501 ( .A(n_493), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_SL g555 ( .A(n_493), .Y(n_555) );
BUFx2_ASAP7_75t_L g580 ( .A(n_493), .Y(n_580) );
INVx2_ASAP7_75t_L g599 ( .A(n_493), .Y(n_599) );
AND2x2_ASAP7_75t_L g661 ( .A(n_493), .B(n_585), .Y(n_661) );
AOI321xp33_ASAP7_75t_L g680 ( .A1(n_501), .A2(n_681), .A3(n_682), .B1(n_683), .B2(n_685), .C(n_686), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_502), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_502), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g674 ( .A(n_502), .B(n_653), .Y(n_674) );
AND2x2_ASAP7_75t_L g707 ( .A(n_502), .B(n_599), .Y(n_707) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_527), .Y(n_504) );
OR2x2_ASAP7_75t_L g609 ( .A(n_505), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_517), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g561 ( .A(n_508), .Y(n_561) );
AND2x2_ASAP7_75t_L g571 ( .A(n_508), .B(n_529), .Y(n_571) );
AND2x2_ASAP7_75t_L g576 ( .A(n_508), .B(n_551), .Y(n_576) );
INVx1_ASAP7_75t_L g593 ( .A(n_508), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_508), .B(n_574), .Y(n_612) );
AND2x2_ASAP7_75t_L g617 ( .A(n_508), .B(n_550), .Y(n_617) );
OR2x2_ASAP7_75t_L g649 ( .A(n_508), .B(n_638), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_508), .B(n_562), .Y(n_688) );
AND2x2_ASAP7_75t_L g722 ( .A(n_508), .B(n_548), .Y(n_722) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_515), .Y(n_508) );
INVx1_ASAP7_75t_L g549 ( .A(n_517), .Y(n_549) );
INVx2_ASAP7_75t_L g564 ( .A(n_517), .Y(n_564) );
AND2x2_ASAP7_75t_L g604 ( .A(n_517), .B(n_575), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_517), .B(n_551), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_524), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B(n_523), .Y(n_520) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g710 ( .A(n_528), .B(n_561), .Y(n_710) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_538), .Y(n_528) );
INVx2_ASAP7_75t_L g551 ( .A(n_529), .Y(n_551) );
AND2x2_ASAP7_75t_L g704 ( .A(n_529), .B(n_564), .Y(n_704) );
AND2x2_ASAP7_75t_L g550 ( .A(n_538), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g565 ( .A(n_538), .Y(n_565) );
INVx1_ASAP7_75t_L g575 ( .A(n_538), .Y(n_575) );
OAI22xp33_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_552), .B1(n_556), .B2(n_560), .Y(n_546) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_547), .A2(n_665), .B1(n_702), .B2(n_703), .Y(n_701) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g616 ( .A(n_549), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_550), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g611 ( .A(n_551), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_551), .B(n_564), .Y(n_638) );
INVx1_ASAP7_75t_L g654 ( .A(n_551), .Y(n_654) );
AND2x2_ASAP7_75t_L g595 ( .A(n_553), .B(n_596), .Y(n_595) );
INVx3_ASAP7_75t_SL g634 ( .A(n_553), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_553), .B(n_559), .Y(n_711) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g720 ( .A(n_556), .Y(n_720) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_557), .B(n_653), .Y(n_695) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx3_ASAP7_75t_SL g600 ( .A(n_559), .Y(n_600) );
NAND2x1_ASAP7_75t_SL g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AND2x2_ASAP7_75t_L g621 ( .A(n_561), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g628 ( .A(n_561), .B(n_565), .Y(n_628) );
AND2x2_ASAP7_75t_L g633 ( .A(n_561), .B(n_574), .Y(n_633) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_561), .Y(n_682) );
OAI311xp33_ASAP7_75t_L g705 ( .A1(n_562), .A2(n_706), .A3(n_708), .B1(n_709), .C1(n_719), .Y(n_705) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g718 ( .A(n_563), .B(n_591), .Y(n_718) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g574 ( .A(n_564), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g622 ( .A(n_564), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g677 ( .A(n_564), .Y(n_677) );
INVx1_ASAP7_75t_L g570 ( .A(n_565), .Y(n_570) );
INVx1_ASAP7_75t_L g590 ( .A(n_565), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_565), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g623 ( .A(n_565), .Y(n_623) );
AOI221xp5_ASAP7_75t_SL g566 ( .A1(n_567), .A2(n_569), .B1(n_577), .B2(n_582), .C(n_587), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx4_ASAP7_75t_L g591 ( .A(n_571), .Y(n_591) );
AND2x2_ASAP7_75t_L g685 ( .A(n_571), .B(n_604), .Y(n_685) );
AND2x2_ASAP7_75t_L g692 ( .A(n_571), .B(n_574), .Y(n_692) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_574), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g603 ( .A(n_576), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_579), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g728 ( .A(n_581), .B(n_672), .Y(n_728) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g713 ( .A(n_585), .B(n_641), .Y(n_713) );
OAI211xp5_ASAP7_75t_L g678 ( .A1(n_586), .A2(n_679), .B(n_680), .C(n_693), .Y(n_678) );
AOI21xp33_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_592), .B(n_594), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp67_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g657 ( .A(n_591), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g686 ( .A1(n_592), .A2(n_687), .B1(n_688), .B2(n_689), .C(n_690), .Y(n_686) );
AND2x2_ASAP7_75t_L g663 ( .A(n_593), .B(n_604), .Y(n_663) );
AND2x2_ASAP7_75t_L g716 ( .A(n_593), .B(n_611), .Y(n_716) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_596), .B(n_634), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_601), .B(n_603), .C(n_605), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g644 ( .A(n_599), .B(n_602), .Y(n_644) );
OR2x2_ASAP7_75t_L g687 ( .A(n_599), .B(n_641), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_600), .B(n_666), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_600), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g631 ( .A(n_601), .Y(n_631) );
INVx1_ASAP7_75t_L g697 ( .A(n_604), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_609), .B1(n_612), .B2(n_613), .Y(n_605) );
INVx1_ASAP7_75t_L g620 ( .A(n_606), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_607), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g683 ( .A(n_608), .B(n_684), .Y(n_683) );
INVxp67_ASAP7_75t_L g669 ( .A(n_610), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_611), .B(n_697), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g670 ( .A1(n_612), .A2(n_671), .B1(n_673), .B2(n_675), .Y(n_670) );
INVx1_ASAP7_75t_L g679 ( .A(n_615), .Y(n_679) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g721 ( .A(n_616), .B(n_716), .Y(n_721) );
AOI222xp33_ASAP7_75t_L g650 ( .A1(n_617), .A2(n_651), .B1(n_654), .B2(n_655), .C1(n_658), .C2(n_659), .Y(n_650) );
NAND4xp25_ASAP7_75t_SL g618 ( .A(n_619), .B(n_639), .C(n_650), .D(n_662), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_624), .B2(n_629), .C(n_630), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_622), .B(n_657), .Y(n_656) );
INVxp67_ASAP7_75t_L g648 ( .A(n_623), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_624), .A2(n_694), .B1(n_696), .B2(n_698), .C(n_701), .Y(n_693) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g636 ( .A(n_628), .B(n_637), .Y(n_636) );
OAI21xp33_ASAP7_75t_L g690 ( .A1(n_629), .A2(n_691), .B(n_692), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_634), .B2(n_635), .Y(n_630) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI21xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B(n_645), .Y(n_639) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g681 ( .A(n_652), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_653), .B(n_672), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_653), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_657), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g689 ( .A(n_661), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_667), .B2(n_669), .C(n_670), .Y(n_662) );
INVxp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI222xp33_ASAP7_75t_L g709 ( .A1(n_672), .A2(n_710), .B1(n_711), .B2(n_712), .C1(n_714), .C2(n_717), .Y(n_709) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_676), .B(n_716), .Y(n_715) );
INVxp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g708 ( .A(n_682), .Y(n_708) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVxp33_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .B1(n_722), .B2(n_723), .C(n_726), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVxp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g739 ( .A(n_733), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_734), .Y(n_740) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
endmodule