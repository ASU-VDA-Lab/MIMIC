module fake_jpeg_9337_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_19),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_0),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_20),
.Y(n_27)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_8),
.A2(n_1),
.B1(n_6),
.B2(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_9),
.C(n_12),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_29),
.C(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_9),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_18),
.C(n_22),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_29),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_18),
.B(n_17),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_13),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_24),
.C(n_31),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_41),
.C(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_45),
.B(n_40),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_47),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_49),
.A2(n_48),
.B(n_31),
.Y(n_50)
);

AOI21x1_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_23),
.B(n_29),
.Y(n_51)
);


endmodule