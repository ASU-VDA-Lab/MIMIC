module fake_jpeg_17945_n_330 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_45),
.Y(n_69)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_42),
.B(n_26),
.Y(n_110)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_17),
.B(n_13),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_46),
.B(n_49),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_17),
.B(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_50),
.B(n_52),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_29),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_18),
.B(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_21),
.B(n_11),
.Y(n_57)
);

BUFx2_ASAP7_75t_R g58 ( 
.A(n_22),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_58),
.B(n_15),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_21),
.B(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_29),
.B(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_65),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_16),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_70),
.B(n_83),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_72),
.B(n_87),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_33),
.B(n_31),
.C(n_19),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_74),
.A2(n_79),
.B(n_107),
.C(n_119),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_15),
.C(n_64),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_76),
.B(n_99),
.C(n_22),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_22),
.B(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_31),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_28),
.B1(n_36),
.B2(n_34),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_37),
.B1(n_9),
.B2(n_7),
.Y(n_123)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_89),
.B(n_90),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_40),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_48),
.A2(n_28),
.B1(n_34),
.B2(n_32),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_1),
.B(n_2),
.Y(n_121)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_51),
.A2(n_15),
.B1(n_28),
.B2(n_23),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_105),
.B1(n_3),
.B2(n_4),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_15),
.C(n_32),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g101 ( 
.A(n_63),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_101),
.Y(n_156)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_53),
.A2(n_37),
.B1(n_25),
.B2(n_23),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_45),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_113),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_7),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_66),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_68),
.Y(n_115)
);

OR2x2_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_54),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_58),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_119),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_33),
.B1(n_19),
.B2(n_7),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_121),
.A2(n_129),
.B1(n_143),
.B2(n_148),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_37),
.B1(n_23),
.B2(n_15),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_122),
.A2(n_123),
.B1(n_136),
.B2(n_147),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_153),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_125),
.B(n_130),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_71),
.A2(n_116),
.B1(n_84),
.B2(n_100),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_71),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_78),
.Y(n_130)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_4),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_139),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_138),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_6),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_93),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_150),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_84),
.B1(n_100),
.B2(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_155),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_103),
.A2(n_80),
.B1(n_97),
.B2(n_74),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_91),
.B1(n_98),
.B2(n_92),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_69),
.A2(n_72),
.B(n_87),
.C(n_89),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_145),
.B(n_163),
.C(n_154),
.D(n_132),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_81),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_88),
.A2(n_94),
.B1(n_112),
.B2(n_107),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_152),
.B(n_159),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_77),
.A2(n_85),
.B(n_75),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_154),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_75),
.A2(n_79),
.B(n_110),
.C(n_119),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_96),
.B(n_109),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_162),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_109),
.A2(n_27),
.B1(n_76),
.B2(n_110),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_95),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_160)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_137),
.A3(n_139),
.B1(n_157),
.B2(n_131),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_76),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

BUFx4f_ASAP7_75t_SL g165 ( 
.A(n_96),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_166),
.B(n_162),
.Y(n_169)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_138),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_190),
.C(n_182),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_178),
.A2(n_207),
.B1(n_197),
.B2(n_199),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_180),
.A2(n_193),
.B(n_165),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_146),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_190),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_133),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_188),
.B(n_192),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_130),
.B(n_166),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_125),
.B(n_141),
.Y(n_192)
);

AND2x4_ASAP7_75t_L g193 ( 
.A(n_121),
.B(n_145),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_125),
.B(n_144),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_194),
.B(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_156),
.B(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_199),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_124),
.B(n_135),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_200),
.B(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_135),
.Y(n_201)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_126),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_132),
.B(n_149),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_134),
.Y(n_205)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

OAI32xp33_ASAP7_75t_L g207 ( 
.A1(n_160),
.A2(n_143),
.A3(n_164),
.B1(n_142),
.B2(n_127),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_231),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_215),
.C(n_230),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_167),
.Y(n_213)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_165),
.C(n_142),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_220),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_127),
.Y(n_217)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_217),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_219),
.A2(n_236),
.B(n_205),
.Y(n_246)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_224),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_174),
.A2(n_173),
.B1(n_178),
.B2(n_183),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_222),
.A2(n_223),
.B1(n_218),
.B2(n_212),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_174),
.A2(n_183),
.B1(n_207),
.B2(n_203),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_193),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_240),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_169),
.B(n_186),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_177),
.B(n_170),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_189),
.A2(n_168),
.B1(n_195),
.B2(n_176),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_237),
.B1(n_239),
.B2(n_215),
.Y(n_260)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_172),
.A2(n_180),
.B(n_195),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_168),
.A2(n_176),
.B1(n_172),
.B2(n_187),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_175),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_210),
.B(n_231),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_197),
.C(n_204),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_244),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_242),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_226),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_257),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_246),
.B(n_261),
.Y(n_279)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_196),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_256),
.B(n_265),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_223),
.A2(n_171),
.B1(n_184),
.B2(n_239),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_251),
.Y(n_281)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_219),
.A2(n_236),
.B(n_229),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_184),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_209),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_259),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_263),
.B1(n_265),
.B2(n_258),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_SL g264 ( 
.A1(n_218),
.A2(n_208),
.B(n_235),
.C(n_214),
.Y(n_264)
);

AO21x1_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_208),
.B(n_225),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_227),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_238),
.Y(n_270)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_267),
.A2(n_270),
.B(n_274),
.Y(n_297)
);

OA21x2_ASAP7_75t_SL g272 ( 
.A1(n_246),
.A2(n_228),
.B(n_224),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_264),
.Y(n_292)
);

OA21x2_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_225),
.B(n_221),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_211),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_254),
.C(n_252),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_247),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_285),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_266),
.A2(n_256),
.B1(n_244),
.B2(n_263),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_280),
.B1(n_258),
.B2(n_261),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_249),
.A2(n_262),
.B1(n_241),
.B2(n_265),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_278),
.A2(n_274),
.B1(n_272),
.B2(n_286),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_264),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_248),
.Y(n_295)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_247),
.Y(n_286)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_282),
.Y(n_287)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_243),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_290),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_268),
.B1(n_277),
.B2(n_267),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_292),
.A2(n_293),
.B1(n_296),
.B2(n_298),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_264),
.B(n_254),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_267),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_242),
.B1(n_255),
.B2(n_270),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_284),
.B(n_280),
.Y(n_298)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_271),
.Y(n_302)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_308),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_291),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_307),
.B(n_282),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_295),
.B1(n_297),
.B2(n_292),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_312),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_288),
.C(n_290),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_306),
.B(n_283),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_303),
.A3(n_309),
.B1(n_308),
.B2(n_310),
.C1(n_304),
.C2(n_301),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_322),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_317),
.A2(n_298),
.B1(n_297),
.B2(n_311),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_319),
.B(n_315),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_323),
.B(n_325),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_283),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_313),
.C(n_305),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_323),
.B(n_321),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_328),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_327),
.Y(n_330)
);


endmodule