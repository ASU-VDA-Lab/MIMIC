module fake_aes_12693_n_703 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_703);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_703;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_490;
wire n_247;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g87 ( .A(n_66), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_48), .Y(n_88) );
INVx2_ASAP7_75t_SL g89 ( .A(n_78), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_60), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_29), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_80), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_75), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_25), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_27), .Y(n_95) );
BUFx6f_ASAP7_75t_L g96 ( .A(n_17), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_19), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_32), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_21), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_28), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_71), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_67), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_63), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_4), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_12), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_38), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_10), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_43), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_15), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_35), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_77), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_47), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_6), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_55), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_3), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_76), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_70), .Y(n_117) );
INVxp67_ASAP7_75t_L g118 ( .A(n_15), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_18), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_51), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_42), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_5), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_46), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_23), .Y(n_124) );
OR2x2_ASAP7_75t_L g125 ( .A(n_26), .B(n_0), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_79), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_110), .Y(n_127) );
AOI22xp5_ASAP7_75t_SL g128 ( .A1(n_105), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_128) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_123), .B(n_86), .Y(n_129) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_110), .A2(n_53), .B(n_84), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_89), .B(n_1), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_102), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_112), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_112), .Y(n_134) );
BUFx12f_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
INVx5_ASAP7_75t_L g138 ( .A(n_96), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_107), .B(n_2), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_105), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_140) );
INVx2_ASAP7_75t_SL g141 ( .A(n_88), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_90), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_96), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_92), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_104), .B(n_6), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_96), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_139), .B(n_107), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_141), .B(n_122), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_132), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_141), .B(n_122), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_133), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_136), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_133), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_133), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_142), .B(n_100), .Y(n_155) );
INVx4_ASAP7_75t_L g156 ( .A(n_130), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_129), .B(n_91), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_133), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_133), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_142), .B(n_93), .Y(n_160) );
OR2x6_ASAP7_75t_L g161 ( .A(n_140), .B(n_125), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_136), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_137), .B(n_94), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_129), .B(n_94), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_133), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
NAND2x1p5_ASAP7_75t_L g168 ( .A(n_129), .B(n_97), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_143), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_127), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_135), .B(n_95), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_139), .A2(n_115), .B1(n_118), .B2(n_113), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_143), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_137), .B(n_95), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_127), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_164), .B(n_135), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_160), .A2(n_144), .B(n_137), .C(n_127), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_148), .B(n_135), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_170), .Y(n_181) );
NAND2xp33_ASAP7_75t_SL g182 ( .A(n_157), .B(n_120), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_150), .B(n_131), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_170), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_147), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_177), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_168), .A2(n_131), .B1(n_144), .B2(n_145), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_168), .A2(n_120), .B1(n_128), .B2(n_145), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_165), .A2(n_109), .B1(n_140), .B2(n_144), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_176), .B(n_119), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_147), .B(n_119), .Y(n_192) );
INVx4_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_155), .B(n_126), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_152), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_168), .B(n_126), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_174), .B(n_98), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_152), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_161), .A2(n_134), .B1(n_113), .B2(n_96), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_177), .Y(n_200) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_156), .A2(n_130), .B(n_106), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_149), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_152), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_171), .B(n_99), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_162), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_162), .B(n_101), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_161), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_163), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_163), .B(n_103), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_161), .A2(n_134), .B(n_117), .C(n_116), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_163), .B(n_134), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_163), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_156), .B(n_108), .Y(n_215) );
INVx2_ASAP7_75t_SL g216 ( .A(n_156), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_161), .B(n_111), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_185), .B(n_161), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g219 ( .A1(n_189), .A2(n_128), .B1(n_130), .B2(n_113), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_200), .Y(n_220) );
NAND3xp33_ASAP7_75t_L g221 ( .A(n_199), .B(n_130), .C(n_114), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_185), .A2(n_121), .B(n_124), .C(n_146), .Y(n_222) );
O2A1O1Ixp5_ASAP7_75t_L g223 ( .A1(n_201), .A2(n_154), .B(n_151), .C(n_153), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_SL g224 ( .A1(n_179), .A2(n_159), .B(n_151), .C(n_153), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_200), .B(n_113), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_183), .B(n_130), .Y(n_226) );
NAND3xp33_ASAP7_75t_L g227 ( .A(n_212), .B(n_159), .C(n_158), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_209), .B(n_181), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_181), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_217), .B(n_146), .Y(n_230) );
AOI21x1_ASAP7_75t_L g231 ( .A1(n_204), .A2(n_166), .B(n_158), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_202), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_216), .A2(n_215), .B(n_187), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_182), .A2(n_146), .B1(n_166), .B2(n_138), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_216), .A2(n_154), .B(n_172), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_192), .B(n_7), .Y(n_236) );
NOR2xp33_ASAP7_75t_SL g237 ( .A(n_202), .B(n_154), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_187), .A2(n_172), .B(n_173), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_184), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_180), .B(n_7), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_187), .A2(n_175), .B(n_173), .Y(n_241) );
AO22x1_ASAP7_75t_L g242 ( .A1(n_196), .A2(n_138), .B1(n_143), .B2(n_146), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_178), .B(n_8), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_188), .B(n_138), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_184), .A2(n_175), .B(n_173), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_187), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_186), .Y(n_247) );
NOR2xp67_ASAP7_75t_L g248 ( .A(n_193), .B(n_186), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_191), .B(n_138), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_187), .A2(n_204), .B(n_195), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_220), .Y(n_251) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_223), .A2(n_213), .B(n_198), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_226), .A2(n_208), .B(n_206), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_218), .B(n_190), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_231), .A2(n_198), .B(n_207), .Y(n_255) );
INVxp67_ASAP7_75t_SL g256 ( .A(n_220), .Y(n_256) );
INVx5_ASAP7_75t_L g257 ( .A(n_246), .Y(n_257) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_231), .A2(n_210), .B(n_207), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_233), .A2(n_214), .B(n_203), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_228), .A2(n_182), .B1(n_194), .B2(n_197), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_228), .B(n_193), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_229), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_229), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_239), .A2(n_210), .B(n_205), .C(n_211), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_235), .A2(n_193), .B(n_175), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_239), .B(n_8), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_250), .A2(n_169), .B(n_167), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_247), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_246), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_232), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_221), .A2(n_169), .B(n_167), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_247), .A2(n_169), .B(n_167), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_219), .B(n_9), .Y(n_273) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_271), .A2(n_245), .B(n_241), .Y(n_274) );
AOI21xp33_ASAP7_75t_SL g275 ( .A1(n_273), .A2(n_236), .B(n_240), .Y(n_275) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_271), .A2(n_238), .B(n_244), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_254), .B(n_243), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_262), .B(n_248), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_257), .B(n_237), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_263), .B(n_234), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_255), .A2(n_225), .B(n_249), .Y(n_281) );
OAI21x1_ASAP7_75t_SL g282 ( .A1(n_266), .A2(n_222), .B(n_230), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_253), .A2(n_224), .B(n_248), .Y(n_283) );
AO31x2_ASAP7_75t_L g284 ( .A1(n_264), .A2(n_227), .A3(n_242), .B(n_138), .Y(n_284) );
AO21x2_ASAP7_75t_L g285 ( .A1(n_255), .A2(n_227), .B(n_242), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_258), .A2(n_58), .B(n_85), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_268), .B(n_9), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_251), .Y(n_288) );
NOR2xp67_ASAP7_75t_SL g289 ( .A(n_257), .B(n_138), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_251), .Y(n_290) );
OAI21x1_ASAP7_75t_SL g291 ( .A1(n_259), .A2(n_10), .B(n_11), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_260), .B(n_11), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_270), .B(n_12), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_258), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_251), .Y(n_295) );
AO21x2_ASAP7_75t_L g296 ( .A1(n_291), .A2(n_264), .B(n_252), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_288), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_278), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_294), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_294), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_288), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_287), .B(n_261), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_294), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_278), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_287), .B(n_256), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_290), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_284), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_290), .Y(n_308) );
OAI21x1_ASAP7_75t_L g309 ( .A1(n_276), .A2(n_252), .B(n_265), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_295), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_295), .B(n_257), .Y(n_311) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_279), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_291), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_276), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_284), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_286), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_285), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_284), .B(n_257), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_286), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
OR2x6_ASAP7_75t_L g321 ( .A(n_282), .B(n_269), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_293), .B(n_257), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_284), .B(n_269), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_284), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_284), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_282), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_292), .B(n_269), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_310), .B(n_285), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_297), .B(n_277), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_297), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_310), .B(n_280), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_301), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_318), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_310), .B(n_269), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_301), .B(n_13), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_306), .B(n_13), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_306), .B(n_14), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_304), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_318), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_318), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_299), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_308), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_318), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_308), .B(n_14), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_299), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_304), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_305), .A2(n_275), .B1(n_283), .B2(n_289), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_304), .B(n_275), .Y(n_348) );
AND2x4_ASAP7_75t_SL g349 ( .A(n_311), .B(n_289), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_298), .B(n_16), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_321), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_299), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_324), .B(n_274), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_324), .B(n_274), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_298), .B(n_16), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_325), .B(n_323), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_300), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_325), .B(n_281), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_323), .B(n_281), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_323), .B(n_17), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_300), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_300), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_298), .B(n_20), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_298), .B(n_22), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_303), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_303), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_326), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_303), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_317), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_313), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_313), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_307), .B(n_24), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_326), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_326), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_305), .B(n_307), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_315), .B(n_138), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_321), .Y(n_377) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_314), .Y(n_378) );
AND2x2_ASAP7_75t_SL g379 ( .A(n_315), .B(n_30), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_321), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_311), .B(n_272), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_321), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_360), .B(n_302), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_360), .B(n_302), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_356), .B(n_317), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_356), .B(n_317), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_330), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_375), .B(n_320), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_356), .B(n_320), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_346), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_341), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_338), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_341), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_339), .B(n_321), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_360), .B(n_322), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_329), .B(n_327), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_330), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_338), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_359), .B(n_320), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_341), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_369), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_332), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_329), .B(n_327), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_369), .Y(n_404) );
INVx4_ASAP7_75t_L g405 ( .A(n_379), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_359), .B(n_296), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_369), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_359), .B(n_296), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_362), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_332), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_333), .B(n_296), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_333), .B(n_296), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_342), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_362), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_342), .Y(n_415) );
AOI21xp33_ASAP7_75t_L g416 ( .A1(n_348), .A2(n_312), .B(n_321), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_343), .B(n_319), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_343), .B(n_319), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_340), .B(n_316), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_370), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_375), .B(n_312), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_340), .B(n_316), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_340), .B(n_314), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_339), .B(n_314), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_353), .B(n_314), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_353), .B(n_314), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_370), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_376), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_335), .B(n_314), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_371), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_335), .B(n_309), .Y(n_431) );
AND2x4_ASAP7_75t_SL g432 ( .A(n_339), .B(n_309), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_353), .B(n_309), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_367), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_371), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_339), .B(n_267), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_354), .B(n_31), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_378), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_382), .B(n_33), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_374), .B(n_34), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_345), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_336), .B(n_36), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_345), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_352), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_354), .B(n_37), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_374), .B(n_39), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_362), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_365), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_365), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_365), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_367), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_366), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_378), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_366), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_354), .B(n_40), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_352), .Y(n_456) );
NOR2xp67_ASAP7_75t_L g457 ( .A(n_350), .B(n_41), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_357), .B(n_361), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_328), .B(n_44), .Y(n_459) );
BUFx2_ASAP7_75t_SL g460 ( .A(n_367), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_328), .B(n_358), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_366), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_358), .B(n_45), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_387), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_428), .B(n_357), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_395), .B(n_348), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_461), .B(n_331), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_461), .B(n_361), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_385), .B(n_331), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_387), .B(n_358), .Y(n_470) );
INVx3_ASAP7_75t_L g471 ( .A(n_434), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_385), .B(n_373), .Y(n_472) );
INVxp67_ASAP7_75t_L g473 ( .A(n_460), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_397), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_440), .B(n_379), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_386), .B(n_373), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_458), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_397), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_434), .B(n_382), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_402), .B(n_368), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_386), .B(n_389), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_389), .B(n_380), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_401), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_410), .B(n_368), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_413), .B(n_368), .Y(n_485) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_405), .A2(n_379), .B1(n_336), .B2(n_337), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_434), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_415), .B(n_376), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_396), .B(n_355), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_399), .B(n_380), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_420), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_390), .B(n_337), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_399), .B(n_351), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_420), .B(n_376), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_392), .B(n_351), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_401), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_398), .B(n_377), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_458), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_451), .B(n_382), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_451), .B(n_382), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_427), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_403), .B(n_355), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_451), .B(n_377), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_427), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_430), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_406), .B(n_372), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_430), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_435), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_435), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_406), .B(n_372), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_441), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_409), .Y(n_512) );
NAND2x1_ASAP7_75t_L g513 ( .A(n_405), .B(n_350), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_441), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_443), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_408), .B(n_349), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_408), .B(n_349), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_409), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_425), .B(n_349), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_443), .B(n_344), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_394), .B(n_378), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_444), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_444), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_425), .B(n_334), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_426), .B(n_334), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_456), .B(n_433), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_456), .B(n_433), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_383), .B(n_344), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_426), .B(n_364), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_417), .B(n_347), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_463), .B(n_364), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_421), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_417), .B(n_347), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_384), .B(n_381), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_421), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_394), .B(n_378), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_388), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_463), .B(n_363), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_388), .B(n_381), .Y(n_539) );
INVxp67_ASAP7_75t_SL g540 ( .A(n_401), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_418), .Y(n_541) );
AO22x1_ASAP7_75t_L g542 ( .A1(n_405), .A2(n_363), .B1(n_378), .B2(n_52), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_418), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_462), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_431), .B(n_378), .Y(n_545) );
INVxp67_ASAP7_75t_SL g546 ( .A(n_404), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_437), .B(n_49), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_394), .B(n_50), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_437), .B(n_54), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_391), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_391), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_532), .B(n_411), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_492), .B(n_405), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_481), .B(n_394), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_468), .B(n_429), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_535), .B(n_412), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_526), .B(n_412), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_487), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_526), .B(n_411), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_467), .B(n_419), .Y(n_560) );
AND2x4_ASAP7_75t_SL g561 ( .A(n_519), .B(n_439), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_542), .A2(n_457), .B(n_440), .Y(n_562) );
NAND2xp33_ASAP7_75t_L g563 ( .A(n_475), .B(n_446), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_492), .Y(n_564) );
OA21x2_ASAP7_75t_L g565 ( .A1(n_473), .A2(n_416), .B(n_407), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_527), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_539), .B(n_422), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_483), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_471), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_469), .B(n_419), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_464), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_496), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_496), .Y(n_573) );
OAI21xp33_ASAP7_75t_L g574 ( .A1(n_530), .A2(n_432), .B(n_424), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_474), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_512), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_518), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_544), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_466), .B(n_455), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_478), .Y(n_580) );
AOI21xp5_ASAP7_75t_SL g581 ( .A1(n_475), .A2(n_439), .B(n_457), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_541), .B(n_445), .Y(n_582) );
OAI32xp33_ASAP7_75t_L g583 ( .A1(n_473), .A2(n_455), .A3(n_445), .B1(n_442), .B2(n_423), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_486), .A2(n_459), .B1(n_439), .B2(n_432), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_524), .B(n_432), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_543), .B(n_459), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_537), .B(n_404), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_486), .A2(n_439), .B1(n_423), .B2(n_424), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_525), .B(n_404), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_490), .B(n_407), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_513), .A2(n_462), .B1(n_409), .B2(n_450), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_477), .B(n_407), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_493), .B(n_438), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_498), .B(n_462), .Y(n_594) );
NOR2xp33_ASAP7_75t_SL g595 ( .A(n_547), .B(n_450), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_491), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_465), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_470), .B(n_450), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_516), .B(n_438), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_534), .B(n_452), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_470), .B(n_452), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_472), .B(n_452), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_501), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_504), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_476), .B(n_454), .Y(n_605) );
BUFx2_ASAP7_75t_SL g606 ( .A(n_548), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_545), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_503), .Y(n_608) );
AOI311xp33_ASAP7_75t_L g609 ( .A1(n_530), .A2(n_436), .A3(n_449), .B(n_448), .C(n_447), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_533), .A2(n_436), .B1(n_393), .B2(n_449), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_497), .B(n_454), .Y(n_611) );
BUFx2_ASAP7_75t_L g612 ( .A(n_503), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_479), .B(n_453), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_511), .B(n_448), .Y(n_614) );
INVx2_ASAP7_75t_SL g615 ( .A(n_479), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_505), .Y(n_616) );
NAND2x1p5_ASAP7_75t_L g617 ( .A(n_548), .B(n_447), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_597), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_584), .A2(n_533), .B1(n_495), .B2(n_517), .Y(n_619) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_588), .A2(n_549), .B(n_531), .Y(n_620) );
OAI22xp33_ASAP7_75t_SL g621 ( .A1(n_595), .A2(n_528), .B1(n_520), .B2(n_488), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_566), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_595), .B(n_500), .Y(n_623) );
AOI211x1_ASAP7_75t_L g624 ( .A1(n_583), .A2(n_488), .B(n_494), .C(n_520), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_567), .Y(n_625) );
AOI222xp33_ASAP7_75t_L g626 ( .A1(n_564), .A2(n_494), .B1(n_482), .B2(n_506), .C1(n_510), .C2(n_508), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_609), .B(n_499), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_553), .A2(n_507), .B1(n_509), .B2(n_514), .C(n_523), .Y(n_628) );
AOI21xp33_ASAP7_75t_L g629 ( .A1(n_574), .A2(n_489), .B(n_502), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_612), .B(n_500), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_558), .B(n_554), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_571), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_606), .A2(n_499), .B1(n_538), .B2(n_546), .Y(n_633) );
OAI21xp33_ASAP7_75t_L g634 ( .A1(n_557), .A2(n_529), .B(n_485), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_565), .B(n_515), .C(n_522), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g636 ( .A1(n_617), .A2(n_546), .B1(n_540), .B2(n_484), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_557), .A2(n_559), .B1(n_552), .B2(n_556), .C(n_579), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_575), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_580), .Y(n_639) );
OAI322xp33_ASAP7_75t_L g640 ( .A1(n_610), .A2(n_484), .A3(n_480), .B1(n_485), .B2(n_551), .C1(n_550), .C2(n_540), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_608), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_613), .B(n_536), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_559), .B(n_480), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_581), .A2(n_521), .B(n_414), .Y(n_644) );
INVxp67_ASAP7_75t_L g645 ( .A(n_569), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_608), .Y(n_646) );
INVxp67_ASAP7_75t_L g647 ( .A(n_572), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_596), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_573), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_556), .B(n_400), .Y(n_650) );
CKINVDCx14_ASAP7_75t_R g651 ( .A(n_560), .Y(n_651) );
OA21x2_ASAP7_75t_L g652 ( .A1(n_635), .A2(n_627), .B(n_647), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_641), .Y(n_653) );
OAI31xp33_ASAP7_75t_L g654 ( .A1(n_621), .A2(n_591), .A3(n_562), .B(n_615), .Y(n_654) );
AOI322xp5_ASAP7_75t_L g655 ( .A1(n_651), .A2(n_570), .A3(n_563), .B1(n_585), .B2(n_589), .C1(n_590), .C2(n_586), .Y(n_655) );
OAI21xp5_ASAP7_75t_SL g656 ( .A1(n_620), .A2(n_591), .B(n_561), .Y(n_656) );
XOR2x2_ASAP7_75t_L g657 ( .A(n_633), .B(n_599), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_619), .A2(n_555), .B1(n_605), .B2(n_602), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_622), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_623), .A2(n_587), .B(n_592), .Y(n_660) );
AOI221x1_ASAP7_75t_L g661 ( .A1(n_621), .A2(n_616), .B1(n_603), .B2(n_604), .C(n_613), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_624), .A2(n_598), .B1(n_601), .B2(n_587), .C(n_611), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_626), .A2(n_593), .B1(n_582), .B2(n_607), .Y(n_663) );
O2A1O1Ixp33_ASAP7_75t_SL g664 ( .A1(n_645), .A2(n_646), .B(n_636), .C(n_629), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_618), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_637), .B(n_568), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_640), .A2(n_592), .B(n_614), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_643), .B(n_600), .Y(n_668) );
NAND4xp25_ASAP7_75t_L g669 ( .A(n_644), .B(n_614), .C(n_594), .D(n_438), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_634), .A2(n_565), .B1(n_577), .B2(n_576), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g671 ( .A1(n_631), .A2(n_578), .B(n_453), .C(n_59), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_625), .A2(n_56), .B1(n_57), .B2(n_61), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_628), .B(n_62), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_640), .A2(n_64), .B(n_65), .Y(n_674) );
AOI222xp33_ASAP7_75t_L g675 ( .A1(n_632), .A2(n_68), .B1(n_69), .B2(n_72), .C1(n_73), .C2(n_74), .Y(n_675) );
AO22x1_ASAP7_75t_L g676 ( .A1(n_630), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_638), .B(n_639), .Y(n_677) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_649), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_642), .B(n_650), .Y(n_679) );
AOI211xp5_ASAP7_75t_L g680 ( .A1(n_642), .A2(n_627), .B(n_621), .C(n_633), .Y(n_680) );
OAI221xp5_ASAP7_75t_SL g681 ( .A1(n_648), .A2(n_620), .B1(n_619), .B2(n_651), .C(n_584), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_680), .B(n_652), .C(n_654), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_659), .Y(n_683) );
OAI21xp33_ASAP7_75t_SL g684 ( .A1(n_655), .A2(n_669), .B(n_679), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_652), .B(n_681), .C(n_664), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_677), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_665), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_683), .Y(n_688) );
AND5x1_ASAP7_75t_L g689 ( .A(n_684), .B(n_674), .C(n_670), .D(n_663), .E(n_671), .Y(n_689) );
NAND4xp25_ASAP7_75t_SL g690 ( .A(n_685), .B(n_661), .C(n_667), .D(n_666), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_686), .B(n_662), .Y(n_691) );
NOR2x1_ASAP7_75t_L g692 ( .A(n_690), .B(n_682), .Y(n_692) );
AND2x4_ASAP7_75t_L g693 ( .A(n_689), .B(n_653), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_691), .B(n_687), .Y(n_694) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_694), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_692), .Y(n_696) );
AO22x2_ASAP7_75t_L g697 ( .A1(n_696), .A2(n_693), .B1(n_688), .B2(n_656), .Y(n_697) );
OAI22x1_ASAP7_75t_L g698 ( .A1(n_695), .A2(n_678), .B1(n_672), .B2(n_673), .Y(n_698) );
INVx3_ASAP7_75t_L g699 ( .A(n_697), .Y(n_699) );
AOI21xp33_ASAP7_75t_SL g700 ( .A1(n_699), .A2(n_698), .B(n_675), .Y(n_700) );
OAI21xp5_ASAP7_75t_L g701 ( .A1(n_700), .A2(n_699), .B(n_657), .Y(n_701) );
OR2x6_ASAP7_75t_L g702 ( .A(n_701), .B(n_676), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_702), .A2(n_658), .B1(n_668), .B2(n_660), .Y(n_703) );
endmodule