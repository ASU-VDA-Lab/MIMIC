module fake_jpeg_3418_n_236 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_7),
.B(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_47),
.B(n_50),
.Y(n_92)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_15),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_0),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_75),
.Y(n_80)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_40),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g105 ( 
.A(n_57),
.Y(n_105)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_59),
.B(n_65),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_32),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_42),
.B1(n_33),
.B2(n_31),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_21),
.B(n_12),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_2),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_71),
.Y(n_89)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_3),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_21),
.B(n_14),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_72),
.B(n_61),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_3),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_74),
.B(n_35),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_29),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_23),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_33),
.B1(n_31),
.B2(n_27),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_78),
.A2(n_117),
.B1(n_104),
.B2(n_102),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_82),
.A2(n_90),
.B1(n_101),
.B2(n_105),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_26),
.B1(n_27),
.B2(n_23),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_84),
.A2(n_94),
.B1(n_99),
.B2(n_106),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_90),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_44),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_4),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_4),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_4),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_100),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_44),
.A2(n_35),
.B1(n_18),
.B2(n_20),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_5),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_5),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_63),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_56),
.A2(n_35),
.B1(n_18),
.B2(n_20),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_5),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_118),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_70),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_53),
.A2(n_54),
.B1(n_66),
.B2(n_67),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_131),
.Y(n_158)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_80),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_139),
.Y(n_150)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_92),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_141),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_89),
.A2(n_87),
.B1(n_103),
.B2(n_79),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_138),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_88),
.A2(n_78),
.B(n_93),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_91),
.B(n_139),
.Y(n_161)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_87),
.A2(n_108),
.B(n_97),
.C(n_105),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_142),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_113),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_111),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_144),
.A2(n_116),
.B1(n_109),
.B2(n_91),
.Y(n_149)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_146),
.Y(n_156)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_104),
.B1(n_81),
.B2(n_107),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_148),
.B1(n_120),
.B2(n_145),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_147),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_153),
.B1(n_166),
.B2(n_138),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_116),
.B1(n_111),
.B2(n_109),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_124),
.Y(n_185)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_91),
.B1(n_137),
.B2(n_134),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_167),
.B1(n_158),
.B2(n_159),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_137),
.A2(n_136),
.B1(n_133),
.B2(n_120),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_123),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_122),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_177),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_123),
.C(n_126),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_184),
.C(n_127),
.Y(n_187)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_173),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_130),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_176),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_155),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_128),
.Y(n_178)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_121),
.B(n_125),
.C(n_146),
.D(n_154),
.Y(n_197)
);

OAI21x1_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_182),
.B(n_185),
.Y(n_194)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

INVx4_ASAP7_75t_SL g181 ( 
.A(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_167),
.B1(n_158),
.B2(n_162),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_119),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_183),
.A2(n_163),
.B(n_156),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_135),
.C(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_151),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_184),
.C(n_180),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_159),
.B(n_166),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_188),
.A2(n_195),
.B(n_197),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_169),
.B(n_168),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_196),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_168),
.B(n_163),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_151),
.B(n_152),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_182),
.B1(n_175),
.B2(n_181),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_204),
.A2(n_207),
.B1(n_188),
.B2(n_195),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_175),
.B1(n_176),
.B2(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_208),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_181),
.B1(n_172),
.B2(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_209),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_193),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_177),
.B1(n_152),
.B2(n_143),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_191),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_216),
.Y(n_222)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_215),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_191),
.A3(n_187),
.B1(n_211),
.B2(n_203),
.C1(n_197),
.C2(n_210),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_218),
.C(n_203),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_221),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_193),
.C(n_204),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_210),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_224),
.B(n_219),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_222),
.A2(n_214),
.B1(n_215),
.B2(n_206),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_206),
.B(n_219),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_226),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_232),
.B1(n_223),
.B2(n_226),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_230),
.B(n_227),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_234),
.A2(n_231),
.B1(n_228),
.B2(n_143),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_173),
.Y(n_236)
);


endmodule