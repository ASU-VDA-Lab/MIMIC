module real_jpeg_20585_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_255;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_0),
.A2(n_28),
.B1(n_31),
.B2(n_48),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_1),
.A2(n_46),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_1),
.A2(n_28),
.B1(n_31),
.B2(n_46),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_2),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_2),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_2),
.A2(n_56),
.B1(n_57),
.B2(n_75),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_2),
.A2(n_28),
.B1(n_31),
.B2(n_75),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_75),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_3),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_4),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_4),
.A2(n_32),
.B1(n_56),
.B2(n_57),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_4),
.A2(n_32),
.B1(n_39),
.B2(n_40),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_5),
.A2(n_69),
.B1(n_74),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_5),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_136),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_136),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_5),
.A2(n_28),
.B1(n_31),
.B2(n_136),
.Y(n_193)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_6),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_6),
.A2(n_26),
.B(n_127),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_6),
.A2(n_177),
.B1(n_178),
.B2(n_180),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_7),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_7),
.A2(n_36),
.B1(n_69),
.B2(n_74),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_7),
.A2(n_36),
.B1(n_56),
.B2(n_57),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_7),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_149)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_9),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_9),
.A2(n_14),
.B(n_28),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_9),
.A2(n_39),
.B1(n_40),
.B2(n_124),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_9),
.A2(n_27),
.B1(n_193),
.B2(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_9),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_9),
.B(n_56),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_9),
.A2(n_56),
.B(n_220),
.Y(n_224)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_11),
.A2(n_69),
.B1(n_74),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_11),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_11),
.A2(n_56),
.B1(n_57),
.B2(n_109),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_11),
.A2(n_28),
.B1(n_31),
.B2(n_109),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_109),
.Y(n_211)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_13),
.A2(n_56),
.B1(n_57),
.B2(n_68),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_14),
.A2(n_39),
.B(n_42),
.C(n_43),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_39),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_14),
.A2(n_28),
.B1(n_31),
.B2(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_15),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_139),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_137),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_19),
.B(n_111),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_89),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_79),
.B2(n_80),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_49),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_24),
.B(n_37),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_27),
.A2(n_29),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_27),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_27),
.A2(n_98),
.B1(n_101),
.B2(n_126),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_27),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_27),
.A2(n_101),
.B1(n_179),
.B2(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_27),
.A2(n_33),
.B(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_29),
.B(n_124),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_30),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_31),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_34),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_35),
.A2(n_100),
.B(n_177),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_38),
.A2(n_47),
.B(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_38),
.A2(n_85),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_38),
.A2(n_43),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_38),
.A2(n_43),
.B1(n_189),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_38),
.A2(n_43),
.B1(n_211),
.B2(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_38),
.A2(n_227),
.B(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_40),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

AOI32xp33_ASAP7_75t_L g219 ( 
.A1(n_39),
.A2(n_54),
.A3(n_57),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_40),
.A2(n_44),
.B(n_124),
.C(n_185),
.Y(n_184)
);

NAND2xp33_ASAP7_75t_SL g221 ( 
.A(n_40),
.B(n_52),
.Y(n_221)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_43),
.A2(n_45),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_43),
.B(n_124),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_64),
.B1(n_65),
.B2(n_78),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_50),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B(n_58),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_52),
.B(n_56),
.C(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_63),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_51),
.B(n_104),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_51),
.A2(n_60),
.B1(n_130),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_51),
.A2(n_60),
.B1(n_152),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_51),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_51),
.A2(n_60),
.B1(n_165),
.B2(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_56),
.Y(n_61)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_68),
.Y(n_122)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_57),
.A2(n_71),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_59),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_59),
.A2(n_129),
.B(n_131),
.Y(n_128)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_73),
.B(n_76),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_73),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_66),
.A2(n_108),
.B1(n_110),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_67),
.A2(n_72),
.B1(n_123),
.B2(n_135),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_71),
.C(n_72),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g123 ( 
.A(n_69),
.B(n_124),
.CON(n_123),
.SN(n_123)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_88),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_87),
.B(n_149),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_102),
.C(n_106),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_91),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_106),
.B1(n_107),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_110),
.B(n_124),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_118),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_112),
.A2(n_116),
.B1(n_117),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_112),
.Y(n_257)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_118),
.A2(n_119),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_128),
.C(n_132),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_125),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_132),
.B1(n_133),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_169),
.B(n_252),
.C(n_258),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_158),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_141),
.B(n_158),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_154),
.B2(n_157),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_144),
.B(n_145),
.C(n_157),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_153),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_153),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_159),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_163),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_167),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_164),
.B(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_166),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_251),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_245),
.B(n_250),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_232),
.B(n_244),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_214),
.B(n_231),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_202),
.B(n_213),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_190),
.B(n_201),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_182),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_182),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_186),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_195),
.B(n_200),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_194),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_203),
.B(n_204),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_212),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_210),
.C(n_212),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_216),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_222),
.B1(n_229),
.B2(n_230),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_217),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_223),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_233),
.B(n_234),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_241),
.C(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_254),
.Y(n_258)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);


endmodule