module real_jpeg_16904_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_572;
wire n_405;
wire n_412;
wire n_548;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_1),
.Y(n_106)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_1),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_3),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_3),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_3),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_3),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_4),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_4),
.A2(n_52),
.B1(n_96),
.B2(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_4),
.A2(n_52),
.B1(n_205),
.B2(n_209),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_4),
.A2(n_52),
.B1(n_261),
.B2(n_266),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_5),
.A2(n_48),
.B1(n_121),
.B2(n_124),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_5),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_5),
.A2(n_124),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_5),
.A2(n_124),
.B1(n_273),
.B2(n_277),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_5),
.A2(n_124),
.B1(n_339),
.B2(n_342),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_6),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_6),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_6),
.A2(n_129),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_6),
.A2(n_129),
.B1(n_238),
.B2(n_241),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_6),
.A2(n_129),
.B1(n_351),
.B2(n_354),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_7),
.Y(n_220)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_7),
.Y(n_349)
);

BUFx5_ASAP7_75t_L g405 ( 
.A(n_7),
.Y(n_405)
);

BUFx5_ASAP7_75t_L g497 ( 
.A(n_7),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_8),
.A2(n_127),
.B1(n_306),
.B2(n_308),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_8),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_8),
.A2(n_308),
.B1(n_395),
.B2(n_397),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_8),
.A2(n_205),
.B1(n_308),
.B2(n_451),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_8),
.A2(n_308),
.B1(n_490),
.B2(n_493),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_43),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_9),
.A2(n_38),
.B1(n_89),
.B2(n_92),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_9),
.A2(n_38),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_9),
.A2(n_38),
.B1(n_226),
.B2(n_229),
.Y(n_225)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_10),
.Y(n_150)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_10),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_10),
.Y(n_240)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_10),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_10),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_10),
.Y(n_469)
);

BUFx5_ASAP7_75t_L g524 ( 
.A(n_10),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_11),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_11),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_11),
.A2(n_169),
.B1(n_285),
.B2(n_318),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_11),
.A2(n_285),
.B1(n_456),
.B2(n_457),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g517 ( 
.A1(n_11),
.A2(n_285),
.B1(n_518),
.B2(n_520),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_12),
.Y(n_313)
);

OAI32xp33_ASAP7_75t_L g322 ( 
.A1(n_13),
.A2(n_126),
.A3(n_323),
.B1(n_325),
.B2(n_331),
.Y(n_322)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_13),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_13),
.A2(n_43),
.B1(n_330),
.B2(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_13),
.B(n_27),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_13),
.B(n_77),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_13),
.B(n_133),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_13),
.B(n_507),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_SL g526 ( 
.A1(n_13),
.A2(n_326),
.B1(n_330),
.B2(n_365),
.Y(n_526)
);

OAI32xp33_ASAP7_75t_L g528 ( 
.A1(n_13),
.A2(n_529),
.A3(n_532),
.B1(n_535),
.B2(n_536),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_15),
.Y(n_117)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_16),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_16),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_16),
.Y(n_265)
);

BUFx4f_ASAP7_75t_L g505 ( 
.A(n_16),
.Y(n_505)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_579),
.Y(n_22)
);

OAI221xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_65),
.B1(n_68),
.B2(n_294),
.C(n_573),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_24),
.B(n_65),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_25),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_25),
.B(n_70),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_46),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_26),
.A2(n_58),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_37),
.Y(n_26)
);

OR2x6_ASAP7_75t_L g58 ( 
.A(n_27),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_27),
.B(n_47),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_27),
.A2(n_57),
.B1(n_304),
.B2(n_309),
.Y(n_303)
);

AO22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_29),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_30),
.Y(n_176)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_31),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_33),
.Y(n_531)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_41),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_43),
.Y(n_130)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_45),
.Y(n_286)
);

OAI21x1_ASAP7_75t_SL g165 ( 
.A1(n_46),
.A2(n_66),
.B(n_120),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_57),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_50),
.Y(n_307)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_51),
.Y(n_312)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_56),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_66),
.B(n_67),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_58),
.A2(n_66),
.B1(n_120),
.B2(n_125),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_58),
.A2(n_125),
.B(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_58),
.A2(n_67),
.B(n_157),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_58),
.A2(n_66),
.B1(n_305),
.B2(n_361),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_58),
.A2(n_66),
.B1(n_282),
.B2(n_310),
.Y(n_383)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_160),
.C(n_180),
.Y(n_68)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g573 ( 
.A1(n_69),
.A2(n_160),
.B(n_574),
.C(n_577),
.D(n_578),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_156),
.C(n_158),
.Y(n_70)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_71),
.B(n_156),
.CI(n_158),
.CON(n_179),
.SN(n_179)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_118),
.C(n_131),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_72),
.A2(n_73),
.B1(n_131),
.B2(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_94),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_75),
.A2(n_101),
.B(n_316),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_88),
.Y(n_75)
);

OAI22x1_ASAP7_75t_L g288 ( 
.A1(n_76),
.A2(n_102),
.B1(n_195),
.B2(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_76),
.A2(n_102),
.B1(n_317),
.B2(n_364),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_76),
.A2(n_102),
.B1(n_364),
.B2(n_394),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_76),
.A2(n_102),
.B1(n_394),
.B2(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_103),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_77),
.A2(n_101),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_77),
.B(n_95),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_77),
.A2(n_101),
.B1(n_168),
.B2(n_194),
.Y(n_193)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_84),
.B2(n_86),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_81),
.A2(n_145),
.B1(n_146),
.B2(n_148),
.Y(n_144)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_83),
.Y(n_211)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_83),
.Y(n_276)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_88),
.A2(n_102),
.B(n_178),
.Y(n_384)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_89),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_90),
.Y(n_320)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_95),
.Y(n_289)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_97),
.Y(n_396)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21x1_ASAP7_75t_SL g167 ( 
.A1(n_101),
.A2(n_168),
.B(n_177),
.Y(n_167)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_109),
.B2(n_114),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_117),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_117),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_122),
.A2(n_311),
.B1(n_313),
.B2(n_314),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_165),
.C(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_132),
.B(n_167),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_143),
.B(n_151),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_133),
.B(n_204),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_133),
.B(n_272),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_133),
.A2(n_143),
.B1(n_445),
.B2(n_450),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_133),
.A2(n_143),
.B1(n_450),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_134),
.B(n_152),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_134),
.A2(n_237),
.B1(n_242),
.B2(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_134),
.A2(n_242),
.B1(n_516),
.B2(n_517),
.Y(n_515)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_138),
.B1(n_140),
.B2(n_142),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_136),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_137),
.Y(n_224)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_140),
.Y(n_456)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_141),
.Y(n_228)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_141),
.Y(n_344)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_141),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_141),
.Y(n_481)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_141),
.Y(n_492)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_142),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_143),
.B(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_143),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_143),
.A2(n_201),
.B(n_558),
.Y(n_557)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_149),
.Y(n_452)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_150),
.Y(n_435)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_151),
.Y(n_359)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_155),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_179),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_161),
.B(n_179),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.C(n_166),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_165),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_185),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_176),
.Y(n_199)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_176),
.Y(n_367)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g581 ( 
.A(n_179),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_246),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_181),
.A2(n_575),
.B(n_576),
.Y(n_574)
);

NOR2xp67_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_182),
.B(n_186),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.C(n_212),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_188),
.A2(n_191),
.B1(n_192),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_188),
.Y(n_293)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_189),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

OA21x2_ASAP7_75t_SL g250 ( 
.A1(n_192),
.A2(n_200),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_200),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_203),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_205),
.B(n_330),
.Y(n_440)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_212),
.A2(n_213),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_233),
.B(n_244),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_215),
.B1(n_244),
.B2(n_245),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_214),
.A2(n_215),
.B1(n_236),
.B2(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_221),
.B(n_225),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_222),
.Y(n_221)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_220),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_221),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_221),
.Y(n_337)
);

AOI21x1_ASAP7_75t_L g454 ( 
.A1(n_221),
.A2(n_455),
.B(n_462),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_221),
.A2(n_475),
.B1(n_489),
.B2(n_494),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_221),
.A2(n_330),
.B1(n_489),
.B2(n_496),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_222),
.Y(n_493)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_224),
.Y(n_341)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_224),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_225),
.Y(n_546)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_232),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_236),
.Y(n_414)
);

OA21x2_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_242),
.B(n_243),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_242),
.A2(n_243),
.B(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_290),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_247),
.B(n_290),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.C(n_252),
.Y(n_247)
);

XNOR2x1_ASAP7_75t_L g424 ( 
.A(n_248),
.B(n_250),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_252),
.B(n_424),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_281),
.C(n_287),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g415 ( 
.A(n_253),
.B(n_416),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_270),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_254),
.B(n_270),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_259),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_255),
.Y(n_462)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_259),
.A2(n_338),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_260),
.B(n_371),
.Y(n_370)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_264),
.Y(n_269)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_264),
.Y(n_461)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_276),
.Y(n_534)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2x1_ASAP7_75t_L g416 ( 
.A(n_281),
.B(n_288),
.Y(n_416)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_567),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_425),
.Y(n_296)
);

NOR3xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_408),
.C(n_421),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_386),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_375),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_300),
.B(n_375),
.C(n_569),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_357),
.C(n_368),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_301),
.B(n_407),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_321),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_315),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_303),
.B(n_315),
.C(n_321),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_311),
.Y(n_362)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_313),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_313),
.A2(n_314),
.B1(n_318),
.B2(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_313),
.A2(n_314),
.B1(n_466),
.B2(n_468),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_313),
.A2(n_314),
.B1(n_476),
.B2(n_480),
.Y(n_475)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_336),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_322),
.B(n_336),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_329),
.Y(n_398)
);

OAI21xp33_ASAP7_75t_SL g445 ( 
.A1(n_330),
.A2(n_440),
.B(n_446),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_330),
.B(n_432),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_345),
.B2(n_350),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_337),
.A2(n_350),
.B(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_337),
.A2(n_474),
.B1(n_482),
.B2(n_483),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_337),
.A2(n_370),
.B(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_344),
.Y(n_356)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_348),
.Y(n_372)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_357),
.B(n_368),
.Y(n_407)
);

MAJx2_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.C(n_363),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_363),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_360),
.B(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_SL g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_373),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_373),
.Y(n_381)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_376),
.B(n_379),
.C(n_385),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_380),
.B2(n_385),
.Y(n_377)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_378),
.Y(n_385)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_R g418 ( 
.A(n_381),
.B(n_383),
.C(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_384),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_406),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_387),
.B(n_406),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_390),
.C(n_392),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_388),
.B(n_563),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_390),
.A2(n_391),
.B1(n_392),
.B2(n_564),
.Y(n_563)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_392),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_399),
.C(n_401),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g552 ( 
.A(n_393),
.B(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_399),
.A2(n_400),
.B1(n_401),
.B2(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_401),
.Y(n_554)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g567 ( 
.A1(n_409),
.A2(n_568),
.B(n_570),
.C(n_571),
.D(n_572),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_410),
.B(n_411),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_417),
.B1(n_418),
.B2(n_420),
.Y(n_411)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_412),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_415),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_413),
.B(n_415),
.C(n_417),
.Y(n_422)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_421),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_422),
.B(n_423),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_561),
.B(n_566),
.Y(n_425)
);

AOI21x1_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_548),
.B(n_560),
.Y(n_426)
);

OAI21x1_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_511),
.B(n_547),
.Y(n_427)
);

AOI21x1_ASAP7_75t_SL g428 ( 
.A1(n_429),
.A2(n_471),
.B(n_510),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_453),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_430),
.B(n_453),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_443),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_431),
.A2(n_443),
.B1(n_444),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_431),
.Y(n_485)
);

OAI32xp33_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_436),
.A3(n_438),
.B1(n_440),
.B2(n_441),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_437),
.B(n_442),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_463),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_454),
.B(n_464),
.C(n_470),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_455),
.Y(n_482)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_470),
.Y(n_463)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_465),
.Y(n_516)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_468),
.Y(n_519)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_472),
.A2(n_486),
.B(n_509),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_484),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_473),
.B(n_484),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

AOI21x1_ASAP7_75t_L g486 ( 
.A1(n_487),
.A2(n_499),
.B(n_508),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_488),
.B(n_498),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_488),
.B(n_498),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx6_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

BUFx12f_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_500),
.B(n_501),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_506),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_513),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_512),
.B(n_513),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_527),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_525),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_515),
.B(n_525),
.C(n_527),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_517),
.Y(n_558)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_545),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_528),
.B(n_545),
.Y(n_556)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_540),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_550),
.Y(n_548)
);

NOR2xp67_ASAP7_75t_SL g560 ( 
.A(n_549),
.B(n_550),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_551),
.A2(n_552),
.B1(n_555),
.B2(n_559),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_551),
.B(n_556),
.C(n_557),
.Y(n_565)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_555),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_557),
.Y(n_555)
);

NOR2xp67_ASAP7_75t_SL g561 ( 
.A(n_562),
.B(n_565),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_562),
.B(n_565),
.Y(n_566)
);


endmodule