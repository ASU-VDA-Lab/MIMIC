module fake_jpeg_1441_n_682 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_682);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_682;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_540;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_587;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g161 ( 
.A(n_60),
.Y(n_161)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_61),
.Y(n_211)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_10),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_63),
.B(n_64),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_11),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_29),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_65),
.A2(n_27),
.B(n_55),
.Y(n_147)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_66),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_67),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_29),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_69),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_70),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_71),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_22),
.B(n_8),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_72),
.B(n_75),
.Y(n_133)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_74),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_76),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_77),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_78),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_79),
.Y(n_217)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_81),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_21),
.B(n_8),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_86),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_33),
.B(n_8),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_83),
.B(n_89),
.Y(n_146)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_85),
.Y(n_222)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_87),
.Y(n_218)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_88),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_36),
.B(n_12),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_37),
.B(n_12),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_109),
.Y(n_148)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_95),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_97),
.Y(n_224)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_106),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_28),
.Y(n_101)
);

BUFx24_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_102),
.Y(n_190)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_28),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_111),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_21),
.B(n_12),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_110),
.Y(n_225)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_44),
.Y(n_115)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_123),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_59),
.B(n_12),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_58),
.Y(n_165)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_57),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_126),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_57),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_127),
.B(n_47),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_128),
.Y(n_189)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_34),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_39),
.Y(n_130)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_39),
.Y(n_131)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

BUFx16f_ASAP7_75t_L g132 ( 
.A(n_34),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_132),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_143),
.B(n_163),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_147),
.A2(n_174),
.B1(n_179),
.B2(n_197),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_72),
.B(n_27),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_165),
.B(n_167),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_68),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_84),
.B(n_32),
.C(n_47),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_169),
.B(n_202),
.C(n_210),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_70),
.A2(n_47),
.B1(n_56),
.B2(n_58),
.Y(n_174)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_176),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_61),
.B(n_52),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_178),
.B(n_188),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_71),
.A2(n_34),
.B1(n_50),
.B2(n_52),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_76),
.A2(n_56),
.B1(n_55),
.B2(n_49),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_184),
.A2(n_125),
.B1(n_0),
.B2(n_3),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_101),
.B(n_35),
.Y(n_188)
);

HAxp5_ASAP7_75t_SL g193 ( 
.A(n_65),
.B(n_50),
.CON(n_193),
.SN(n_193)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_193),
.B(n_195),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_77),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_199),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_62),
.B(n_49),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_79),
.A2(n_43),
.B1(n_41),
.B2(n_40),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_73),
.Y(n_198)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_100),
.B(n_43),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_96),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_200),
.B(n_201),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_97),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_90),
.B(n_50),
.C(n_34),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_95),
.Y(n_203)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_60),
.B(n_35),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_206),
.B(n_207),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_131),
.B(n_60),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_99),
.Y(n_209)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_87),
.A2(n_41),
.B1(n_40),
.B2(n_50),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_115),
.B(n_50),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_119),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_130),
.B(n_34),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_214),
.B(n_219),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_88),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_215),
.A2(n_119),
.B1(n_78),
.B2(n_113),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_108),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_110),
.Y(n_220)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_220),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_102),
.B(n_19),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_223),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_116),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_118),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_229),
.Y(n_275)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_122),
.Y(n_228)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_228),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_129),
.B(n_19),
.Y(n_229)
);

BUFx16f_ASAP7_75t_L g231 ( 
.A(n_136),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_231),
.Y(n_341)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_145),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_232),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_152),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_234),
.B(n_242),
.Y(n_329)
);

CKINVDCx12_ASAP7_75t_R g235 ( 
.A(n_150),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_235),
.Y(n_373)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_236),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_237),
.B(n_298),
.Y(n_321)
);

INVx13_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_238),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_240),
.A2(n_267),
.B1(n_290),
.B2(n_307),
.Y(n_314)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_150),
.Y(n_241)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_241),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_159),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_145),
.Y(n_243)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_243),
.Y(n_347)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_150),
.Y(n_246)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_246),
.Y(n_357)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_247),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_179),
.A2(n_78),
.B1(n_112),
.B2(n_105),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_248),
.A2(n_293),
.B1(n_294),
.B2(n_310),
.Y(n_315)
);

CKINVDCx12_ASAP7_75t_R g250 ( 
.A(n_134),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_250),
.Y(n_326)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_160),
.Y(n_251)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_251),
.Y(n_313)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_153),
.Y(n_252)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_252),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_180),
.Y(n_254)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_254),
.Y(n_319)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_175),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_255),
.Y(n_330)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_257),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_204),
.Y(n_259)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_259),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_260),
.A2(n_308),
.B1(n_161),
.B2(n_173),
.Y(n_323)
);

INVx8_ASAP7_75t_L g261 ( 
.A(n_156),
.Y(n_261)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_261),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_168),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_262),
.B(n_300),
.Y(n_369)
);

CKINVDCx12_ASAP7_75t_R g264 ( 
.A(n_207),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_264),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_174),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_133),
.B(n_148),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_268),
.B(n_271),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_146),
.B(n_181),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_0),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_272),
.B(n_280),
.Y(n_352)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_187),
.Y(n_273)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_273),
.Y(n_362)
);

CKINVDCx6p67_ASAP7_75t_R g274 ( 
.A(n_158),
.Y(n_274)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

INVx3_ASAP7_75t_SL g276 ( 
.A(n_153),
.Y(n_276)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_276),
.Y(n_372)
);

BUFx4f_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_277),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_142),
.B(n_14),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_285),
.Y(n_318)
);

CKINVDCx6p67_ASAP7_75t_R g279 ( 
.A(n_158),
.Y(n_279)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_279),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_169),
.B(n_0),
.Y(n_280)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_191),
.Y(n_282)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_282),
.Y(n_317)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_172),
.Y(n_284)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_139),
.B(n_151),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_211),
.Y(n_286)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_204),
.Y(n_287)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_287),
.Y(n_368)
);

INVx3_ASAP7_75t_SL g288 ( 
.A(n_190),
.Y(n_288)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_288),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_202),
.B(n_0),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_289),
.B(n_301),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_197),
.A2(n_14),
.B1(n_3),
.B2(n_4),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_166),
.Y(n_291)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_291),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_135),
.B(n_15),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_295),
.Y(n_327)
);

CKINVDCx6p67_ASAP7_75t_R g293 ( 
.A(n_161),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_193),
.A2(n_208),
.B1(n_173),
.B2(n_226),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_218),
.B(n_5),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_192),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_296),
.B(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_155),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_166),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_149),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_147),
.B(n_0),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_149),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_302),
.B(n_303),
.Y(n_343)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_192),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_157),
.B(n_13),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_R g359 ( 
.A(n_304),
.B(n_156),
.Y(n_359)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_140),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_305),
.B(n_306),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_218),
.B(n_14),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_184),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_210),
.A2(n_16),
.B1(n_17),
.B2(n_215),
.Y(n_308)
);

CKINVDCx12_ASAP7_75t_R g309 ( 
.A(n_161),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_312),
.Y(n_334)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_183),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_185),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_311),
.A2(n_189),
.B1(n_216),
.B2(n_162),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_226),
.B(n_190),
.Y(n_312)
);

AOI22x1_ASAP7_75t_L g322 ( 
.A1(n_301),
.A2(n_140),
.B1(n_186),
.B2(n_164),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_322),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_323),
.A2(n_332),
.B1(n_274),
.B2(n_279),
.Y(n_377)
);

AO22x1_ASAP7_75t_SL g324 ( 
.A1(n_308),
.A2(n_185),
.B1(n_170),
.B2(n_171),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_324),
.B(n_335),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_283),
.A2(n_154),
.B1(n_217),
.B2(n_212),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_325),
.A2(n_340),
.B1(n_345),
.B2(n_349),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_249),
.A2(n_208),
.B(n_182),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_SL g331 ( 
.A(n_249),
.B(n_189),
.C(n_182),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_331),
.B(n_367),
.C(n_349),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_283),
.A2(n_217),
.B1(n_212),
.B2(n_205),
.Y(n_332)
);

AO22x1_ASAP7_75t_SL g335 ( 
.A1(n_260),
.A2(n_137),
.B1(n_138),
.B2(n_177),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_299),
.A2(n_186),
.B1(n_137),
.B2(n_138),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_342),
.A2(n_360),
.B1(n_279),
.B2(n_293),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_299),
.A2(n_154),
.B1(n_205),
.B2(n_225),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_230),
.A2(n_191),
.B1(n_164),
.B2(n_144),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_346),
.Y(n_388)
);

OAI22x1_ASAP7_75t_L g349 ( 
.A1(n_280),
.A2(n_189),
.B1(n_216),
.B2(n_144),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_253),
.B(n_216),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_350),
.B(n_274),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_266),
.A2(n_225),
.B1(n_141),
.B2(n_196),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_353),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_272),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_275),
.A2(n_224),
.B1(n_141),
.B2(n_196),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_289),
.A2(n_156),
.B(n_162),
.Y(n_363)
);

AOI21xp33_ASAP7_75t_L g393 ( 
.A1(n_363),
.A2(n_274),
.B(n_279),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_258),
.A2(n_162),
.B(n_177),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_369),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_375),
.B(n_400),
.Y(n_429)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_376),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_377),
.A2(n_325),
.B1(n_363),
.B2(n_332),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_378),
.Y(n_439)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_343),
.Y(n_380)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_380),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_270),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_381),
.B(n_387),
.Y(n_446)
);

BUFx24_ASAP7_75t_SL g383 ( 
.A(n_320),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_383),
.B(n_396),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_384),
.A2(n_393),
.B(n_334),
.Y(n_426)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_385),
.Y(n_440)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_372),
.Y(n_386)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_386),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_263),
.Y(n_387)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_372),
.Y(n_389)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_389),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_351),
.B(n_268),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_390),
.B(n_407),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_352),
.B(n_271),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_391),
.B(n_398),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_351),
.B(n_237),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g459 ( 
.A(n_394),
.B(n_303),
.C(n_245),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_395),
.A2(n_405),
.B1(n_417),
.B2(n_423),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g396 ( 
.A(n_331),
.B(n_239),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_397),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_352),
.B(n_304),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_333),
.Y(n_399)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_399),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_330),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_366),
.B(n_265),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_401),
.B(n_406),
.Y(n_456)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_403),
.Y(n_432)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_404),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_359),
.A2(n_244),
.B1(n_298),
.B2(n_291),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_281),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_321),
.B(n_281),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_338),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_408),
.B(n_410),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_409),
.Y(n_438)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_338),
.Y(n_410)
);

INVx8_ASAP7_75t_L g411 ( 
.A(n_336),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_411),
.B(n_413),
.Y(n_452)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_371),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_355),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_414),
.B(n_415),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_327),
.B(n_252),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_321),
.B(n_256),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_370),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g417 ( 
.A1(n_314),
.A2(n_245),
.B1(n_310),
.B2(n_233),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_326),
.B(n_231),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_418),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_345),
.A2(n_293),
.B1(n_277),
.B2(n_282),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_419),
.A2(n_373),
.B1(n_374),
.B2(n_277),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_361),
.B(n_231),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_421),
.A2(n_422),
.B(n_341),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_321),
.B(n_293),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_355),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_424),
.A2(n_451),
.B1(n_392),
.B2(n_388),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_394),
.B(n_328),
.C(n_350),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_425),
.B(n_428),
.C(n_435),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_426),
.A2(n_443),
.B(n_463),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_367),
.C(n_313),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_430),
.B(n_453),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_431),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_420),
.A2(n_322),
.B1(n_323),
.B2(n_315),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_433),
.A2(n_450),
.B1(n_455),
.B2(n_379),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_398),
.B(n_334),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_401),
.B(n_339),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_436),
.B(n_449),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_384),
.A2(n_353),
.B(n_346),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_391),
.B(n_354),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_420),
.A2(n_322),
.B1(n_335),
.B2(n_324),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_382),
.A2(n_335),
.B1(n_324),
.B2(n_232),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g453 ( 
.A1(n_382),
.A2(n_317),
.B(n_365),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_388),
.A2(n_368),
.B1(n_337),
.B2(n_319),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_377),
.A2(n_357),
.B1(n_373),
.B2(n_316),
.Y(n_457)
);

BUFx12f_ASAP7_75t_L g484 ( 
.A(n_457),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_458),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_459),
.B(n_397),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_SL g463 ( 
.A1(n_409),
.A2(n_357),
.B1(n_316),
.B2(n_358),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_464),
.B(n_375),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_465),
.B(n_468),
.Y(n_503)
);

A2O1A1O1Ixp25_ASAP7_75t_L g466 ( 
.A1(n_447),
.A2(n_406),
.B(n_396),
.C(n_378),
.D(n_387),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_448),
.Y(n_467)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_467),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_381),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_469),
.A2(n_424),
.B1(n_450),
.B2(n_444),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_471),
.A2(n_453),
.B1(n_435),
.B2(n_428),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_380),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_472),
.B(n_475),
.Y(n_510)
);

CKINVDCx14_ASAP7_75t_R g474 ( 
.A(n_429),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_474),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_446),
.B(n_390),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_421),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_476),
.Y(n_532)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_448),
.Y(n_477)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_477),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_427),
.B(n_446),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_478),
.B(n_485),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_433),
.A2(n_392),
.B1(n_415),
.B2(n_422),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_479),
.Y(n_504)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_432),
.Y(n_480)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_480),
.Y(n_516)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_432),
.Y(n_481)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_481),
.Y(n_519)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_442),
.Y(n_483)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_483),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_427),
.B(n_400),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_442),
.Y(n_486)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_486),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_429),
.B(n_447),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_488),
.B(n_489),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_416),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_426),
.A2(n_407),
.B(n_399),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_490),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_461),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_491),
.B(n_437),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g539 ( 
.A(n_493),
.B(n_499),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_441),
.B(n_365),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_494),
.B(n_495),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_449),
.B(n_376),
.Y(n_495)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_462),
.Y(n_497)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_497),
.Y(n_506)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_462),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_498),
.B(n_500),
.Y(n_528)
);

MAJx2_ASAP7_75t_L g499 ( 
.A(n_438),
.B(n_402),
.C(n_403),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_452),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_439),
.A2(n_423),
.B(n_414),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_501),
.A2(n_458),
.B(n_443),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_456),
.B(n_413),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_459),
.C(n_430),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_505),
.A2(n_513),
.B(n_476),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_445),
.Y(n_508)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_508),
.B(n_514),
.C(n_527),
.Y(n_560)
);

AO22x1_ASAP7_75t_L g513 ( 
.A1(n_476),
.A2(n_477),
.B1(n_467),
.B2(n_451),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_470),
.B(n_445),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_515),
.B(n_493),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_517),
.A2(n_526),
.B1(n_492),
.B2(n_484),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_518),
.A2(n_529),
.B1(n_484),
.B2(n_440),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_496),
.B(n_425),
.C(n_459),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_522),
.B(n_537),
.C(n_538),
.Y(n_548)
);

CKINVDCx14_ASAP7_75t_R g524 ( 
.A(n_488),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_524),
.A2(n_501),
.B1(n_482),
.B2(n_487),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_479),
.A2(n_461),
.B1(n_453),
.B2(n_460),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_480),
.B(n_460),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_466),
.B(n_385),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_481),
.B(n_452),
.Y(n_530)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_530),
.Y(n_542)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_531),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_491),
.B(n_389),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_533),
.B(n_535),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_500),
.B(n_502),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_496),
.B(n_434),
.C(n_437),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_499),
.B(n_434),
.C(n_358),
.Y(n_538)
);

XOR2x1_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_490),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_540),
.B(n_541),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_528),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_543),
.A2(n_552),
.B1(n_558),
.B2(n_562),
.Y(n_572)
);

AO21x1_ASAP7_75t_L g588 ( 
.A1(n_545),
.A2(n_557),
.B(n_507),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_503),
.B(n_510),
.Y(n_546)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_546),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_522),
.B(n_482),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_547),
.B(n_550),
.Y(n_584)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_549),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_537),
.B(n_489),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_515),
.B(n_487),
.C(n_473),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_551),
.B(n_556),
.C(n_570),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_528),
.Y(n_552)
);

NOR2x1_ASAP7_75t_L g553 ( 
.A(n_536),
.B(n_469),
.Y(n_553)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_553),
.Y(n_590)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_516),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_554),
.A2(n_563),
.B1(n_564),
.B2(n_567),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_518),
.B(n_473),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_555),
.B(n_505),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_539),
.B(n_471),
.C(n_497),
.Y(n_556)
);

FAx1_ASAP7_75t_SL g557 ( 
.A(n_511),
.B(n_498),
.CI(n_486),
.CON(n_557),
.SN(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_520),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_539),
.B(n_483),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_559),
.B(n_569),
.Y(n_585)
);

AO22x1_ASAP7_75t_L g561 ( 
.A1(n_504),
.A2(n_492),
.B1(n_484),
.B2(n_440),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_561),
.A2(n_532),
.B(n_525),
.Y(n_587)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_516),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_SL g565 ( 
.A(n_509),
.B(n_504),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_SL g578 ( 
.A(n_565),
.B(n_513),
.Y(n_578)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_519),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_503),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_568),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_538),
.B(n_386),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_536),
.B(n_296),
.C(n_362),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_530),
.B(n_362),
.C(n_454),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_571),
.B(n_534),
.C(n_523),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_573),
.B(n_595),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_561),
.A2(n_517),
.B1(n_513),
.B2(n_532),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_576),
.A2(n_545),
.B1(n_540),
.B2(n_553),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_560),
.A2(n_525),
.B1(n_520),
.B2(n_510),
.Y(n_577)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_577),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_578),
.B(n_581),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_548),
.B(n_547),
.C(n_541),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_582),
.B(n_591),
.C(n_570),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_548),
.B(n_531),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_586),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_587),
.A2(n_557),
.B(n_565),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_588),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_562),
.A2(n_519),
.B1(n_507),
.B2(n_512),
.Y(n_589)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_589),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_556),
.B(n_512),
.C(n_509),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_542),
.A2(n_521),
.B1(n_484),
.B2(n_529),
.Y(n_592)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_592),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_544),
.A2(n_534),
.B1(n_523),
.B2(n_506),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_593),
.B(n_594),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_550),
.B(n_521),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_SL g595 ( 
.A(n_559),
.B(n_506),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_566),
.A2(n_454),
.B1(n_408),
.B2(n_411),
.Y(n_596)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_596),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_599),
.B(n_615),
.Y(n_634)
);

INVxp33_ASAP7_75t_L g600 ( 
.A(n_574),
.Y(n_600)
);

INVxp67_ASAP7_75t_SL g623 ( 
.A(n_600),
.Y(n_623)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_583),
.B(n_555),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_602),
.B(n_609),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_603),
.A2(n_619),
.B1(n_579),
.B2(n_590),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_605),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_582),
.B(n_569),
.C(n_551),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_606),
.B(n_614),
.Y(n_637)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_583),
.B(n_573),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_586),
.B(n_571),
.C(n_557),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_584),
.B(n_454),
.C(n_410),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_572),
.A2(n_411),
.B1(n_368),
.B2(n_319),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_616),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g617 ( 
.A(n_575),
.B(n_337),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_617),
.B(n_574),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_SL g618 ( 
.A1(n_587),
.A2(n_347),
.B(n_255),
.Y(n_618)
);

MAJx2_ASAP7_75t_L g631 ( 
.A(n_618),
.B(n_588),
.C(n_578),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g619 ( 
.A1(n_576),
.A2(n_336),
.B1(n_347),
.B2(n_344),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_606),
.B(n_584),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_622),
.B(n_624),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_599),
.B(n_580),
.C(n_591),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_608),
.Y(n_625)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_625),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_626),
.B(n_631),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_610),
.B(n_580),
.C(n_585),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_628),
.B(n_629),
.Y(n_644)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_600),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_601),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_630),
.B(n_632),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_604),
.B(n_594),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_607),
.B(n_609),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_633),
.B(n_607),
.Y(n_640)
);

XOR2xp5_ASAP7_75t_L g635 ( 
.A(n_602),
.B(n_585),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_635),
.B(n_598),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_636),
.B(n_615),
.Y(n_639)
);

OAI21xp33_ASAP7_75t_L g638 ( 
.A1(n_627),
.A2(n_605),
.B(n_603),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_638),
.B(n_640),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_639),
.A2(n_641),
.B1(n_646),
.B2(n_623),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_637),
.A2(n_604),
.B(n_613),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_624),
.B(n_611),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_642),
.B(n_652),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_634),
.B(n_614),
.C(n_612),
.Y(n_645)
);

NOR2xp67_ASAP7_75t_SL g656 ( 
.A(n_645),
.B(n_649),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_626),
.A2(n_597),
.B1(n_612),
.B2(n_616),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_628),
.B(n_581),
.C(n_598),
.Y(n_649)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_651),
.B(n_344),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_620),
.B(n_595),
.C(n_618),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_643),
.B(n_621),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_653),
.B(n_655),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_647),
.B(n_623),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_657),
.B(n_660),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_650),
.A2(n_619),
.B1(n_631),
.B2(n_635),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_659),
.B(n_661),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_644),
.Y(n_660)
);

XOR2xp5_ASAP7_75t_L g662 ( 
.A(n_645),
.B(n_256),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g666 ( 
.A(n_662),
.B(n_663),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_SL g663 ( 
.A1(n_638),
.A2(n_649),
.B(n_648),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_656),
.B(n_648),
.C(n_651),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_664),
.B(n_668),
.Y(n_672)
);

AOI322xp5_ASAP7_75t_L g667 ( 
.A1(n_654),
.A2(n_652),
.A3(n_287),
.B1(n_259),
.B2(n_254),
.C1(n_243),
.C2(n_247),
.Y(n_667)
);

AOI21xp33_ASAP7_75t_L g671 ( 
.A1(n_667),
.A2(n_659),
.B(n_662),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g668 ( 
.A(n_658),
.B(n_269),
.Y(n_668)
);

AOI322xp5_ASAP7_75t_L g675 ( 
.A1(n_671),
.A2(n_673),
.A3(n_674),
.B1(n_669),
.B2(n_667),
.C1(n_666),
.C2(n_238),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_SL g673 ( 
.A1(n_670),
.A2(n_661),
.B(n_305),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_665),
.B(n_257),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_675),
.B(n_676),
.Y(n_677)
);

AOI322xp5_ASAP7_75t_L g676 ( 
.A1(n_672),
.A2(n_669),
.A3(n_177),
.B1(n_348),
.B2(n_273),
.C1(n_236),
.C2(n_261),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g678 ( 
.A(n_675),
.B(n_348),
.C(n_269),
.Y(n_678)
);

XNOR2x2_ASAP7_75t_SL g679 ( 
.A(n_678),
.B(n_246),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_677),
.Y(n_680)
);

OAI221xp5_ASAP7_75t_SL g681 ( 
.A1(n_680),
.A2(n_241),
.B1(n_224),
.B2(n_288),
.C(n_17),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_681),
.A2(n_311),
.B(n_233),
.Y(n_682)
);


endmodule