module fake_netlist_1_10722_n_25 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_25);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
NAND2xp5_ASAP7_75t_L g8 ( .A(n_4), .B(n_1), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_5), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_6), .B(n_3), .Y(n_10) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_7), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_12), .B(n_0), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
AO31x2_ASAP7_75t_L g17 ( .A1(n_15), .A2(n_9), .A3(n_8), .B(n_10), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_18), .B(n_13), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_19), .B(n_17), .Y(n_20) );
AOI21xp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_17), .B(n_1), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
INVxp67_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
BUFx2_ASAP7_75t_SL g25 ( .A(n_24), .Y(n_25) );
endmodule