module fake_jpeg_1785_n_295 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_57),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_43),
.B(n_50),
.Y(n_90)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_44),
.Y(n_83)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_25),
.B(n_1),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_32),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_62),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_28),
.B(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_1),
.Y(n_99)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

BUFx12f_ASAP7_75t_SL g60 ( 
.A(n_29),
.Y(n_60)
);

HAxp5_ASAP7_75t_SL g89 ( 
.A(n_60),
.B(n_64),
.CON(n_89),
.SN(n_89)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

BUFx12f_ASAP7_75t_SL g64 ( 
.A(n_29),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_19),
.Y(n_65)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_41),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_17),
.B1(n_40),
.B2(n_38),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_41),
.B1(n_21),
.B2(n_39),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_68),
.A2(n_93),
.B1(n_105),
.B2(n_107),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_40),
.B(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_74),
.B(n_79),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_36),
.B1(n_39),
.B2(n_37),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_68),
.B1(n_84),
.B2(n_75),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_77),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_88),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_82),
.B(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_36),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_101),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_37),
.B1(n_34),
.B2(n_30),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_SL g94 ( 
.A1(n_42),
.A2(n_47),
.B(n_49),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_47),
.Y(n_114)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_2),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_55),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_66),
.A2(n_52),
.B1(n_56),
.B2(n_63),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_34),
.B1(n_30),
.B2(n_27),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_59),
.A2(n_27),
.B1(n_46),
.B2(n_61),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_24),
.B1(n_5),
.B2(n_6),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_110),
.B(n_144),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_114),
.B(n_129),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_120),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_46),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_82),
.A2(n_24),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_123),
.A2(n_141),
.B1(n_120),
.B2(n_111),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_3),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_3),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_91),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_3),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_134),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_72),
.B(n_81),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_73),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_86),
.B1(n_98),
.B2(n_97),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_7),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_85),
.C(n_71),
.Y(n_157)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_86),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_83),
.B(n_16),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_83),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_103),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_145),
.A2(n_159),
.B1(n_163),
.B2(n_169),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_155),
.Y(n_178)
);

NAND2x1_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_89),
.Y(n_150)
);

XNOR2x1_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_157),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_116),
.A2(n_100),
.B(n_81),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_152),
.A2(n_171),
.B(n_166),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_153),
.A2(n_112),
.B1(n_121),
.B2(n_156),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_69),
.B(n_106),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_118),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_100),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_164),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_95),
.B1(n_72),
.B2(n_102),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_120),
.B(n_85),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_87),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_109),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_87),
.B1(n_12),
.B2(n_14),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_9),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_14),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_166),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_15),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_15),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_158),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_111),
.A2(n_16),
.B1(n_115),
.B2(n_123),
.Y(n_169)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_115),
.A2(n_16),
.B(n_138),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_115),
.A2(n_132),
.B1(n_143),
.B2(n_135),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_131),
.B1(n_136),
.B2(n_133),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_143),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_182),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_150),
.B(n_140),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_198),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_170),
.B(n_139),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_184),
.B(n_193),
.Y(n_211)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_190),
.B1(n_202),
.B2(n_205),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_136),
.B1(n_112),
.B2(n_121),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_146),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_207),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_197),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_150),
.B(n_168),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_149),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_157),
.C(n_177),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_169),
.B1(n_147),
.B2(n_149),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_146),
.B(n_164),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_203),
.B(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_147),
.A2(n_163),
.B1(n_165),
.B2(n_171),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_206),
.A2(n_172),
.B(n_176),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_168),
.B(n_174),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_230),
.B(n_216),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_153),
.B1(n_161),
.B2(n_176),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_212),
.B(n_209),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_221),
.C(n_226),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_191),
.A2(n_145),
.B1(n_173),
.B2(n_177),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_217),
.A2(n_187),
.B1(n_204),
.B2(n_195),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_220),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_172),
.C(n_198),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_199),
.B1(n_205),
.B2(n_190),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_222),
.A2(n_225),
.B1(n_183),
.B2(n_215),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_179),
.A2(n_185),
.B1(n_200),
.B2(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_185),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_227),
.B(n_228),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_201),
.B(n_196),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_231),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_189),
.B(n_188),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_186),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_192),
.B1(n_187),
.B2(n_195),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_233),
.B1(n_239),
.B2(n_249),
.Y(n_255)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_211),
.B(n_208),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_242),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_221),
.C(n_226),
.Y(n_251)
);

NAND2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_238),
.A2(n_240),
.B(n_244),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_230),
.B1(n_212),
.B2(n_225),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_231),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_211),
.B(n_208),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_229),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_248),
.Y(n_261)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_223),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_219),
.B1(n_213),
.B2(n_224),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_259),
.C(n_234),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_236),
.B(n_224),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_251),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_233),
.Y(n_257)
);

INVx11_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_216),
.C(n_214),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_244),
.A2(n_210),
.B(n_214),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_260),
.A2(n_238),
.B(n_237),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_265),
.C(n_271),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g264 ( 
.A(n_253),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_264),
.B(n_250),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_256),
.B(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_259),
.B(n_245),
.CI(n_243),
.CON(n_267),
.SN(n_267)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_261),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_270),
.B(n_262),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_239),
.B(n_232),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_243),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_252),
.A2(n_241),
.B1(n_245),
.B2(n_247),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_270),
.A2(n_252),
.B1(n_256),
.B2(n_258),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_280),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_271),
.B(n_266),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_269),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_255),
.B1(n_262),
.B2(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_279),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_265),
.C(n_263),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_277),
.C(n_273),
.Y(n_289)
);

OAI211xp5_ASAP7_75t_L g287 ( 
.A1(n_283),
.A2(n_284),
.B(n_276),
.C(n_280),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_272),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_287),
.B(n_289),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_276),
.B(n_277),
.C(n_267),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_285),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_291),
.A2(n_288),
.A3(n_267),
.B1(n_285),
.B2(n_268),
.C1(n_281),
.C2(n_217),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_292),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_268),
.Y(n_295)
);


endmodule