module fake_jpeg_10626_n_84 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_84);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_84;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_SL g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_11),
.B(n_23),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_23),
.Y(n_33)
);

CKINVDCx12_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_11),
.B(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_40),
.Y(n_42)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_18),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_25),
.B1(n_16),
.B2(n_24),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_47),
.B1(n_52),
.B2(n_17),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_48),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_23),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_49),
.B(n_51),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_25),
.B1(n_13),
.B2(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2x1_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_26),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_32),
.A2(n_16),
.B1(n_15),
.B2(n_17),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_15),
.B1(n_17),
.B2(n_21),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_21),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g61 ( 
.A(n_53),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_12),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_50),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_64),
.C(n_66),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_47),
.C(n_42),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_47),
.Y(n_65)
);

AOI322xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_54),
.A3(n_60),
.B1(n_57),
.B2(n_18),
.C1(n_20),
.C2(n_12),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_48),
.C(n_29),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_73),
.B1(n_74),
.B2(n_20),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_66),
.B(n_67),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_72),
.B(n_71),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_19),
.Y(n_79)
);

FAx1_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_70),
.CI(n_73),
.CON(n_78),
.SN(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_79),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_78),
.A2(n_77),
.B(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

AOI322xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_81),
.A3(n_3),
.B1(n_5),
.B2(n_8),
.C1(n_10),
.C2(n_0),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);


endmodule