module fake_jpeg_8215_n_113 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_113);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_113;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_27),
.B(n_23),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_13),
.Y(n_39)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_32),
.Y(n_38)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_15),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_43),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_13),
.B1(n_25),
.B2(n_17),
.Y(n_40)
);

NOR2x1p5_ASAP7_75t_SL g63 ( 
.A(n_40),
.B(n_26),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_19),
.B1(n_25),
.B2(n_17),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_50),
.B1(n_35),
.B2(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_58),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_54),
.Y(n_71)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVxp33_ASAP7_75t_SL g77 ( 
.A(n_55),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_30),
.C(n_27),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_22),
.CI(n_14),
.CON(n_70),
.SN(n_70)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_33),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_40),
.Y(n_68)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_61),
.B(n_60),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_69),
.B(n_56),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_53),
.B1(n_48),
.B2(n_59),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_48),
.B(n_22),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_38),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_14),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_12),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_76),
.B(n_72),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_79),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_51),
.C(n_57),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_83),
.C(n_70),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_57),
.B(n_22),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_86),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_67),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_90),
.C(n_83),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_96),
.C(n_99),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_81),
.C(n_70),
.Y(n_96)
);

BUFx4f_ASAP7_75t_SL g97 ( 
.A(n_93),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_91),
.B(n_92),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_98),
.A2(n_12),
.B(n_47),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_92),
.C(n_67),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_101),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_47),
.B(n_46),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_106),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_2),
.C(n_7),
.Y(n_109)
);

AOI31xp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_8),
.A3(n_9),
.B(n_11),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_105),
.B1(n_8),
.B2(n_59),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_108),
.B(n_55),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_65),
.Y(n_113)
);


endmodule