module fake_jpeg_7382_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

OR2x2_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_23),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_25),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_16),
.A2(n_0),
.B1(n_2),
.B2(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_17),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_45),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_22),
.B1(n_16),
.B2(n_27),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_22),
.B1(n_30),
.B2(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_18),
.B1(n_10),
.B2(n_17),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_12),
.B1(n_19),
.B2(n_14),
.Y(n_49)
);

OA21x2_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_32),
.B(n_31),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_40),
.B1(n_47),
.B2(n_41),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_36),
.C(n_26),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_15),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_15),
.B(n_19),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_49),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_54),
.C(n_57),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_55),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_64),
.A2(n_59),
.B(n_65),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_50),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_69),
.C(n_70),
.Y(n_72)
);

AOI322xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_59),
.A3(n_53),
.B1(n_50),
.B2(n_24),
.C1(n_11),
.C2(n_12),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_41),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_15),
.C(n_34),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_72),
.A2(n_64),
.B(n_11),
.C(n_0),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_5),
.A3(n_6),
.B1(n_8),
.B2(n_34),
.C1(n_74),
.C2(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);


endmodule