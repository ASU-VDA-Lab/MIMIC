module real_jpeg_16693_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_249;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_286;
wire n_288;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_293;
wire n_164;
wire n_275;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_185;
wire n_297;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_295;
wire n_128;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_0),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_0),
.A2(n_58),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_1),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g20 ( 
.A1(n_2),
.A2(n_21),
.A3(n_26),
.B1(n_30),
.B2(n_35),
.Y(n_20)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_2),
.A2(n_31),
.B1(n_140),
.B2(n_145),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_2),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_2),
.A2(n_48),
.B1(n_292),
.B2(n_297),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_3),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_3),
.Y(n_247)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_3),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_4),
.A2(n_108),
.B1(n_109),
.B2(n_113),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_4),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_4),
.A2(n_72),
.B1(n_108),
.B2(n_218),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_5),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_5),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_6),
.Y(n_184)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_6),
.Y(n_227)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_7),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_7),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_7),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_7),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_7),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_8),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_8),
.A2(n_85),
.B1(n_162),
.B2(n_167),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_8),
.A2(n_85),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_9),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_9),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_11),
.A2(n_67),
.B1(n_71),
.B2(n_72),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_12),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_13),
.A2(n_151),
.B1(n_154),
.B2(n_156),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_13),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_13),
.A2(n_156),
.B1(n_211),
.B2(n_214),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_13),
.A2(n_156),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_205),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_204),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_157),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_18),
.B(n_157),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_78),
.C(n_119),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_19),
.B(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_46),
.B1(n_76),
.B2(n_77),
.Y(n_19)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_20),
.B(n_77),
.Y(n_194)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_24),
.Y(n_153)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_25),
.Y(n_177)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_29),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_31),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_31),
.B(n_249),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_SL g264 ( 
.A1(n_31),
.A2(n_248),
.B(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_31),
.B(n_223),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_31),
.B(n_118),
.Y(n_300)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_33),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_36),
.A2(n_123),
.B(n_129),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_42),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_40),
.Y(n_125)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_44),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_45),
.Y(n_128)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_45),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_45),
.Y(n_166)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_55),
.B1(n_62),
.B2(n_66),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_47),
.A2(n_66),
.B1(n_182),
.B2(n_185),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_47),
.A2(n_273),
.B1(n_281),
.B2(n_283),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_48),
.A2(n_217),
.B1(n_223),
.B2(n_228),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_48),
.A2(n_64),
.B1(n_274),
.B2(n_292),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_91),
.B1(n_92),
.B2(n_96),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_54),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_55),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_57),
.Y(n_191)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_57),
.Y(n_222)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_57),
.Y(n_294)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_61),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_74),
.Y(n_296)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_75),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_78),
.A2(n_119),
.B1(n_120),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_78),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_89),
.B1(n_107),
.B2(n_117),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_79),
.A2(n_89),
.B1(n_117),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_89),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_89),
.A2(n_117),
.B1(n_210),
.B2(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_98),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_94),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_94),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_99),
.B1(n_101),
.B2(n_104),
.Y(n_98)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_105),
.Y(n_201)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_107),
.Y(n_197)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_118),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_195)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_139),
.B1(n_149),
.B2(n_150),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_121),
.A2(n_149),
.B1(n_150),
.B2(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_132),
.B1(n_134),
.B2(n_136),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_133),
.Y(n_267)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_149),
.Y(n_231)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_192),
.B2(n_193),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_171),
.Y(n_159)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AO22x2_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_180),
.B2(n_181),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_182),
.Y(n_297)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_202),
.B2(n_203),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_235),
.B(n_304),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_232),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_207),
.B(n_232),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_216),
.C(n_229),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_208),
.A2(n_209),
.B1(n_229),
.B2(n_230),
.Y(n_269)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_269),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_217),
.Y(n_283)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_218),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_224),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI21x1_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_270),
.B(n_303),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_268),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_237),
.B(n_268),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_262),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_238),
.A2(n_262),
.B1(n_263),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

OAI32xp33_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.A3(n_245),
.B1(n_248),
.B2(n_253),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_286),
.B(n_302),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_284),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_284),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_298),
.B(n_301),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_300),
.Y(n_301)
);


endmodule