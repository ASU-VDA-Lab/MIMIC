module real_jpeg_11811_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_249;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_286;
wire n_292;
wire n_221;
wire n_215;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_299;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_200;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_195;
wire n_110;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_295;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_3),
.A2(n_37),
.B1(n_41),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_3),
.A2(n_44),
.B1(n_60),
.B2(n_61),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_44),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_4),
.A2(n_55),
.B1(n_57),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_4),
.A2(n_60),
.B1(n_61),
.B2(n_104),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_4),
.A2(n_37),
.B1(n_41),
.B2(n_104),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_104),
.Y(n_252)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_6),
.A2(n_37),
.B1(n_41),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_6),
.A2(n_47),
.B1(n_55),
.B2(n_57),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_47),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_6),
.A2(n_47),
.B1(n_60),
.B2(n_61),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_7),
.A2(n_55),
.B1(n_57),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_7),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_7),
.A2(n_60),
.B1(n_61),
.B2(n_168),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_7),
.A2(n_37),
.B1(n_41),
.B2(n_168),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_168),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_10),
.A2(n_55),
.B1(n_57),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_10),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_145),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_10),
.A2(n_37),
.B1(n_41),
.B2(n_145),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_145),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_11),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_11),
.B(n_106),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_11),
.B(n_27),
.C(n_40),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_11),
.A2(n_37),
.B1(n_41),
.B2(n_160),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_11),
.A2(n_24),
.B1(n_30),
.B2(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_11),
.B(n_82),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_12),
.A2(n_33),
.B1(n_55),
.B2(n_57),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_12),
.A2(n_33),
.B1(n_37),
.B2(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_12),
.A2(n_33),
.B1(n_60),
.B2(n_61),
.Y(n_148)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_14),
.A2(n_60),
.B1(n_61),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_14),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_14),
.A2(n_37),
.B1(n_41),
.B2(n_76),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_14),
.A2(n_55),
.B1(n_57),
.B2(n_76),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_76),
.Y(n_157)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_107),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_19),
.B(n_107),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_66),
.C(n_85),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_20),
.A2(n_21),
.B1(n_66),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_48),
.Y(n_21)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_22),
.A2(n_23),
.B(n_50),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_23),
.A2(n_49),
.B1(n_50),
.B2(n_65),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_23),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_23),
.A2(n_34),
.B1(n_65),
.B2(n_177),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_31),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_24),
.A2(n_136),
.B(n_138),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_24),
.A2(n_30),
.B1(n_250),
.B2(n_258),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_24),
.A2(n_94),
.B(n_252),
.Y(n_272)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_25),
.B(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_25),
.A2(n_29),
.B1(n_137),
.B2(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_25),
.A2(n_32),
.B(n_139),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_25),
.A2(n_29),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_26),
.A2(n_27),
.B1(n_38),
.B2(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_26),
.B(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_29),
.B(n_32),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_30),
.B(n_93),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_30),
.A2(n_91),
.B(n_157),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_30),
.B(n_160),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_34),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_43),
.B(n_45),
.Y(n_34)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_35),
.A2(n_43),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_35),
.A2(n_70),
.B(n_97),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_35),
.A2(n_45),
.B(n_70),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_35),
.A2(n_68),
.B(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_35),
.A2(n_97),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_35),
.A2(n_97),
.B1(n_224),
.B2(n_247),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_36)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

OA22x2_ASAP7_75t_SL g81 ( 
.A1(n_37),
.A2(n_41),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_37),
.A2(n_79),
.B(n_219),
.C(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_37),
.B(n_243),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_SL g40 ( 
.A(n_38),
.Y(n_40)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_41),
.B(n_61),
.C(n_80),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_42),
.A2(n_72),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_72),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_62),
.B(n_63),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_51),
.A2(n_106),
.B1(n_159),
.B2(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_52),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_64),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_52),
.A2(n_59),
.B1(n_103),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_52),
.A2(n_59),
.B1(n_144),
.B2(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_54),
.A2(n_61),
.B(n_159),
.C(n_161),
.Y(n_158)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_55),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

HAxp5_ASAP7_75t_SL g159 ( 
.A(n_57),
.B(n_160),
.CON(n_159),
.SN(n_159)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_57),
.B(n_58),
.C(n_60),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_61),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HAxp5_ASAP7_75t_SL g219 ( 
.A(n_61),
.B(n_160),
.CON(n_219),
.SN(n_219)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_66),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_73),
.B(n_84),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_73),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_71),
.A2(n_96),
.B(n_97),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_81),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_77),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_77),
.A2(n_121),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_77),
.A2(n_82),
.B1(n_196),
.B2(n_219),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_101),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_81),
.A2(n_118),
.B1(n_163),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_81),
.A2(n_118),
.B1(n_187),
.B2(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_82),
.B(n_148),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_110),
.B1(n_111),
.B2(n_126),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_85),
.A2(n_86),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_98),
.C(n_102),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_87),
.A2(n_88),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_95),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_97),
.B(n_160),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_98),
.B(n_102),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_124),
.B2(n_125),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_122),
.B2(n_123),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B(n_120),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_118),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_122),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_293),
.B(n_299),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_179),
.B(n_292),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_169),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_132),
.B(n_169),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_149),
.C(n_151),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_133),
.B(n_149),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_141),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_142),
.C(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_140),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_135),
.B(n_140),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_151),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_162),
.C(n_165),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_152),
.A2(n_153),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_154),
.A2(n_155),
.B1(n_158),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_165),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_178),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_171),
.B(n_176),
.C(n_178),
.Y(n_298)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_207),
.B(n_287),
.C(n_291),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_200),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_200),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_190),
.C(n_193),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_182),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_185),
.C(n_189),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_193),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.C(n_199),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_194),
.B(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_201),
.B(n_205),
.C(n_206),
.Y(n_288)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_281),
.B(n_286),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_236),
.B(n_280),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_226),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_212),
.B(n_226),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_221),
.C(n_222),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_213),
.A2(n_214),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_215),
.B(n_218),
.Y(n_231)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_221),
.B(n_222),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_225),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_227),
.B(n_232),
.C(n_234),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_274),
.B(n_279),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_264),
.B(n_273),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_253),
.B(n_263),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_248),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_248),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_259),
.B(n_262),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_261),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_266),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_272),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_271),
.C(n_272),
.Y(n_278)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_278),
.Y(n_279)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_285),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_289),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_298),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_298),
.Y(n_299)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);


endmodule