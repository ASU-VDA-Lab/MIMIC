module fake_jpeg_21991_n_166 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_166);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_11),
.B(n_1),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_24),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_20),
.Y(n_54)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_28),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_13),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_17),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_35),
.C(n_11),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_32),
.A2(n_25),
.B1(n_17),
.B2(n_22),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_68),
.B1(n_71),
.B2(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_33),
.A2(n_27),
.B1(n_17),
.B2(n_23),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_43),
.B(n_41),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_33),
.A2(n_27),
.B1(n_28),
.B2(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_2),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_70),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_34),
.A2(n_2),
.B1(n_5),
.B2(n_8),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_86),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_82),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_10),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_50),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_45),
.C(n_12),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_12),
.B1(n_13),
.B2(n_55),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_46),
.B1(n_52),
.B2(n_51),
.Y(n_85)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_53),
.C(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_94),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_50),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_112),
.Y(n_117)
);

CKINVDCx12_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_65),
.B1(n_77),
.B2(n_87),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_75),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_107),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_73),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_78),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_101),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_128),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_77),
.C(n_76),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_120),
.C(n_122),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_82),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_105),
.B(n_112),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_81),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_88),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_98),
.B(n_95),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_131),
.B(n_139),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_139),
.C(n_103),
.Y(n_147)
);

OAI21x1_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_96),
.B(n_110),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_106),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_110),
.B1(n_96),
.B2(n_105),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_106),
.C(n_96),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_142),
.Y(n_149)
);

AO221x1_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_121),
.B1(n_127),
.B2(n_126),
.C(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_115),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_148),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_145),
.B1(n_137),
.B2(n_135),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_145),
.C(n_130),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_143),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_135),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_147),
.B(n_148),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_156),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_158),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_149),
.A2(n_133),
.B(n_93),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_91),
.Y(n_161)
);

AO21x2_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_153),
.B(n_162),
.Y(n_164)
);

OAI221xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_156),
.B1(n_152),
.B2(n_153),
.C(n_91),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_163),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_164),
.Y(n_166)
);


endmodule