module real_jpeg_17438_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_0),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_536),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_1),
.B(n_537),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_2),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_2),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_3),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_3),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_3),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_4),
.A2(n_119),
.B1(n_255),
.B2(n_258),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_4),
.A2(n_119),
.B1(n_379),
.B2(n_381),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_4),
.A2(n_119),
.B1(n_345),
.B2(n_452),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_5),
.A2(n_272),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_5),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_5),
.A2(n_326),
.B1(n_425),
.B2(n_437),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_5),
.A2(n_326),
.B1(n_513),
.B2(n_515),
.Y(n_512)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_6),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_7),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_7),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_8),
.A2(n_201),
.B1(n_204),
.B2(n_207),
.Y(n_200)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_8),
.A2(n_207),
.B1(n_421),
.B2(n_424),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g479 ( 
.A1(n_8),
.A2(n_207),
.B1(n_480),
.B2(n_482),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_9),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_9),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_9),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g388 ( 
.A(n_9),
.Y(n_388)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_9),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_10),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_10),
.A2(n_68),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_10),
.A2(n_46),
.B1(n_68),
.B2(n_380),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_10),
.A2(n_68),
.B1(n_489),
.B2(n_491),
.Y(n_488)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_11),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_11),
.Y(n_348)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_11),
.Y(n_355)
);

OAI32xp33_ASAP7_75t_L g29 ( 
.A1(n_12),
.A2(n_30),
.A3(n_36),
.B1(n_39),
.B2(n_44),
.Y(n_29)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_12),
.A2(n_43),
.B1(n_148),
.B2(n_152),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_12),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_12),
.B(n_122),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_12),
.B(n_287),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_12),
.B(n_242),
.Y(n_304)
);

OAI32xp33_ASAP7_75t_L g327 ( 
.A1(n_12),
.A2(n_328),
.A3(n_331),
.B1(n_336),
.B2(n_343),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_12),
.A2(n_43),
.B1(n_364),
.B2(n_366),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_13),
.A2(n_159),
.B1(n_164),
.B2(n_166),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_13),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_13),
.A2(n_166),
.B1(n_244),
.B2(n_250),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_13),
.A2(n_166),
.B1(n_289),
.B2(n_293),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_13),
.A2(n_166),
.B1(n_371),
.B2(n_373),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_14),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_15),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_15),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_15),
.A2(n_77),
.B1(n_387),
.B2(n_389),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_15),
.A2(n_77),
.B1(n_446),
.B2(n_448),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_15),
.A2(n_77),
.B1(n_526),
.B2(n_529),
.Y(n_525)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_17),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_17),
.Y(n_357)
);

BUFx8_ASAP7_75t_L g359 ( 
.A(n_17),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g528 ( 
.A(n_17),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_502),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_463),
.B(n_500),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_396),
.B(n_459),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_314),
.B(n_395),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_219),
.B(n_313),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_168),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_27),
.B(n_168),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_83),
.C(n_120),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_28),
.B(n_311),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_53),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_29),
.B(n_53),
.Y(n_170)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_34),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_34),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_35),
.Y(n_139)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_35),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_35),
.Y(n_189)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_37),
.Y(n_179)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_43),
.B(n_96),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_SL g239 ( 
.A1(n_43),
.A2(n_230),
.B(n_240),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_43),
.A2(n_55),
.B1(n_286),
.B2(n_288),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_43),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_48),
.Y(n_163)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_48),
.Y(n_330)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_63),
.B(n_70),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_54),
.A2(n_270),
.B1(n_279),
.B2(n_280),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_54),
.A2(n_200),
.B1(n_322),
.B2(n_324),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_54),
.A2(n_70),
.B(n_324),
.Y(n_417)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_55),
.B(n_71),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_55),
.A2(n_254),
.B(n_260),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_55),
.A2(n_271),
.B1(n_288),
.B2(n_301),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_55),
.A2(n_64),
.B(n_470),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_58),
.Y(n_206)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_61),
.Y(n_303)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_64),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_65),
.Y(n_325)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_66),
.Y(n_259)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_66),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_67),
.Y(n_276)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_69),
.Y(n_226)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_76),
.Y(n_203)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_76),
.Y(n_257)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_76),
.Y(n_292)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_82),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_83),
.B(n_120),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_97),
.B1(n_104),
.B2(n_115),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_84),
.A2(n_174),
.B(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_84),
.A2(n_97),
.B1(n_435),
.B2(n_436),
.Y(n_434)
);

OA21x2_ASAP7_75t_L g473 ( 
.A1(n_84),
.A2(n_385),
.B(n_436),
.Y(n_473)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_85),
.A2(n_172),
.B(n_173),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_85),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_85),
.A2(n_105),
.B1(n_242),
.B2(n_243),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_85),
.B(n_386),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_97),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_90),
.B1(n_92),
.B2(n_96),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_88),
.Y(n_225)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVxp67_ASAP7_75t_SL g251 ( 
.A(n_89),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_91),
.Y(n_229)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_97),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_97),
.Y(n_242)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_108),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_108),
.Y(n_438)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_109),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_110),
.A2(n_111),
.B1(n_213),
.B2(n_217),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_110),
.A2(n_111),
.B1(n_272),
.B2(n_277),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_110),
.A2(n_111),
.B1(n_374),
.B2(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_116),
.Y(n_241)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_147),
.B1(n_158),
.B2(n_167),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_121),
.A2(n_167),
.B1(n_212),
.B2(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_121),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_121),
.A2(n_413),
.B(n_444),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_121),
.A2(n_167),
.B1(n_478),
.B2(n_479),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_132),
.Y(n_121)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_122),
.B(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_122),
.A2(n_410),
.B1(n_511),
.B2(n_512),
.Y(n_510)
);

AO22x2_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_137),
.B1(n_140),
.B2(n_143),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_139),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_139),
.Y(n_449)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_139),
.Y(n_514)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_146),
.Y(n_342)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_146),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_146),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_149),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AO22x2_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_209)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_163),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_167),
.B(n_413),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_180),
.B1(n_181),
.B2(n_218),
.Y(n_168)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_170),
.B(n_171),
.C(n_180),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_173),
.B(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_209),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_192),
.B2(n_193),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_183),
.B(n_193),
.C(n_209),
.Y(n_318)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_185),
.B(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_185),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_185),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_185),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_185),
.B(n_525),
.Y(n_524)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

INVx3_ASAP7_75t_SL g362 ( 
.A(n_188),
.Y(n_362)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_189),
.Y(n_447)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_200),
.B(n_208),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_SL g263 ( 
.A(n_197),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_197),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_199),
.Y(n_323)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_203),
.Y(n_293)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_208),
.B(n_261),
.Y(n_433)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_308),
.B(n_312),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_267),
.B(n_307),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_252),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_222),
.B(n_252),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_237),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_223),
.A2(n_237),
.B1(n_238),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_223),
.Y(n_282)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_226),
.A3(n_227),
.B1(n_230),
.B2(n_231),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_242),
.B(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_242),
.B(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_264),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_253),
.B(n_265),
.C(n_266),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

OAI21x1_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_283),
.B(n_306),
.Y(n_267)
);

NOR2x1_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_281),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_281),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_299),
.B(n_305),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_294),
.Y(n_284)
);

INVx6_ASAP7_75t_L g471 ( 
.A(n_286),
.Y(n_471)
);

BUFx12f_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_304),
.Y(n_305)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_309),
.B(n_310),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_394),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_315),
.B(n_394),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_349),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_318),
.B(n_319),
.C(n_349),
.Y(n_456)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_327),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_321),
.B(n_327),
.Y(n_414)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_334),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_334),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_342),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_347),
.Y(n_343)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_376),
.Y(n_349)
);

MAJx2_ASAP7_75t_L g415 ( 
.A(n_350),
.B(n_377),
.C(n_384),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_363),
.B1(n_370),
.B2(n_375),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_351),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_351),
.A2(n_375),
.B1(n_406),
.B2(n_451),
.Y(n_450)
);

OAI21x1_ASAP7_75t_SL g486 ( 
.A1(n_351),
.A2(n_451),
.B(n_487),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_351),
.A2(n_523),
.B(n_524),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_356),
.B1(n_358),
.B2(n_360),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx12f_ASAP7_75t_L g365 ( 
.A(n_357),
.Y(n_365)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_359),
.Y(n_374)
);

BUFx12f_ASAP7_75t_L g530 ( 
.A(n_359),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_365),
.Y(n_408)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_368),
.Y(n_372)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_369),
.Y(n_453)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_369),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_384),
.Y(n_376)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_378),
.Y(n_411)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_455),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_429),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_399),
.B(n_429),
.C(n_462),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_415),
.C(n_416),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_400),
.B(n_458),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_414),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_409),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_402),
.B(n_409),
.C(n_414),
.Y(n_430)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_411),
.B(n_412),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_415),
.B(n_416),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_418),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_428),
.Y(n_418)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_420),
.Y(n_435)
);

BUFx2_ASAP7_75t_SL g421 ( 
.A(n_422),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVxp33_ASAP7_75t_L g518 ( 
.A(n_428),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_439),
.C(n_454),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_439),
.B1(n_440),
.B2(n_454),
.Y(n_431)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_432),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_433),
.B(n_434),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_440),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_441),
.B(n_497),
.C(n_498),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_450),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_443),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_445),
.Y(n_478)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_450),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_457),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_460),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_465),
.B(n_466),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_467),
.A2(n_495),
.B1(n_496),
.B2(n_499),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_467),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_475),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_475),
.C(n_495),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_469),
.A2(n_472),
.B1(n_473),
.B2(n_474),
.Y(n_468)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_469),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_469),
.A2(n_474),
.B1(n_522),
.B2(n_531),
.Y(n_521)
);

NOR2x1_ASAP7_75t_L g532 ( 
.A(n_469),
.B(n_473),
.Y(n_532)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

XNOR2x1_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_494),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_486),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_477),
.Y(n_507)
);

INVxp33_ASAP7_75t_SL g511 ( 
.A(n_479),
.Y(n_511)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_486),
.B(n_494),
.C(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_488),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVxp33_ASAP7_75t_SL g500 ( 
.A(n_501),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_535),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_505),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_504),
.B(n_505),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_508),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_509),
.A2(n_520),
.B1(n_533),
.B2(n_534),
.Y(n_508)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_509),
.Y(n_533)
);

OAI21xp33_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_517),
.B(n_519),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_510),
.B(n_517),
.Y(n_519)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_520),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_532),
.Y(n_520)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_522),
.Y(n_531)
);

INVx6_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);


endmodule