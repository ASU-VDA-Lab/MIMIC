module fake_jpeg_8203_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_18),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_46),
.Y(n_73)
);

BUFx3_ASAP7_75t_SL g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_44),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_20),
.B(n_7),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_19),
.B(n_0),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_52),
.Y(n_84)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_61),
.Y(n_95)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_74),
.B1(n_37),
.B2(n_39),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_34),
.C(n_17),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_72),
.C(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_34),
.C(n_17),
.Y(n_72)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_17),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_78),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_35),
.B1(n_30),
.B2(n_16),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_79),
.A2(n_30),
.B1(n_16),
.B2(n_28),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_89),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_43),
.C(n_6),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_82),
.B(n_97),
.Y(n_128)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_92),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_87),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_40),
.Y(n_89)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_63),
.Y(n_92)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_94),
.Y(n_119)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_25),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_101),
.Y(n_138)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_32),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_108),
.Y(n_125)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_74),
.A2(n_35),
.B1(n_30),
.B2(n_32),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_35),
.B(n_16),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_28),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_28),
.Y(n_115)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_106),
.B1(n_37),
.B2(n_38),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_118),
.A2(n_126),
.B1(n_87),
.B2(n_96),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_45),
.B1(n_35),
.B2(n_44),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_136),
.B1(n_143),
.B2(n_86),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_40),
.C(n_64),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_144),
.C(n_147),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_83),
.A2(n_45),
.B1(n_19),
.B2(n_33),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_49),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_116),
.A2(n_25),
.B1(n_20),
.B2(n_22),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_93),
.A2(n_33),
.B(n_61),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_153),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_85),
.C(n_99),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_152),
.C(n_158),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_180),
.B1(n_123),
.B2(n_124),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_100),
.C(n_107),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_159),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_162),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_164),
.B1(n_181),
.B2(n_131),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_84),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_88),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_117),
.C(n_114),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_165),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_112),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_132),
.A2(n_91),
.B1(n_102),
.B2(n_94),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_65),
.C(n_110),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_65),
.C(n_49),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_172),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_128),
.B(n_20),
.Y(n_169)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_122),
.B(n_22),
.Y(n_170)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_146),
.B(n_25),
.Y(n_171)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_65),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_23),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_134),
.A2(n_98),
.B1(n_111),
.B2(n_33),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_177),
.B1(n_161),
.B2(n_120),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_127),
.B(n_22),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_111),
.B1(n_21),
.B2(n_27),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_119),
.B(n_21),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_178),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_129),
.A2(n_27),
.B1(n_21),
.B2(n_24),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_27),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_24),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_SL g183 ( 
.A1(n_152),
.A2(n_124),
.B(n_123),
.C(n_34),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_183),
.A2(n_203),
.B(n_211),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_SL g228 ( 
.A1(n_185),
.A2(n_193),
.B(n_173),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_121),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_186),
.B(n_207),
.C(n_212),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_189),
.B(n_195),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_157),
.A2(n_145),
.B1(n_141),
.B2(n_131),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_194),
.A2(n_165),
.B1(n_179),
.B2(n_150),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_149),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_164),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_209),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_199),
.A2(n_210),
.B1(n_7),
.B2(n_14),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_145),
.B1(n_120),
.B2(n_130),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_166),
.B1(n_175),
.B2(n_153),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_34),
.B(n_31),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_31),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_208),
.B(n_0),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_163),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_177),
.A2(n_24),
.B1(n_31),
.B2(n_105),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_31),
.B(n_1),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_81),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_156),
.Y(n_217)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_217),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_206),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_218),
.B(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_187),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_230),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

AO32x1_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_199),
.A3(n_211),
.B1(n_215),
.B2(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_228),
.B1(n_241),
.B2(n_183),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_202),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_231),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_8),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_239),
.C(n_213),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_202),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_233),
.A2(n_240),
.B1(n_227),
.B2(n_222),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_8),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_1),
.C(n_2),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_198),
.A2(n_203),
.B1(n_183),
.B2(n_196),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_186),
.B(n_1),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_242),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_9),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_243),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_198),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_247),
.C(n_254),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_265),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_196),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_239),
.C(n_219),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_226),
.A2(n_210),
.B1(n_201),
.B2(n_191),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_232),
.C(n_207),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_216),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_257),
.A2(n_10),
.B(n_11),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_201),
.B1(n_192),
.B2(n_3),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_1),
.C(n_2),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_264),
.C(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_3),
.C(n_4),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_217),
.B(n_242),
.Y(n_265)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_279),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_276),
.C(n_278),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_225),
.B1(n_221),
.B2(n_223),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

FAx1_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_234),
.CI(n_238),
.CON(n_271),
.SN(n_271)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_263),
.B(n_258),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_250),
.Y(n_272)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_273),
.B(n_264),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_218),
.B1(n_231),
.B2(n_236),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_274),
.B(n_282),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_234),
.C(n_240),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_3),
.C(n_5),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_6),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_248),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_259),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_246),
.C(n_252),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_253),
.Y(n_297)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_284),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_288),
.B(n_297),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_246),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_268),
.C(n_281),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_277),
.A2(n_263),
.B(n_256),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_295),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_294),
.A2(n_271),
.B1(n_280),
.B2(n_268),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_256),
.B(n_260),
.Y(n_295)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_273),
.B(n_255),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_278),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_302),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_299),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_292),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_309),
.C(n_311),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_291),
.B(n_290),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_280),
.C(n_271),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_12),
.C(n_14),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_15),
.C(n_5),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_314),
.C(n_294),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_15),
.C(n_5),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_320),
.Y(n_330)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_318),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_301),
.Y(n_319)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_288),
.C(n_286),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_296),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_321),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_SL g322 ( 
.A1(n_306),
.A2(n_287),
.B(n_291),
.C(n_286),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_314),
.Y(n_326)
);

AOI21xp33_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_312),
.B(n_15),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_313),
.B1(n_304),
.B2(n_311),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_317),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_316),
.Y(n_331)
);

AOI21xp33_ASAP7_75t_L g334 ( 
.A1(n_328),
.A2(n_326),
.B(n_330),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_322),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_334),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_329),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_337),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_335),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_339),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_340),
.B(n_327),
.Y(n_341)
);


endmodule