module fake_aes_2961_n_40 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
wire n_39;
OA21x2_ASAP7_75t_L g11 ( .A1(n_6), .A2(n_4), .B(n_0), .Y(n_11) );
NOR2xp67_ASAP7_75t_L g12 ( .A(n_0), .B(n_10), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_9), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_7), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_5), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_17), .B(n_1), .Y(n_18) );
AOI22xp33_ASAP7_75t_SL g19 ( .A1(n_17), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_19) );
NOR2xp33_ASAP7_75t_L g20 ( .A(n_14), .B(n_4), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_14), .B(n_5), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_15), .B(n_8), .Y(n_22) );
NOR2xp33_ASAP7_75t_L g23 ( .A(n_18), .B(n_13), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_20), .A2(n_15), .B1(n_16), .B2(n_11), .Y(n_24) );
OR2x6_ASAP7_75t_L g25 ( .A(n_21), .B(n_16), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_22), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
OAI221xp5_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_19), .B1(n_20), .B2(n_11), .C(n_12), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_27), .B(n_25), .Y(n_31) );
OAI22xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_29), .B1(n_28), .B2(n_24), .Y(n_32) );
INVx2_ASAP7_75t_L g33 ( .A(n_30), .Y(n_33) );
AOI22xp33_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_31), .B1(n_23), .B2(n_11), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_33), .B(n_31), .Y(n_35) );
XOR2xp5_ASAP7_75t_L g36 ( .A(n_32), .B(n_31), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
NOR3xp33_ASAP7_75t_L g38 ( .A(n_36), .B(n_12), .C(n_11), .Y(n_38) );
NOR3x2_ASAP7_75t_L g39 ( .A(n_38), .B(n_11), .C(n_7), .Y(n_39) );
AOI22xp5_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_34), .B1(n_37), .B2(n_6), .Y(n_40) );
endmodule