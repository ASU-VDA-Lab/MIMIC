module fake_jpeg_22486_n_171 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_171);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_33),
.B(n_41),
.Y(n_67)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_2),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_15),
.B(n_3),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_3),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_23),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_28),
.B1(n_17),
.B2(n_20),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_47),
.A2(n_48),
.B1(n_60),
.B2(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_17),
.B1(n_26),
.B2(n_21),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_49),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_14),
.B1(n_34),
.B2(n_21),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_66),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_68),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_20),
.B1(n_21),
.B2(n_26),
.Y(n_60)
);

AO21x1_ASAP7_75t_SL g96 ( 
.A1(n_62),
.A2(n_31),
.B(n_25),
.Y(n_96)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_71),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_26),
.Y(n_66)
);

OR2x2_ASAP7_75t_SL g68 ( 
.A(n_37),
.B(n_14),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_29),
.Y(n_87)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_15),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_74),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_35),
.A2(n_20),
.B1(n_19),
.B2(n_27),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_36),
.A2(n_15),
.B1(n_27),
.B2(n_25),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_4),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_66),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_23),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_77),
.B(n_78),
.Y(n_121)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_50),
.B(n_29),
.Y(n_79)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_92),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_16),
.C(n_24),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_65),
.C(n_59),
.Y(n_112)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_96),
.C(n_99),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_16),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_67),
.B(n_31),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_19),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_66),
.B1(n_75),
.B2(n_61),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_75),
.B1(n_47),
.B2(n_48),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_62),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_120),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_57),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_90),
.C(n_91),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_53),
.B(n_55),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_100),
.B(n_92),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_81),
.A2(n_60),
.B1(n_55),
.B2(n_65),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_113),
.C(n_116),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_4),
.Y(n_113)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_82),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_84),
.C(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_5),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_129),
.B(n_112),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_126),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_94),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_128),
.C(n_133),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_86),
.C(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_86),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_138),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_83),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_132),
.B(n_135),
.Y(n_140)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_96),
.B(n_83),
.C(n_101),
.D(n_76),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_5),
.B(n_6),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_110),
.B(n_102),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_6),
.Y(n_135)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_6),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_143),
.A2(n_147),
.B(n_122),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_111),
.B1(n_106),
.B2(n_121),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_125),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_154),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_150),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_155),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_128),
.C(n_108),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_140),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_156),
.A2(n_141),
.B(n_144),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_146),
.B(n_149),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_161),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_156),
.A2(n_147),
.B(n_145),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_159),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_158),
.A2(n_157),
.B1(n_148),
.B2(n_139),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_160),
.B1(n_104),
.B2(n_117),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_142),
.B(n_114),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_167),
.C(n_11),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_9),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_168),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_12),
.Y(n_171)
);


endmodule