module fake_netlist_5_1810_n_4989 (n_137, n_294, n_431, n_318, n_380, n_419, n_611, n_444, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_515, n_57, n_353, n_351, n_367, n_620, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_629, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_600, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_50, n_337, n_430, n_313, n_631, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_613, n_241, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_4989);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_611;
input n_444;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_600;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_613;
input n_241;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_4989;

wire n_924;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_977;
wire n_4706;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_790;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_2395;
wire n_2347;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_671;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_1462;
wire n_4211;
wire n_3448;
wire n_3019;
wire n_2096;
wire n_877;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_1696;
wire n_2483;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_1860;
wire n_4615;
wire n_1107;
wire n_1728;
wire n_2076;
wire n_668;
wire n_2147;
wire n_3010;
wire n_2770;
wire n_4131;
wire n_2584;
wire n_3188;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_1242;
wire n_3283;
wire n_2323;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_731;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_3214;
wire n_1517;
wire n_2091;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_1449;
wire n_4678;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_3947;
wire n_3490;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_2384;
wire n_882;
wire n_3156;
wire n_696;
wire n_3376;
wire n_646;
wire n_4468;
wire n_3653;
wire n_3702;
wire n_1040;
wire n_4976;
wire n_2202;
wire n_2648;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_2276;
wire n_2089;
wire n_3420;
wire n_1561;
wire n_1165;
wire n_1034;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_845;
wire n_4255;
wire n_1796;
wire n_901;
wire n_4484;
wire n_3668;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_637;
wire n_2079;
wire n_2238;
wire n_1151;
wire n_1405;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_2859;
wire n_1075;
wire n_3395;
wire n_4917;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_2968;
wire n_1585;
wire n_2684;
wire n_3593;
wire n_1599;
wire n_4421;
wire n_4836;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_4532;
wire n_3339;
wire n_3349;
wire n_3735;
wire n_2248;
wire n_3007;
wire n_1000;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_2100;
wire n_3487;
wire n_3310;
wire n_2258;
wire n_748;
wire n_1667;
wire n_1058;
wire n_838;
wire n_3983;
wire n_1053;
wire n_1224;
wire n_4405;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_1014;
wire n_4969;
wire n_1241;
wire n_4504;
wire n_1385;
wire n_793;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_2987;
wire n_1527;
wire n_4567;
wire n_4164;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_2175;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_4471;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_3208;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_3649;
wire n_4302;
wire n_2514;
wire n_4786;
wire n_3257;
wire n_1027;
wire n_4160;
wire n_2293;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_1276;
wire n_1412;
wire n_3981;
wire n_1199;
wire n_1038;
wire n_1841;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_870;
wire n_1711;
wire n_1891;
wire n_3526;
wire n_2546;
wire n_965;
wire n_3790;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_4028;
wire n_1690;
wire n_3819;
wire n_2449;
wire n_1194;
wire n_2297;
wire n_4186;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2876;
wire n_4099;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2479;
wire n_1464;
wire n_4295;
wire n_649;
wire n_1444;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_3068;
wire n_2871;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_3317;
wire n_1121;
wire n_4391;
wire n_949;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1001;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_3455;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_1994;
wire n_1195;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_2796;
wire n_757;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_3095;
wire n_2805;
wire n_1145;
wire n_4918;
wire n_1153;
wire n_3856;
wire n_741;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_1207;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_2857;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_940;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_2947;
wire n_978;
wire n_4299;
wire n_4801;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_3378;
wire n_1431;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_660;
wire n_4294;
wire n_1732;
wire n_4125;
wire n_4232;
wire n_4949;
wire n_2941;
wire n_2457;
wire n_4790;
wire n_962;
wire n_723;
wire n_2536;
wire n_1336;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_3058;
wire n_4365;
wire n_1878;
wire n_3505;
wire n_4610;
wire n_3730;
wire n_4489;
wire n_974;
wire n_727;
wire n_4967;
wire n_957;
wire n_3001;
wire n_3945;
wire n_4542;
wire n_2261;
wire n_2729;
wire n_3597;
wire n_1612;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_4534;
wire n_4500;
wire n_3185;
wire n_1300;
wire n_1127;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_4329;
wire n_1006;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_2231;
wire n_2017;
wire n_2604;
wire n_4257;
wire n_3453;
wire n_2390;
wire n_3213;
wire n_1041;
wire n_3077;
wire n_1562;
wire n_3474;
wire n_3984;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_4189;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_860;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_948;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_4037;
wire n_2922;
wire n_3499;
wire n_3275;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_1552;
wire n_3618;
wire n_2593;
wire n_3683;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_824;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_815;
wire n_4594;
wire n_3424;
wire n_1381;
wire n_1037;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_3171;
wire n_1437;
wire n_645;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_1123;
wire n_1467;
wire n_2163;
wire n_634;
wire n_2254;
wire n_1382;
wire n_925;
wire n_3546;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_950;
wire n_4443;
wire n_4507;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_3244;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_912;
wire n_968;
wire n_4452;
wire n_4348;
wire n_4355;
wire n_3494;
wire n_885;
wire n_2125;
wire n_3771;
wire n_683;
wire n_3110;
wire n_1057;
wire n_1051;
wire n_721;
wire n_1157;
wire n_3073;
wire n_4572;
wire n_802;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_1305;
wire n_3178;
wire n_873;
wire n_2334;
wire n_690;
wire n_4521;
wire n_4488;
wire n_2289;
wire n_3051;
wire n_1343;
wire n_2783;
wire n_2263;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_4519;
wire n_3715;
wire n_972;
wire n_3040;
wire n_1938;
wire n_1200;
wire n_2499;
wire n_3568;
wire n_3737;
wire n_1185;
wire n_991;
wire n_1967;
wire n_1329;
wire n_3255;
wire n_4856;
wire n_2997;
wire n_4400;
wire n_943;
wire n_3326;
wire n_3734;
wire n_650;
wire n_4778;
wire n_2429;
wire n_883;
wire n_856;
wire n_1793;
wire n_4352;
wire n_4441;
wire n_918;
wire n_4761;
wire n_942;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_2094;
wire n_1096;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_3831;
wire n_3801;
wire n_2043;
wire n_2751;
wire n_4893;
wire n_1549;
wire n_1934;
wire n_4948;
wire n_4000;
wire n_655;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_1807;
wire n_2618;
wire n_2559;
wire n_763;
wire n_4748;
wire n_2295;
wire n_3931;
wire n_1219;
wire n_4010;
wire n_2840;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_2795;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_789;
wire n_4247;
wire n_4933;
wire n_4018;
wire n_3900;
wire n_1105;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_3872;
wire n_4336;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_836;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_3877;
wire n_2995;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_1102;
wire n_4052;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_2633;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_1164;
wire n_2097;
wire n_4304;
wire n_3911;
wire n_1303;
wire n_4431;
wire n_4192;
wire n_3736;
wire n_4805;
wire n_4885;
wire n_1661;
wire n_3565;
wire n_4701;
wire n_2575;
wire n_861;
wire n_1658;
wire n_1904;
wire n_1345;
wire n_1899;
wire n_1003;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_1726;
wire n_4631;
wire n_3035;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_3639;
wire n_708;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_1915;
wire n_1109;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_1399;
wire n_1979;
wire n_2924;
wire n_4111;
wire n_2484;
wire n_808;
wire n_797;
wire n_1025;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_4538;
wire n_766;
wire n_1117;
wire n_2754;
wire n_687;
wire n_1742;
wire n_2489;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_2866;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_827;
wire n_4878;
wire n_1703;
wire n_1650;
wire n_1137;
wire n_3934;
wire n_4985;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_653;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_850;
wire n_3074;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_3768;
wire n_2861;
wire n_1372;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_4022;
wire n_1531;
wire n_840;
wire n_1334;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_2817;
wire n_3139;
wire n_2598;
wire n_4601;
wire n_2687;
wire n_1120;
wire n_1890;
wire n_714;
wire n_4220;
wire n_1944;
wire n_909;
wire n_1497;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_1889;
wire n_1489;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_1569;
wire n_2188;
wire n_756;
wire n_1429;
wire n_4644;
wire n_4456;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_2898;
wire n_2717;
wire n_1861;
wire n_760;
wire n_3691;
wire n_3628;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_2573;
wire n_4435;
wire n_2939;
wire n_3807;
wire n_2447;
wire n_4764;
wire n_886;
wire n_1221;
wire n_2774;
wire n_1707;
wire n_853;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_751;
wire n_4827;
wire n_2488;
wire n_3477;
wire n_2476;
wire n_704;
wire n_4399;
wire n_2781;
wire n_2778;
wire n_771;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_2691;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_2526;
wire n_2703;
wire n_2167;
wire n_3391;
wire n_4259;
wire n_2709;
wire n_816;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_1339;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_2173;
wire n_1842;
wire n_871;
wire n_3738;
wire n_685;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_1555;
wire n_3245;
wire n_4417;
wire n_4899;
wire n_796;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1012;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_740;
wire n_3509;
wire n_3352;
wire n_3076;
wire n_3535;
wire n_2182;
wire n_1061;
wire n_3251;
wire n_2931;
wire n_1193;
wire n_3118;
wire n_3511;
wire n_1226;
wire n_3443;
wire n_2146;
wire n_1487;
wire n_3644;
wire n_3336;
wire n_3935;
wire n_781;
wire n_3521;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_3114;
wire n_3125;
wire n_4981;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_4430;
wire n_4081;
wire n_1103;
wire n_3132;
wire n_4407;
wire n_648;
wire n_3951;
wire n_4894;
wire n_3238;
wire n_3210;
wire n_2036;
wire n_3267;
wire n_695;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_3884;
wire n_3726;
wire n_805;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_3577;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_1160;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_1074;
wire n_3347;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_1448;
wire n_4288;
wire n_3567;
wire n_1634;
wire n_3939;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_666;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_2920;
wire n_4265;
wire n_1186;
wire n_1018;
wire n_2247;
wire n_713;
wire n_1622;
wire n_1180;
wire n_3705;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_2268;
wire n_3778;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_3795;
wire n_4419;
wire n_4477;
wire n_3179;
wire n_3256;
wire n_667;
wire n_2386;
wire n_1501;
wire n_3086;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_1099;
wire n_2568;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_1021;
wire n_4639;
wire n_3713;
wire n_3663;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_819;
wire n_2302;
wire n_951;
wire n_1494;
wire n_2069;
wire n_3434;
wire n_1806;
wire n_933;
wire n_1563;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_755;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_2482;
wire n_2677;
wire n_3832;
wire n_3987;
wire n_902;
wire n_1698;
wire n_2329;
wire n_1098;
wire n_2142;
wire n_3332;
wire n_1135;
wire n_3048;
wire n_3937;
wire n_2203;
wire n_4525;
wire n_1243;
wire n_3782;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_3786;
wire n_2888;
wire n_3638;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_3022;
wire n_4264;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_2149;
wire n_1078;
wire n_3060;
wire n_4276;
wire n_3013;
wire n_1984;
wire n_2408;
wire n_1877;
wire n_3049;
wire n_1723;
wire n_4485;
wire n_4626;
wire n_1036;
wire n_1097;
wire n_798;
wire n_2659;
wire n_1414;
wire n_4975;
wire n_1852;
wire n_3089;
wire n_2470;
wire n_3985;
wire n_1391;
wire n_670;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_663;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_813;
wire n_1284;
wire n_3440;
wire n_1748;
wire n_4569;
wire n_2699;
wire n_4897;
wire n_888;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_2615;
wire n_3940;
wire n_1064;
wire n_858;
wire n_2985;
wire n_691;
wire n_2753;
wire n_1582;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_3141;
wire n_3164;
wire n_3570;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_3936;
wire n_4503;
wire n_3507;
wire n_3821;
wire n_2700;
wire n_1211;
wire n_3367;
wire n_4464;
wire n_907;
wire n_3096;
wire n_3496;
wire n_4114;
wire n_989;
wire n_2544;
wire n_2356;
wire n_892;
wire n_4556;
wire n_2620;
wire n_1581;
wire n_4089;
wire n_2919;
wire n_4327;
wire n_953;
wire n_4218;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_963;
wire n_1052;
wire n_954;
wire n_4353;
wire n_2042;
wire n_884;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_1856;
wire n_4959;
wire n_4161;
wire n_832;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_2462;
wire n_1532;
wire n_3625;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_686;
wire n_2837;
wire n_847;
wire n_4844;
wire n_2979;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_702;
wire n_2548;
wire n_822;
wire n_2108;
wire n_3640;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_1779;
wire n_4738;
wire n_1369;
wire n_3909;
wire n_3207;
wire n_3944;
wire n_809;
wire n_4434;
wire n_4837;
wire n_3042;
wire n_1942;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_2222;
wire n_3510;
wire n_3218;
wire n_2667;
wire n_3150;
wire n_747;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_851;
wire n_843;
wire n_705;
wire n_3775;
wire n_4133;
wire n_678;
wire n_4184;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_2181;
wire n_1829;
wire n_4030;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_4820;
wire n_3770;
wire n_1308;
wire n_4938;
wire n_4179;
wire n_3469;
wire n_677;
wire n_2723;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_3855;
wire n_1008;
wire n_2054;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_3158;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_3113;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_4404;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_878;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_906;
wire n_919;
wire n_4356;
wire n_658;
wire n_2061;
wire n_4432;
wire n_2378;
wire n_1740;
wire n_1586;
wire n_4291;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_3545;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1095;
wire n_1614;
wire n_2339;
wire n_4637;
wire n_4935;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_3741;
wire n_3410;
wire n_2029;
wire n_995;
wire n_1609;
wire n_1887;
wire n_4413;
wire n_1073;
wire n_2346;
wire n_662;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_1215;
wire n_1592;
wire n_2882;
wire n_1721;
wire n_2338;
wire n_3672;
wire n_3197;
wire n_3109;
wire n_2721;
wire n_1043;
wire n_3002;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_2081;
wire n_4570;
wire n_2156;
wire n_4296;
wire n_1820;
wire n_2418;
wire n_2179;
wire n_1416;
wire n_1724;
wire n_2521;
wire n_3458;
wire n_1420;
wire n_1132;
wire n_3330;
wire n_4606;
wire n_4774;
wire n_2477;
wire n_3887;
wire n_4093;
wire n_1486;
wire n_4672;
wire n_3519;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_4766;
wire n_2896;
wire n_652;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_1349;
wire n_4460;
wire n_1031;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_834;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1965;
wire n_1902;
wire n_1941;
wire n_3938;
wire n_2878;
wire n_874;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_3189;
wire n_2066;
wire n_993;
wire n_3154;
wire n_1551;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4349;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1084;
wire n_970;
wire n_1935;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_1205;
wire n_3242;
wire n_3525;
wire n_3486;
wire n_2405;
wire n_3995;
wire n_2088;
wire n_2953;
wire n_4036;
wire n_921;
wire n_1795;
wire n_2578;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_2656;
wire n_1080;
wire n_1274;
wire n_3524;
wire n_1708;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2092;
wire n_2075;
wire n_3658;
wire n_1776;
wire n_4807;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_890;
wire n_1919;
wire n_960;
wire n_4230;
wire n_3419;
wire n_1290;
wire n_1047;
wire n_2053;
wire n_1958;
wire n_1252;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_1808;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_967;
wire n_2731;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_3979;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_4840;
wire n_3162;
wire n_983;
wire n_2760;
wire n_3377;
wire n_3749;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_762;
wire n_1283;
wire n_2637;
wire n_4384;
wire n_4423;
wire n_4096;
wire n_2881;
wire n_1203;
wire n_3282;
wire n_821;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_2475;
wire n_4598;
wire n_4478;
wire n_2646;
wire n_1605;
wire n_1228;
wire n_3920;
wire n_4890;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_828;
wire n_779;
wire n_4106;
wire n_3717;
wire n_2743;
wire n_2675;
wire n_1439;
wire n_3052;
wire n_945;
wire n_3743;
wire n_1932;
wire n_4721;
wire n_984;
wire n_694;
wire n_1983;
wire n_4029;
wire n_1594;
wire n_900;
wire n_3870;
wire n_4496;
wire n_3529;
wire n_1147;
wire n_1977;
wire n_2153;
wire n_4338;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_1470;
wire n_1735;
wire n_2318;
wire n_833;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_1201;
wire n_1114;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_669;
wire n_1176;
wire n_1149;
wire n_1020;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_2446;
wire n_3488;
wire n_1035;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_661;
wire n_4668;
wire n_4953;
wire n_3898;
wire n_849;
wire n_1786;
wire n_4274;
wire n_2627;
wire n_4759;
wire n_1413;
wire n_801;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_3552;
wire n_875;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_2361;
wire n_1173;
wire n_1603;
wire n_1401;
wire n_969;
wire n_4113;
wire n_1019;
wire n_1998;
wire n_4686;
wire n_3759;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_3933;
wire n_3206;
wire n_3966;
wire n_1702;
wire n_4183;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4872;
wire n_4233;
wire n_3192;
wire n_3764;
wire n_4709;
wire n_2649;
wire n_1187;
wire n_1929;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_1174;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_2252;
wire n_4819;
wire n_1685;
wire n_917;
wire n_1714;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_3390;
wire n_1573;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_1737;
wire n_774;
wire n_2493;
wire n_4930;
wire n_1059;
wire n_1133;
wire n_4537;
wire n_2885;
wire n_3318;
wire n_4070;
wire n_4282;
wire n_3485;
wire n_4180;
wire n_665;
wire n_3839;
wire n_1440;
wire n_3333;
wire n_2845;
wire n_4143;
wire n_4659;
wire n_2602;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_1812;
wire n_4105;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_2401;
wire n_3135;
wire n_2003;
wire n_1457;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3438;
wire n_4098;
wire n_872;
wire n_1297;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_1184;
wire n_2184;
wire n_985;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_676;
wire n_4442;
wire n_4698;
wire n_642;
wire n_1602;
wire n_1178;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_3397;
wire n_3740;
wire n_1081;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_703;
wire n_1318;
wire n_780;
wire n_2977;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_3600;
wire n_4134;
wire n_1388;
wire n_2836;
wire n_672;
wire n_1625;
wire n_2130;
wire n_898;
wire n_3239;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_4740;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_4049;
wire n_941;
wire n_3862;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_4724;
wire n_1238;
wire n_1772;
wire n_752;
wire n_1476;
wire n_1108;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_862;
wire n_3584;
wire n_3756;
wire n_2889;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_2260;
wire n_1813;
wire n_4833;
wire n_3056;
wire n_2345;
wire n_1172;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_3289;
wire n_1973;
wire n_786;
wire n_1142;
wire n_2579;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2984;
wire n_3364;
wire n_1873;
wire n_3201;
wire n_1087;
wire n_3472;
wire n_2874;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_4968;
wire n_1272;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_3050;
wire n_1478;
wire n_3903;
wire n_4834;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_4171;
wire n_4045;
wire n_1367;
wire n_4562;
wire n_3634;
wire n_1460;
wire n_2834;
wire n_2531;
wire n_2702;
wire n_2030;
wire n_903;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_2234;
wire n_4804;
wire n_2209;
wire n_4270;
wire n_2797;
wire n_1255;
wire n_2321;
wire n_722;
wire n_3680;
wire n_844;
wire n_3497;
wire n_1601;
wire n_2940;
wire n_2612;
wire n_1495;
wire n_4566;
wire n_979;
wire n_2841;
wire n_3322;
wire n_4576;
wire n_846;
wire n_2427;
wire n_2505;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_2594;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_3112;
wire n_2349;
wire n_1379;
wire n_3874;
wire n_4676;
wire n_4544;
wire n_2170;
wire n_1091;
wire n_641;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_3266;
wire n_4646;
wire n_1130;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_2426;
wire n_657;
wire n_4320;
wire n_4881;
wire n_3613;
wire n_3444;
wire n_1181;
wire n_1505;
wire n_4012;
wire n_651;
wire n_4636;
wire n_4584;
wire n_807;
wire n_3910;
wire n_4711;
wire n_835;
wire n_3319;
wire n_3335;
wire n_3413;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_1138;
wire n_927;
wire n_2689;
wire n_3259;
wire n_4191;
wire n_4293;
wire n_2010;
wire n_3688;
wire n_3016;
wire n_1693;
wire n_2599;
wire n_904;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_1271;
wire n_1542;
wire n_1423;
wire n_1166;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2200;
wire n_3261;
wire n_1161;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_1150;
wire n_3127;
wire n_1780;
wire n_3732;
wire n_4250;
wire n_1055;
wire n_3596;
wire n_4699;
wire n_3906;
wire n_4127;
wire n_880;
wire n_3297;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_4202;
wire n_2853;
wire n_1323;
wire n_688;
wire n_3766;
wire n_1353;
wire n_800;
wire n_2880;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_4038;
wire n_4109;
wire n_915;
wire n_864;
wire n_1264;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_3621;
wire n_1580;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1607;
wire n_2538;
wire n_2105;
wire n_3163;
wire n_1118;
wire n_1686;
wire n_947;
wire n_3710;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_1230;
wire n_4144;
wire n_2165;
wire n_929;
wire n_3379;
wire n_4374;
wire n_3532;
wire n_1124;
wire n_2127;
wire n_1818;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1257;
wire n_1182;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_4548;
wire n_3258;
wire n_4622;
wire n_1016;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_4816;
wire n_1483;
wire n_2983;
wire n_3810;
wire n_1289;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_4483;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_2651;
wire n_4358;
wire n_3656;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1374;
wire n_4793;
wire n_4168;
wire n_3446;
wire n_955;
wire n_3028;
wire n_4806;
wire n_1146;
wire n_4350;
wire n_897;
wire n_1428;
wire n_1216;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1931;
wire n_4187;
wire n_1070;
wire n_4166;
wire n_1030;
wire n_3222;
wire n_1071;
wire n_1267;
wire n_1801;
wire n_1513;
wire n_2970;
wire n_2235;
wire n_673;
wire n_837;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_680;
wire n_1473;
wire n_3755;
wire n_4258;
wire n_4498;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_3563;
wire n_2506;
wire n_675;
wire n_4064;
wire n_4936;
wire n_1556;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_2944;
wire n_881;
wire n_2407;
wire n_4907;
wire n_3262;
wire n_1450;
wire n_4006;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_889;
wire n_2358;
wire n_973;
wire n_3716;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_736;
wire n_2750;
wire n_3899;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_2557;
wire n_1248;
wire n_4850;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_2590;
wire n_2330;
wire n_2942;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_944;
wire n_3889;
wire n_4256;
wire n_4224;
wire n_3508;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_857;
wire n_2636;
wire n_1951;
wire n_1825;
wire n_1883;
wire n_2759;
wire n_4415;
wire n_4702;
wire n_4252;
wire n_4457;
wire n_971;
wire n_1393;
wire n_2319;
wire n_3481;
wire n_2808;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_4491;
wire n_2930;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_1662;
wire n_1481;
wire n_4001;
wire n_3047;
wire n_868;
wire n_2454;
wire n_4371;
wire n_914;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_4194;
wire n_759;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1766;
wire n_1571;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_4082;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_3279;
wire n_2621;
wire n_1537;
wire n_4262;
wire n_2671;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_1647;
wire n_4685;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_4014;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_1233;
wire n_1615;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_1333;
wire n_1443;
wire n_1539;
wire n_946;
wire n_4892;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_689;
wire n_738;
wire n_1624;
wire n_4970;
wire n_640;
wire n_3816;
wire n_1279;
wire n_4108;
wire n_4486;
wire n_2960;
wire n_1090;
wire n_633;
wire n_4627;
wire n_758;
wire n_2290;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_1049;
wire n_2145;
wire n_1639;
wire n_1068;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_2039;
wire n_4961;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_3396;
wire n_1445;
wire n_4023;
wire n_4420;
wire n_1923;
wire n_1017;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1828;
wire n_2320;
wire n_1045;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_1033;
wire n_4396;
wire n_636;
wire n_4367;
wire n_2087;
wire n_1009;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_1578;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_2725;
wire n_3883;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_773;
wire n_743;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_3466;
wire n_4962;
wire n_1237;
wire n_2595;
wire n_761;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_3586;
wire n_1390;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_3065;
wire n_4361;
wire n_1093;
wire n_4614;
wire n_1265;
wire n_2681;
wire n_3103;
wire n_765;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_1015;
wire n_1651;
wire n_2775;
wire n_4693;
wire n_1101;
wire n_1106;
wire n_4326;
wire n_3557;
wire n_2230;
wire n_4744;
wire n_2851;
wire n_4305;
wire n_1455;
wire n_767;
wire n_2490;
wire n_1407;
wire n_4213;
wire n_2849;
wire n_3692;
wire n_2204;
wire n_4929;
wire n_729;
wire n_1961;
wire n_4964;
wire n_911;
wire n_1430;
wire n_4802;
wire n_1354;
wire n_4139;
wire n_1044;
wire n_3029;
wire n_2508;
wire n_4031;
wire n_2416;
wire n_3881;
wire n_2461;
wire n_2243;
wire n_4583;
wire n_4210;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_2890;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_716;
wire n_1630;
wire n_4891;
wire n_701;
wire n_1023;
wire n_803;
wire n_1092;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_3993;
wire n_4940;
wire n_1056;
wire n_3588;
wire n_2308;
wire n_4590;
wire n_4830;
wire n_4664;
wire n_3860;
wire n_1029;
wire n_1206;
wire n_3160;
wire n_2191;
wire n_2428;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_1060;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_4297;
wire n_1632;
wire n_1085;
wire n_1066;
wire n_3800;
wire n_2403;
wire n_4608;
wire n_2792;
wire n_2870;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_4172;
wire n_4791;
wire n_4536;
wire n_2463;
wire n_4773;
wire n_4497;
wire n_2472;
wire n_4611;
wire n_4755;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_1560;
wire n_4362;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_4422;
wire n_2589;
wire n_1363;
wire n_1301;
wire n_3482;
wire n_2233;
wire n_1312;
wire n_804;
wire n_4555;
wire n_2827;
wire n_1504;
wire n_3956;
wire n_3572;
wire n_992;
wire n_4215;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_842;
wire n_2082;
wire n_1643;
wire n_3167;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3854;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3078;
wire n_894;
wire n_3253;
wire n_4027;
wire n_2280;
wire n_831;
wire n_4599;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_1881;
wire n_988;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_3950;
wire n_4458;
wire n_4121;
wire n_1616;
wire n_4476;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_4860;
wire n_4359;
wire n_635;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_1848;
wire n_2126;
wire n_4573;
wire n_4118;
wire n_4803;
wire n_4079;
wire n_4091;
wire n_681;
wire n_1638;
wire n_2002;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_830;
wire n_3085;
wire n_1655;
wire n_749;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_4316;
wire n_939;
wire n_3697;
wire n_1232;
wire n_734;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_2711;
wire n_1653;
wire n_1506;
wire n_990;
wire n_2867;
wire n_1894;
wire n_975;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_4253;
wire n_2608;
wire n_2657;
wire n_770;
wire n_2852;
wire n_2392;
wire n_711;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_1516;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_3402;
wire n_4679;
wire n_4115;
wire n_726;
wire n_2988;
wire n_1731;
wire n_818;
wire n_1970;
wire n_2766;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_1993;
wire n_3835;
wire n_2205;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_1912;
wire n_3401;
wire n_3226;
wire n_1410;
wire n_707;
wire n_3902;
wire n_4730;
wire n_937;
wire n_2779;
wire n_1584;
wire n_3654;
wire n_2164;
wire n_2115;
wire n_2232;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_2811;
wire n_3348;
wire n_895;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_1543;
wire n_1991;
wire n_2224;
wire n_732;
wire n_4743;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_2692;
wire n_2008;
wire n_4654;
wire n_799;
wire n_1213;
wire n_4733;
wire n_3792;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_869;
wire n_3312;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_3285;
wire n_3968;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_684;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_664;
wire n_2480;
wire n_2363;
wire n_643;
wire n_4072;
wire n_916;
wire n_1115;
wire n_4781;
wire n_3606;
wire n_2550;
wire n_4424;
wire n_823;
wire n_725;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_3878;
wire n_4450;
wire n_3553;
wire n_719;
wire n_4746;
wire n_1683;
wire n_1530;
wire n_997;
wire n_932;
wire n_3131;
wire n_1409;
wire n_3850;
wire n_788;
wire n_4459;
wire n_1268;
wire n_2996;
wire n_1320;
wire n_4050;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_1063;
wire n_4853;
wire n_981;
wire n_867;
wire n_2422;
wire n_2239;
wire n_2950;
wire n_3852;
wire n_812;
wire n_4520;
wire n_2057;
wire n_4008;
wire n_905;
wire n_782;
wire n_3858;
wire n_1901;
wire n_4502;
wire n_3032;
wire n_4851;
wire n_1330;
wire n_3072;
wire n_3313;
wire n_3081;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_769;
wire n_4571;
wire n_2006;
wire n_934;
wire n_1618;
wire n_826;
wire n_2343;
wire n_3439;
wire n_654;
wire n_2535;
wire n_4205;
wire n_2726;
wire n_4723;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_1083;
wire n_4739;
wire n_2376;
wire n_3017;
wire n_787;
wire n_2456;
wire n_3904;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_4879;
wire n_930;
wire n_3926;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_2764;
wire n_1498;
wire n_4225;
wire n_682;
wire n_2567;
wire n_3102;
wire n_922;
wire n_1648;
wire n_4153;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_839;
wire n_2964;
wire n_3769;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_2442;
wire n_928;
wire n_1943;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_1396;
wire n_1348;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_4839;
wire n_1028;
wire n_4016;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_632;
wire n_4231;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_4083;
wire n_1937;
wire n_4461;
wire n_3234;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_3512;
wire n_4939;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_2503;
wire n_1540;
wire n_1936;
wire n_2027;
wire n_2642;
wire n_720;
wire n_2500;
wire n_1918;
wire n_863;
wire n_4831;
wire n_2513;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_2414;
wire n_1402;
wire n_3662;
wire n_4319;
wire n_644;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_2004;
wire n_3694;
wire n_2586;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_1196;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_811;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_4474;
wire n_1089;
wire n_1004;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_2704;
wire n_4214;
wire n_4884;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_4580;
wire n_1263;
wire n_1126;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_1859;
wire n_1677;
wire n_2955;
wire n_4112;
wire n_4337;
wire n_4138;
wire n_1528;
wire n_1292;
wire n_2520;
wire n_1198;
wire n_956;
wire n_2134;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_3595;
wire n_1347;
wire n_4238;
wire n_1451;
wire n_1022;
wire n_1545;
wire n_2374;
wire n_859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_2396;
wire n_1799;
wire n_854;
wire n_4734;
wire n_674;
wire n_1939;
wire n_2486;
wire n_4635;
wire n_1152;
wire n_3501;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_4242;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_1705;
wire n_659;
wire n_4561;
wire n_2639;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_1261;
wire n_938;
wire n_3186;
wire n_4955;
wire n_1154;
wire n_4501;
wire n_3696;
wire n_1280;
wire n_3650;
wire n_2761;
wire n_3157;
wire n_709;
wire n_2537;
wire n_2144;
wire n_920;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_4197;
wire n_4829;
wire n_1949;
wire n_976;
wire n_1946;
wire n_2936;
wire n_775;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_2141;
wire n_4369;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_1850;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_2663;
wire n_1394;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_4944;
wire n_926;
wire n_2180;
wire n_2249;
wire n_4135;
wire n_1218;
wire n_2632;
wire n_1547;
wire n_777;
wire n_1755;
wire n_958;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_4716;
wire n_4942;
wire n_2432;
wire n_1521;
wire n_3405;
wire n_4745;
wire n_2337;
wire n_1167;
wire n_1384;
wire n_3907;
wire n_923;
wire n_4629;
wire n_2932;
wire n_2980;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_4752;
wire n_1750;
wire n_1459;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_4552;
wire n_3885;
wire n_2713;
wire n_2644;
wire n_1197;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_3427;
wire n_4067;
wire n_1403;
wire n_4042;
wire n_4176;
wire n_4385;
wire n_3320;
wire n_2688;
wire n_1202;
wire n_1463;
wire n_3651;
wire n_4333;
wire n_3359;
wire n_2865;
wire n_2706;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_4246;
wire n_3580;
wire n_2139;
wire n_4609;
wire n_2674;
wire n_1565;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_4462;
wire n_4472;
wire n_647;
wire n_3433;
wire n_1072;
wire n_2305;
wire n_2450;
wire n_3447;
wire n_3305;
wire n_4151;
wire n_4148;
wire n_1712;
wire n_3528;
wire n_4373;
wire n_4934;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_4630;
wire n_4643;
wire n_4331;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_1775;
wire n_3296;
wire n_1368;
wire n_2762;
wire n_4683;
wire n_728;
wire n_1162;
wire n_1847;
wire n_2767;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_3923;
wire n_931;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_639;
wire n_1629;
wire n_2801;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_1997;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_1259;
wire n_4553;
wire n_706;
wire n_746;
wire n_784;
wire n_3978;
wire n_4809;
wire n_1244;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_1788;
wire n_2491;
wire n_913;
wire n_3833;
wire n_865;
wire n_697;
wire n_1222;
wire n_1679;
wire n_4841;
wire n_776;
wire n_2022;
wire n_3814;
wire n_1415;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_3513;
wire n_3133;
wire n_4645;
wire n_1191;
wire n_2992;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_2517;
wire n_3128;
wire n_744;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_1529;
wire n_2469;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_3000;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1839;
wire n_1837;
wire n_4557;
wire n_4451;
wire n_2875;
wire n_936;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_3471;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_1656;
wire n_3564;
wire n_1158;
wire n_3988;
wire n_3457;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_3630;
wire n_3271;
wire n_4771;
wire n_908;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_724;
wire n_1781;
wire n_2084;
wire n_3648;
wire n_3075;
wire n_3173;
wire n_4692;
wire n_959;
wire n_3031;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_1169;
wire n_2666;
wire n_3385;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_2314;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_1079;
wire n_1593;
wire n_3767;
wire n_2299;
wire n_2873;
wire n_2540;
wire n_4589;
wire n_4578;
wire n_1640;
wire n_2162;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_742;
wire n_750;
wire n_2168;
wire n_2790;
wire n_3629;
wire n_3021;
wire n_2359;
wire n_3674;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_2312;
wire n_3015;
wire n_1171;
wire n_1920;
wire n_1065;
wire n_4147;
wire n_2048;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_1309;
wire n_4974;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_3276;
wire n_3787;
wire n_2124;
wire n_1119;
wire n_1240;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_4285;
wire n_4651;
wire n_700;
wire n_4818;
wire n_4514;
wire n_1366;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_1568;
wire n_2110;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_1591;
wire n_2033;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_1249;
wire n_1111;
wire n_2132;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_1140;
wire n_891;
wire n_3387;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_2831;
wire n_1456;
wire n_4882;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_987;
wire n_4545;
wire n_3037;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_1131;
wire n_2467;
wire n_1094;
wire n_2288;
wire n_4063;
wire n_1209;
wire n_3592;
wire n_4650;
wire n_4888;
wire n_1435;
wire n_879;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_1645;
wire n_4041;
wire n_2858;
wire n_4060;
wire n_996;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_3097;
wire n_4541;
wire n_3824;
wire n_3388;
wire n_4494;
wire n_3059;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_3589;
wire n_952;
wire n_2534;
wire n_1229;
wire n_4799;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_2789;
wire n_4775;
wire n_2216;
wire n_1897;
wire n_764;
wire n_1424;
wire n_2933;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_4455;
wire n_2328;
wire n_4248;
wire n_4754;
wire n_4554;
wire n_4845;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_1141;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_1432;
wire n_3875;
wire n_4003;
wire n_2402;
wire n_4301;
wire n_841;
wire n_1050;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_1844;
wire n_3777;
wire n_4784;
wire n_2999;
wire n_1644;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_3080;
wire n_4199;
wire n_2701;
wire n_3362;
wire n_1631;
wire n_3105;
wire n_1179;
wire n_753;
wire n_1048;
wire n_4286;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_692;
wire n_820;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_3417;
wire n_1143;
wire n_1579;
wire n_4034;
wire n_1688;
wire n_3327;
wire n_4689;
wire n_3067;
wire n_2755;
wire n_3237;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_3400;
wire n_4550;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_3382;
wire n_3574;
wire n_2169;
wire n_1557;
wire n_4201;
wire n_896;
wire n_3316;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_2192;
wire n_964;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_4416;
wire n_3372;
wire n_4539;
wire n_814;
wire n_2707;
wire n_2471;
wire n_1472;
wire n_1671;
wire n_3230;
wire n_1062;
wire n_3342;
wire n_4682;
wire n_3708;
wire n_1204;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_3861;
wire n_4736;
wire n_3780;
wire n_783;
wire n_1928;
wire n_1188;
wire n_3957;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_3608;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_4040;
wire n_2207;
wire n_2619;
wire n_2444;
wire n_1110;
wire n_3123;
wire n_1088;
wire n_3393;
wire n_638;
wire n_866;
wire n_4887;
wire n_4617;
wire n_3520;
wire n_2492;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_693;
wire n_4792;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_4290;
wire n_1375;
wire n_3727;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_1371;
wire n_4956;
wire n_2206;
wire n_3182;
wire n_2564;
wire n_4947;
wire n_876;
wire n_4656;
wire n_1190;
wire n_3896;
wire n_3958;
wire n_3450;
wire n_966;
wire n_4729;
wire n_4987;
wire n_4971;
wire n_1116;
wire n_2000;
wire n_1212;
wire n_2074;
wire n_3174;
wire n_982;
wire n_1453;
wire n_2217;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_3408;
wire n_899;
wire n_2722;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_1628;
wire n_3432;
wire n_1514;
wire n_1771;
wire n_1005;
wire n_679;
wire n_710;
wire n_3090;
wire n_1168;
wire n_2437;
wire n_3762;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_910;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_3972;
wire n_3308;
wire n_791;
wire n_1533;
wire n_4772;
wire n_3467;
wire n_4322;
wire n_1720;
wire n_2830;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_4677;
wire n_3901;
wire n_715;
wire n_1480;
wire n_3757;
wire n_3381;
wire n_1782;
wire n_2245;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_810;
wire n_2965;
wire n_3635;
wire n_1144;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_1170;
wire n_2213;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_855;
wire n_1461;
wire n_3204;
wire n_2136;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_3005;
wire n_1235;
wire n_4380;
wire n_980;
wire n_698;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1783;
wire n_2601;
wire n_3043;
wire n_998;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_4880;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_1417;
wire n_1295;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_1762;
wire n_1013;
wire n_718;
wire n_3023;
wire n_4193;
wire n_4075;
wire n_3104;
wire n_4737;
wire n_3647;
wire n_825;
wire n_2819;
wire n_737;
wire n_3609;
wire n_4136;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_3720;
wire n_4535;
wire n_733;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_4794;
wire n_3959;
wire n_792;
wire n_3140;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_4196;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_3069;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_3084;
wire n_1727;
wire n_2735;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_2411;
wire n_1046;
wire n_3761;
wire n_4889;
wire n_2014;
wire n_2986;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4828;
wire n_4558;
wire n_2172;
wire n_4722;
wire n_1129;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_961;
wire n_2250;
wire n_1225;
wire n_4092;
wire n_3908;
wire n_2423;
wire n_3671;
wire n_994;
wire n_3344;
wire n_2194;
wire n_848;
wire n_4465;
wire n_3302;
wire n_1223;
wire n_2680;
wire n_1567;
wire n_3122;
wire n_4808;
wire n_3842;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_1797;
wire n_2957;
wire n_2357;
wire n_1250;
wire n_3309;
wire n_772;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_2570;
wire n_1086;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_2744;
wire n_4287;
wire n_2397;
wire n_2208;
wire n_3063;
wire n_3617;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_1113;
wire n_1277;
wire n_2591;
wire n_3384;
wire n_852;
wire n_4602;
wire n_4449;
wire n_1864;
wire n_1337;
wire n_4445;
wire n_699;
wire n_1627;
wire n_1245;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_2278;
wire n_4915;
wire n_2135;
wire n_3493;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_1076;
wire n_2823;
wire n_1408;
wire n_1761;
wire n_730;
wire n_795;
wire n_4345;
wire n_3281;
wire n_656;
wire n_3307;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_1526;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_712;
wire n_1583;
wire n_2826;
wire n_3539;
wire n_1042;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_4124;
wire n_4492;
wire n_2708;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_3721;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1234;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_1032;
wire n_2614;
wire n_2991;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_3473;
wire n_4560;
wire n_2839;
wire n_1588;
wire n_2237;
wire n_3463;
wire n_3699;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_2728;
wire n_3857;

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_541),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_472),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_174),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_271),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_530),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_118),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_149),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_101),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_547),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_590),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_97),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_117),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_513),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_125),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_83),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_624),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_105),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_298),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_252),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_534),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_129),
.Y(n_652)
);

CKINVDCx16_ASAP7_75t_R g653 ( 
.A(n_239),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_402),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_209),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_231),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_403),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_5),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_62),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_126),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_296),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_367),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_334),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_124),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_564),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_298),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_475),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_254),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_337),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_122),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_124),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_309),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_416),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_137),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_7),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_211),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_286),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_199),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_556),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_300),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_77),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_247),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_279),
.Y(n_683)
);

BUFx5_ASAP7_75t_L g684 ( 
.A(n_378),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_463),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_329),
.Y(n_686)
);

BUFx10_ASAP7_75t_L g687 ( 
.A(n_312),
.Y(n_687)
);

CKINVDCx16_ASAP7_75t_R g688 ( 
.A(n_362),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_4),
.Y(n_689)
);

BUFx2_ASAP7_75t_SL g690 ( 
.A(n_157),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_463),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_119),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_434),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_282),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_418),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_332),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_612),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_430),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_223),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_366),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_433),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_23),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_167),
.Y(n_703)
);

CKINVDCx16_ASAP7_75t_R g704 ( 
.A(n_147),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_343),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_360),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_12),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_438),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_385),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_160),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_214),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_621),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_385),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_60),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_281),
.Y(n_715)
);

CKINVDCx16_ASAP7_75t_R g716 ( 
.A(n_331),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_478),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_343),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_184),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_134),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_74),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_591),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_490),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_475),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_33),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_35),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_275),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_575),
.Y(n_728)
);

BUFx10_ASAP7_75t_L g729 ( 
.A(n_228),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_569),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_527),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_406),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_119),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_13),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_449),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_527),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_578),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_501),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_184),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_520),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_165),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_359),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_231),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_26),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_239),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_151),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_182),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_72),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_525),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_306),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_49),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_219),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_242),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_269),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_74),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_553),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_143),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_327),
.Y(n_758)
);

CKINVDCx14_ASAP7_75t_R g759 ( 
.A(n_266),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_88),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_525),
.Y(n_761)
);

BUFx5_ASAP7_75t_L g762 ( 
.A(n_380),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_172),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_464),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_320),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_307),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_340),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_484),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_308),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_397),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_563),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_211),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_450),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_61),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_446),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_172),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_616),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_561),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_468),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_429),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_375),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_109),
.Y(n_782)
);

BUFx10_ASAP7_75t_L g783 ( 
.A(n_25),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_601),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_436),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_240),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_388),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_442),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_406),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_413),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_549),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_368),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_460),
.Y(n_793)
);

CKINVDCx14_ASAP7_75t_R g794 ( 
.A(n_503),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_26),
.Y(n_795)
);

CKINVDCx16_ASAP7_75t_R g796 ( 
.A(n_391),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_523),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_103),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_539),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_529),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_510),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_528),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_530),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_375),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_450),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_392),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_297),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_404),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_607),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_346),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_402),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_155),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_496),
.Y(n_813)
);

CKINVDCx14_ASAP7_75t_R g814 ( 
.A(n_83),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_175),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_473),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_49),
.Y(n_817)
);

BUFx10_ASAP7_75t_L g818 ( 
.A(n_23),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_276),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_12),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_284),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_474),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_266),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_204),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_108),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_558),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_279),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_55),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_114),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_425),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_147),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_283),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_303),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_511),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_87),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_90),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_535),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_179),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_347),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_623),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_156),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_97),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_236),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_139),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_360),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_458),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_305),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_464),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_149),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_403),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_103),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_47),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_271),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_367),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_330),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_362),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_80),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_518),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_388),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_577),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_259),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_69),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_92),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_417),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_597),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_468),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_96),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_398),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_515),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_547),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_289),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_18),
.Y(n_872)
);

BUFx10_ASAP7_75t_L g873 ( 
.A(n_583),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_503),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_27),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_132),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_502),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_31),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_430),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_222),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_31),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_357),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_324),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_284),
.Y(n_884)
);

INVx4_ASAP7_75t_R g885 ( 
.A(n_550),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_128),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_619),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_498),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_75),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_364),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_155),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_295),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_419),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_109),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_539),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_488),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_133),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_390),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_629),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_55),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_121),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_582),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_352),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_584),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_304),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_296),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_608),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_152),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_427),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_106),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_321),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_614),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_504),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_132),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_563),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_5),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_434),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_502),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_351),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_166),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_461),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_574),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_497),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_179),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_96),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_562),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_107),
.Y(n_927)
);

CKINVDCx14_ASAP7_75t_R g928 ( 
.A(n_264),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_461),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_413),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_192),
.Y(n_931)
);

CKINVDCx16_ASAP7_75t_R g932 ( 
.A(n_508),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_192),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_123),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_217),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_295),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_61),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_357),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_116),
.Y(n_939)
);

CKINVDCx14_ASAP7_75t_R g940 ( 
.A(n_312),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_596),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_520),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_160),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_342),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_221),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_256),
.Y(n_946)
);

CKINVDCx16_ASAP7_75t_R g947 ( 
.A(n_157),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_223),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_207),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_69),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_588),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_602),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_277),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_66),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_626),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_13),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_429),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_129),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_143),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_329),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_500),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_215),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_512),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_581),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_425),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_348),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_631),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_318),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_121),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_334),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_459),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_148),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_110),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_219),
.Y(n_974)
);

CKINVDCx14_ASAP7_75t_R g975 ( 
.A(n_243),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_500),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_529),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_168),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_85),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_27),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_407),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_276),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_370),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_130),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_609),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_414),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_21),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_33),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_146),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_439),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_484),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_68),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_495),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_315),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_421),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_230),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_269),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_627),
.Y(n_998)
);

BUFx10_ASAP7_75t_L g999 ( 
.A(n_85),
.Y(n_999)
);

INVxp33_ASAP7_75t_SL g1000 ( 
.A(n_181),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_471),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_19),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_630),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_56),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_196),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_416),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_153),
.Y(n_1007)
);

BUFx5_ASAP7_75t_L g1008 ( 
.A(n_570),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_611),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_605),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_311),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_350),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_205),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_387),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_105),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_114),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_164),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_506),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_66),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_120),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_410),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_355),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_428),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_532),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_435),
.Y(n_1025)
);

BUFx10_ASAP7_75t_L g1026 ( 
.A(n_272),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_524),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_455),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_300),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_164),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_191),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_180),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_175),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_593),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_368),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_325),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_111),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_552),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_153),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_449),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_441),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_580),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_335),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_221),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_76),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_485),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_393),
.Y(n_1048)
);

CKINVDCx14_ASAP7_75t_R g1049 ( 
.A(n_4),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_439),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_365),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_466),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_567),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_215),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_163),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_247),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_498),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_462),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_912),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_684),
.Y(n_1060)
);

CKINVDCx16_ASAP7_75t_R g1061 ( 
.A(n_653),
.Y(n_1061)
);

INVxp33_ASAP7_75t_L g1062 ( 
.A(n_1048),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_759),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_684),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_684),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_684),
.Y(n_1066)
);

INVxp33_ASAP7_75t_SL g1067 ( 
.A(n_782),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_684),
.Y(n_1068)
);

INVxp67_ASAP7_75t_L g1069 ( 
.A(n_782),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_684),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_794),
.Y(n_1071)
);

INVxp67_ASAP7_75t_SL g1072 ( 
.A(n_777),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_899),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_777),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_814),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_684),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_928),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_684),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_684),
.Y(n_1079)
);

INVxp33_ASAP7_75t_SL g1080 ( 
.A(n_845),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_762),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_940),
.Y(n_1082)
);

INVxp67_ASAP7_75t_SL g1083 ( 
.A(n_717),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_762),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_762),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_762),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_762),
.Y(n_1087)
);

CKINVDCx16_ASAP7_75t_R g1088 ( 
.A(n_653),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_975),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_1049),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_762),
.Y(n_1091)
);

BUFx2_ASAP7_75t_SL g1092 ( 
.A(n_964),
.Y(n_1092)
);

INVxp67_ASAP7_75t_SL g1093 ( 
.A(n_717),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_641),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_762),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_762),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_762),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_717),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_717),
.Y(n_1099)
);

INVxp33_ASAP7_75t_SL g1100 ( 
.A(n_845),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_717),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_722),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_717),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_964),
.B(n_0),
.Y(n_1104)
);

INVxp33_ASAP7_75t_SL g1105 ( 
.A(n_1053),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1051),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_1053),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1051),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1051),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1051),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_728),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1051),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1051),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_694),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_688),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_694),
.Y(n_1116)
);

INVxp33_ASAP7_75t_L g1117 ( 
.A(n_635),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_694),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_694),
.Y(n_1119)
);

INVxp67_ASAP7_75t_SL g1120 ( 
.A(n_694),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_701),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_701),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_701),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_701),
.Y(n_1124)
);

INVxp33_ASAP7_75t_SL g1125 ( 
.A(n_690),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_688),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_730),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_701),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_713),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_704),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_647),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_704),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_647),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_873),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_712),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_716),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_899),
.Y(n_1137)
);

INVxp67_ASAP7_75t_SL g1138 ( 
.A(n_713),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_712),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_737),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_637),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_737),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_951),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_713),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_873),
.Y(n_1145)
);

INVxp33_ASAP7_75t_SL g1146 ( 
.A(n_690),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_951),
.Y(n_1147)
);

INVxp33_ASAP7_75t_SL g1148 ( 
.A(n_632),
.Y(n_1148)
);

INVxp67_ASAP7_75t_SL g1149 ( 
.A(n_713),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_952),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_716),
.Y(n_1151)
);

INVxp67_ASAP7_75t_SL g1152 ( 
.A(n_713),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_952),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1009),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_725),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1009),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_637),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_655),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_635),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_R g1160 ( 
.A(n_1000),
.B(n_0),
.Y(n_1160)
);

INVxp67_ASAP7_75t_SL g1161 ( 
.A(n_725),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_655),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_709),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_709),
.Y(n_1164)
);

INVxp67_ASAP7_75t_SL g1165 ( 
.A(n_725),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_796),
.Y(n_1166)
);

INVxp33_ASAP7_75t_SL g1167 ( 
.A(n_633),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_725),
.Y(n_1168)
);

INVxp67_ASAP7_75t_SL g1169 ( 
.A(n_725),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_770),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_770),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_868),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_868),
.Y(n_1173)
);

INVxp67_ASAP7_75t_SL g1174 ( 
.A(n_735),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_784),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_735),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_796),
.Y(n_1177)
);

INVxp67_ASAP7_75t_SL g1178 ( 
.A(n_735),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_871),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_735),
.Y(n_1180)
);

INVxp33_ASAP7_75t_SL g1181 ( 
.A(n_639),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_871),
.Y(n_1182)
);

CKINVDCx16_ASAP7_75t_R g1183 ( 
.A(n_932),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_893),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_893),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_903),
.Y(n_1186)
);

CKINVDCx16_ASAP7_75t_R g1187 ( 
.A(n_932),
.Y(n_1187)
);

INVxp33_ASAP7_75t_SL g1188 ( 
.A(n_640),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_903),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_873),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_926),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_926),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_947),
.Y(n_1193)
);

BUFx2_ASAP7_75t_SL g1194 ( 
.A(n_638),
.Y(n_1194)
);

INVxp33_ASAP7_75t_L g1195 ( 
.A(n_636),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_735),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_634),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_958),
.Y(n_1198)
);

INVxp33_ASAP7_75t_L g1199 ( 
.A(n_636),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_756),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_756),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_756),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_661),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_756),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_756),
.Y(n_1205)
);

INVxp33_ASAP7_75t_SL g1206 ( 
.A(n_643),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_828),
.Y(n_1207)
);

INVxp33_ASAP7_75t_L g1208 ( 
.A(n_642),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_828),
.Y(n_1209)
);

INVxp67_ASAP7_75t_SL g1210 ( 
.A(n_828),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_958),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_947),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_646),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_828),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_986),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_986),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_828),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_876),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1006),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1006),
.Y(n_1220)
);

INVxp67_ASAP7_75t_SL g1221 ( 
.A(n_876),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1030),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1030),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1037),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_648),
.Y(n_1225)
);

CKINVDCx14_ASAP7_75t_R g1226 ( 
.A(n_687),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_876),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_876),
.Y(n_1228)
);

INVxp67_ASAP7_75t_SL g1229 ( 
.A(n_876),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_886),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_886),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_809),
.Y(n_1232)
);

INVxp67_ASAP7_75t_SL g1233 ( 
.A(n_886),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1037),
.Y(n_1234)
);

INVxp67_ASAP7_75t_SL g1235 ( 
.A(n_886),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_886),
.Y(n_1236)
);

INVxp67_ASAP7_75t_SL g1237 ( 
.A(n_920),
.Y(n_1237)
);

INVxp33_ASAP7_75t_SL g1238 ( 
.A(n_651),
.Y(n_1238)
);

INVxp67_ASAP7_75t_SL g1239 ( 
.A(n_920),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_920),
.Y(n_1240)
);

CKINVDCx16_ASAP7_75t_R g1241 ( 
.A(n_687),
.Y(n_1241)
);

INVxp67_ASAP7_75t_SL g1242 ( 
.A(n_920),
.Y(n_1242)
);

INVxp33_ASAP7_75t_L g1243 ( 
.A(n_642),
.Y(n_1243)
);

INVxp67_ASAP7_75t_SL g1244 ( 
.A(n_920),
.Y(n_1244)
);

INVxp33_ASAP7_75t_L g1245 ( 
.A(n_645),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_943),
.Y(n_1246)
);

INVxp33_ASAP7_75t_SL g1247 ( 
.A(n_658),
.Y(n_1247)
);

INVxp33_ASAP7_75t_L g1248 ( 
.A(n_645),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_943),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_943),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_943),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_943),
.Y(n_1252)
);

CKINVDCx14_ASAP7_75t_R g1253 ( 
.A(n_687),
.Y(n_1253)
);

CKINVDCx14_ASAP7_75t_R g1254 ( 
.A(n_687),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_989),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_840),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_989),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_989),
.Y(n_1258)
);

CKINVDCx16_ASAP7_75t_R g1259 ( 
.A(n_705),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_989),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_989),
.Y(n_1261)
);

CKINVDCx16_ASAP7_75t_R g1262 ( 
.A(n_705),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_682),
.Y(n_1263)
);

INVxp67_ASAP7_75t_SL g1264 ( 
.A(n_697),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_662),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_665),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_644),
.Y(n_1267)
);

INVxp67_ASAP7_75t_SL g1268 ( 
.A(n_697),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_649),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_649),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_650),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_650),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_668),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_669),
.Y(n_1274)
);

INVxp67_ASAP7_75t_SL g1275 ( 
.A(n_674),
.Y(n_1275)
);

CKINVDCx16_ASAP7_75t_R g1276 ( 
.A(n_705),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_652),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_899),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1073),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1116),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1101),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1073),
.Y(n_1282)
);

INVx6_ASAP7_75t_L g1283 ( 
.A(n_1073),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1084),
.A2(n_686),
.B(n_644),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1101),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1157),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1116),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1084),
.A2(n_700),
.B(n_686),
.Y(n_1288)
);

BUFx12f_ASAP7_75t_L g1289 ( 
.A(n_1077),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1072),
.B(n_1043),
.Y(n_1290)
);

XOR2xp5_ASAP7_75t_L g1291 ( 
.A(n_1059),
.B(n_752),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1134),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1118),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1112),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1118),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1067),
.A2(n_670),
.B1(n_672),
.B2(n_671),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1092),
.B(n_860),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1115),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1119),
.Y(n_1299)
);

INVx5_ASAP7_75t_L g1300 ( 
.A(n_1073),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1114),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1073),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1112),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1113),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1113),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1074),
.B(n_638),
.Y(n_1306)
);

BUFx12f_ASAP7_75t_L g1307 ( 
.A(n_1077),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1137),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1137),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1124),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1063),
.Y(n_1311)
);

CKINVDCx14_ASAP7_75t_R g1312 ( 
.A(n_1226),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1124),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1137),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1137),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1119),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1155),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1155),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1121),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1120),
.B(n_1128),
.Y(n_1320)
);

CKINVDCx6p67_ASAP7_75t_R g1321 ( 
.A(n_1071),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1115),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1168),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1168),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1176),
.Y(n_1325)
);

BUFx8_ASAP7_75t_SL g1326 ( 
.A(n_1075),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1121),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1094),
.Y(n_1328)
);

INVx5_ASAP7_75t_L g1329 ( 
.A(n_1176),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1180),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1180),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1196),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1060),
.A2(n_749),
.B(n_700),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1194),
.B(n_766),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1196),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1200),
.Y(n_1336)
);

CKINVDCx11_ASAP7_75t_R g1337 ( 
.A(n_1089),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1158),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1098),
.A2(n_1055),
.B(n_654),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1098),
.A2(n_1103),
.B(n_1099),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1122),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1162),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1092),
.B(n_865),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1122),
.Y(n_1344)
);

BUFx8_ASAP7_75t_L g1345 ( 
.A(n_1266),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1138),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1200),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1144),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1149),
.B(n_899),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1227),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1067),
.A2(n_677),
.B1(n_678),
.B2(n_675),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1227),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1080),
.A2(n_680),
.B1(n_683),
.B2(n_679),
.Y(n_1353)
);

AOI22xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1080),
.A2(n_773),
.B1(n_793),
.B2(n_772),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1228),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1228),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1230),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_1230),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1123),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1148),
.B(n_887),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1100),
.A2(n_689),
.B1(n_691),
.B2(n_685),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1064),
.A2(n_771),
.B(n_749),
.Y(n_1362)
);

CKINVDCx16_ASAP7_75t_R g1363 ( 
.A(n_1061),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1123),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1100),
.A2(n_695),
.B1(n_696),
.B2(n_693),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1231),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1129),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1194),
.B(n_766),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1152),
.B(n_899),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1130),
.Y(n_1370)
);

CKINVDCx8_ASAP7_75t_R g1371 ( 
.A(n_1088),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1231),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1099),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1129),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1161),
.B(n_902),
.Y(n_1375)
);

OAI21xp33_ASAP7_75t_L g1376 ( 
.A1(n_1105),
.A2(n_812),
.B(n_780),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1163),
.B(n_780),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1103),
.Y(n_1378)
);

INVx5_ASAP7_75t_L g1379 ( 
.A(n_1134),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1201),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1165),
.B(n_1003),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_1201),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1169),
.B(n_904),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1164),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1106),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1106),
.A2(n_1109),
.B(n_1108),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1170),
.Y(n_1387)
);

INVxp33_ASAP7_75t_SL g1388 ( 
.A(n_1082),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1108),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1202),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1174),
.B(n_1178),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1210),
.B(n_1003),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1221),
.B(n_1003),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1229),
.B(n_1003),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1233),
.B(n_907),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1102),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1148),
.B(n_922),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1109),
.A2(n_1046),
.B(n_1045),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1110),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1171),
.B(n_812),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1110),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1126),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1202),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1126),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1172),
.Y(n_1405)
);

NOR2x1_ASAP7_75t_L g1406 ( 
.A(n_1145),
.B(n_1003),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1132),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1173),
.B(n_852),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1204),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1235),
.B(n_941),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1105),
.A2(n_703),
.B1(n_706),
.B2(n_702),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1204),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1205),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1205),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1207),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1179),
.B(n_852),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1207),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1132),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1209),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1209),
.Y(n_1420)
);

BUFx12f_ASAP7_75t_L g1421 ( 
.A(n_1082),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1214),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1214),
.Y(n_1423)
);

INVx4_ASAP7_75t_L g1424 ( 
.A(n_1145),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1076),
.A2(n_1055),
.B(n_654),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1217),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1217),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1218),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1218),
.Y(n_1429)
);

AND2x6_ASAP7_75t_L g1430 ( 
.A(n_1076),
.B(n_985),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1237),
.B(n_955),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1239),
.B(n_967),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1136),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1182),
.B(n_874),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1242),
.B(n_998),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1244),
.B(n_985),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1136),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1250),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1250),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1252),
.Y(n_1440)
);

XNOR2xp5_ASAP7_75t_L g1441 ( 
.A(n_1197),
.B(n_806),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1310),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1310),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1313),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1286),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1320),
.B(n_1249),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1313),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1286),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1320),
.B(n_1083),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1279),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1317),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1317),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1338),
.Y(n_1453)
);

BUFx8_ASAP7_75t_L g1454 ( 
.A(n_1289),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1279),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1292),
.B(n_1090),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1318),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1338),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1342),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1342),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1384),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1384),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1292),
.B(n_1090),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1320),
.B(n_1093),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1441),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1387),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1387),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1405),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1318),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1284),
.A2(n_1066),
.B(n_1065),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1405),
.Y(n_1471)
);

AND2x6_ASAP7_75t_L g1472 ( 
.A(n_1334),
.B(n_985),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1441),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1279),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1333),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1391),
.B(n_1278),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1279),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1333),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1279),
.Y(n_1479)
);

NOR2x1_ASAP7_75t_L g1480 ( 
.A(n_1424),
.B(n_1111),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1362),
.Y(n_1481)
);

CKINVDCx16_ASAP7_75t_R g1482 ( 
.A(n_1363),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1362),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1282),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1370),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1323),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1284),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1288),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1323),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1375),
.B(n_1264),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1324),
.Y(n_1491)
);

AND2x6_ASAP7_75t_L g1492 ( 
.A(n_1334),
.B(n_985),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1322),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1368),
.B(n_1131),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1288),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1383),
.B(n_1395),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1425),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1368),
.B(n_1133),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1410),
.B(n_1268),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1425),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1425),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1431),
.B(n_1236),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1349),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1282),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1282),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1322),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1425),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1324),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1282),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1280),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1306),
.B(n_1135),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1331),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1331),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1280),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1287),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1287),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1293),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1293),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1306),
.B(n_1139),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1282),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1340),
.A2(n_1070),
.B(n_1068),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1432),
.B(n_1240),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1435),
.B(n_1246),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1290),
.B(n_1167),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1301),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1346),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1332),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1332),
.Y(n_1528)
);

OA21x2_ASAP7_75t_L g1529 ( 
.A1(n_1295),
.A2(n_1079),
.B(n_1078),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1348),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1302),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1295),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1335),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1299),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1335),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1336),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1377),
.B(n_1140),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1336),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1360),
.B(n_1241),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1299),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1297),
.B(n_1167),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1406),
.B(n_1142),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1402),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1316),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1316),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1355),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1302),
.Y(n_1547)
);

INVx4_ASAP7_75t_L g1548 ( 
.A(n_1380),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1319),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1355),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1402),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1343),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1319),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1377),
.B(n_1143),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1366),
.Y(n_1555)
);

AND2x6_ASAP7_75t_L g1556 ( 
.A(n_1436),
.B(n_985),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1366),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1281),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1327),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1281),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1327),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1341),
.Y(n_1562)
);

AND2x6_ASAP7_75t_L g1563 ( 
.A(n_1436),
.B(n_985),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1302),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1285),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1397),
.B(n_1276),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1349),
.B(n_1251),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1349),
.B(n_1147),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1302),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1341),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1407),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1344),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1344),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1285),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1359),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1298),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1359),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1364),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1364),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1367),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1367),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1374),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1374),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1380),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1390),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1390),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1294),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1409),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1302),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1409),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1412),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1309),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1412),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1311),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1420),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1309),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1420),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1309),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1309),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1369),
.B(n_1252),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1294),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1423),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1303),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1400),
.B(n_1150),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1423),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1428),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1428),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_L g1608 ( 
.A(n_1309),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1378),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1369),
.B(n_1153),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1303),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1304),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1378),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1314),
.Y(n_1614)
);

BUFx8_ASAP7_75t_L g1615 ( 
.A(n_1289),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1314),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1378),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1401),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1304),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1314),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1314),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1401),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1401),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1369),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1407),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1440),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1291),
.A2(n_842),
.B1(n_853),
.B2(n_830),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1418),
.Y(n_1628)
);

INVxp67_ASAP7_75t_L g1629 ( 
.A(n_1418),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1381),
.B(n_1154),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1314),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1381),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_L g1633 ( 
.A(n_1315),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1381),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1315),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1305),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1392),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1291),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1305),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1403),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1392),
.B(n_1393),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1373),
.A2(n_1389),
.B(n_1385),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1392),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1403),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1393),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1393),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1379),
.B(n_1259),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_L g1648 ( 
.A(n_1315),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1394),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1379),
.B(n_1262),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1394),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1315),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1394),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1404),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1440),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1440),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1436),
.B(n_1156),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1414),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1339),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1414),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1417),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1339),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1339),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1379),
.B(n_1181),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1339),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1417),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1398),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1398),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1398),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1433),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1379),
.B(n_1181),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1380),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1419),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1379),
.B(n_1255),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1380),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_1315),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_SL g1677 ( 
.A(n_1424),
.B(n_1188),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1400),
.B(n_1184),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1380),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1382),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1419),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1300),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1427),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1424),
.B(n_1188),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1326),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1308),
.B(n_1255),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1388),
.B(n_1206),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1427),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1552),
.B(n_1125),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1541),
.B(n_1125),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1503),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1503),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1642),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1641),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1624),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1685),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1641),
.B(n_1398),
.Y(n_1697)
);

AND2x6_ASAP7_75t_L g1698 ( 
.A(n_1497),
.B(n_1408),
.Y(n_1698)
);

INVxp67_ASAP7_75t_SL g1699 ( 
.A(n_1641),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1632),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1678),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1642),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1496),
.B(n_1388),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1524),
.B(n_1146),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1445),
.B(n_1408),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_1529),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1634),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1637),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1490),
.B(n_1146),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1643),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1645),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1657),
.Y(n_1712)
);

INVx3_ASAP7_75t_L g1713 ( 
.A(n_1657),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1642),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1657),
.B(n_1433),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1568),
.B(n_1437),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1529),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1568),
.Y(n_1718)
);

AND2x6_ASAP7_75t_L g1719 ( 
.A(n_1497),
.B(n_1416),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1499),
.B(n_1525),
.Y(n_1720)
);

BUFx6f_ASAP7_75t_L g1721 ( 
.A(n_1529),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1485),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1646),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1442),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_1477),
.Y(n_1725)
);

OA22x2_ASAP7_75t_L g1726 ( 
.A1(n_1678),
.A2(n_1376),
.B1(n_1069),
.B2(n_1107),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1649),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1651),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1653),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1510),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1477),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1449),
.B(n_1253),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1442),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1526),
.B(n_1206),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1500),
.A2(n_1104),
.B1(n_776),
.B2(n_866),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1443),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1443),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1568),
.B(n_1437),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1448),
.Y(n_1739)
);

INVxp67_ASAP7_75t_L g1740 ( 
.A(n_1485),
.Y(n_1740)
);

INVx4_ASAP7_75t_SL g1741 ( 
.A(n_1556),
.Y(n_1741)
);

INVx4_ASAP7_75t_L g1742 ( 
.A(n_1610),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1610),
.B(n_1371),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1610),
.B(n_1371),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1464),
.B(n_1254),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1630),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1530),
.B(n_1238),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1510),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1630),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1446),
.B(n_1213),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1514),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1453),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1638),
.B(n_1203),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1476),
.B(n_1213),
.Y(n_1754)
);

INVx4_ASAP7_75t_L g1755 ( 
.A(n_1630),
.Y(n_1755)
);

BUFx10_ASAP7_75t_L g1756 ( 
.A(n_1685),
.Y(n_1756)
);

XOR2xp5_ASAP7_75t_L g1757 ( 
.A(n_1482),
.B(n_1328),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1444),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1444),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1514),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1477),
.Y(n_1761)
);

NOR2x1p5_ASAP7_75t_L g1762 ( 
.A(n_1458),
.B(n_1421),
.Y(n_1762)
);

BUFx3_ASAP7_75t_L g1763 ( 
.A(n_1459),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_1493),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1502),
.B(n_1274),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1447),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1594),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1500),
.B(n_1183),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1447),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1539),
.B(n_1238),
.Y(n_1770)
);

INVx3_ASAP7_75t_L g1771 ( 
.A(n_1451),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1501),
.B(n_1187),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1451),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1515),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1452),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1515),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1516),
.Y(n_1777)
);

AND2x6_ASAP7_75t_L g1778 ( 
.A(n_1501),
.B(n_1416),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1516),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1566),
.B(n_1247),
.Y(n_1780)
);

INVx2_ASAP7_75t_SL g1781 ( 
.A(n_1537),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1507),
.A2(n_1175),
.B1(n_1232),
.B2(n_1127),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1522),
.B(n_1274),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1537),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1477),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1594),
.Y(n_1786)
);

BUFx10_ASAP7_75t_L g1787 ( 
.A(n_1465),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1517),
.Y(n_1788)
);

BUFx10_ASAP7_75t_L g1789 ( 
.A(n_1542),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1517),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1518),
.Y(n_1791)
);

BUFx3_ASAP7_75t_L g1792 ( 
.A(n_1460),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1452),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1493),
.B(n_1263),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1518),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1507),
.B(n_1008),
.Y(n_1796)
);

BUFx6f_ASAP7_75t_L g1797 ( 
.A(n_1477),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1593),
.Y(n_1798)
);

BUFx4f_ASAP7_75t_L g1799 ( 
.A(n_1506),
.Y(n_1799)
);

INVx4_ASAP7_75t_L g1800 ( 
.A(n_1479),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1457),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1659),
.A2(n_776),
.B1(n_866),
.B2(n_771),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1542),
.B(n_1008),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1523),
.B(n_1340),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_SL g1805 ( 
.A(n_1454),
.B(n_1307),
.Y(n_1805)
);

OR2x6_ASAP7_75t_L g1806 ( 
.A(n_1506),
.B(n_1307),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1593),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1554),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1479),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1457),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1494),
.B(n_1247),
.Y(n_1811)
);

BUFx4f_ASAP7_75t_L g1812 ( 
.A(n_1543),
.Y(n_1812)
);

INVx4_ASAP7_75t_L g1813 ( 
.A(n_1479),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1494),
.B(n_1498),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1498),
.B(n_1256),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1605),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1511),
.B(n_1312),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1542),
.B(n_1008),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1461),
.B(n_1351),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1543),
.B(n_1177),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1605),
.Y(n_1821)
);

INVx4_ASAP7_75t_L g1822 ( 
.A(n_1479),
.Y(n_1822)
);

BUFx3_ASAP7_75t_L g1823 ( 
.A(n_1462),
.Y(n_1823)
);

INVx3_ASAP7_75t_L g1824 ( 
.A(n_1469),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1659),
.B(n_1008),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1662),
.A2(n_890),
.B1(n_935),
.B2(n_900),
.Y(n_1826)
);

INVx3_ASAP7_75t_L g1827 ( 
.A(n_1469),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1606),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1486),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1606),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1486),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1607),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1466),
.B(n_1467),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1489),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1454),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1607),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1479),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1489),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1511),
.B(n_1340),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1491),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1491),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1626),
.Y(n_1842)
);

AND2x6_ASAP7_75t_L g1843 ( 
.A(n_1662),
.B(n_1434),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1663),
.A2(n_890),
.B1(n_935),
.B2(n_900),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1626),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_SL g1846 ( 
.A(n_1454),
.B(n_1421),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1519),
.B(n_1554),
.Y(n_1847)
);

INVx2_ASAP7_75t_SL g1848 ( 
.A(n_1604),
.Y(n_1848)
);

INVx4_ASAP7_75t_L g1849 ( 
.A(n_1484),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1609),
.Y(n_1850)
);

BUFx3_ASAP7_75t_L g1851 ( 
.A(n_1468),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1508),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1551),
.B(n_1212),
.Y(n_1853)
);

NAND2xp33_ASAP7_75t_L g1854 ( 
.A(n_1663),
.B(n_1008),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1609),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1613),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1613),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1519),
.A2(n_1667),
.B1(n_1668),
.B2(n_1665),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1623),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1508),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1623),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_1471),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1532),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1604),
.B(n_1225),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1512),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_SL g1866 ( 
.A(n_1615),
.B(n_1328),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1665),
.A2(n_978),
.B1(n_897),
.B2(n_945),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1512),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1677),
.A2(n_1166),
.B1(n_1193),
.B2(n_1151),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1534),
.B(n_1434),
.Y(n_1870)
);

INVxp67_ASAP7_75t_SL g1871 ( 
.A(n_1600),
.Y(n_1871)
);

INVx5_ASAP7_75t_L g1872 ( 
.A(n_1556),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1540),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1513),
.Y(n_1874)
);

OAI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1629),
.A2(n_1160),
.B1(n_1062),
.B2(n_1117),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1551),
.B(n_1265),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_SL g1877 ( 
.A(n_1667),
.B(n_1008),
.Y(n_1877)
);

BUFx10_ASAP7_75t_L g1878 ( 
.A(n_1473),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1513),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1571),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1668),
.B(n_1008),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1544),
.Y(n_1882)
);

INVx4_ASAP7_75t_L g1883 ( 
.A(n_1484),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1669),
.B(n_1008),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1545),
.Y(n_1885)
);

INVx4_ASAP7_75t_L g1886 ( 
.A(n_1484),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1669),
.B(n_1617),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1549),
.Y(n_1888)
);

INVx2_ASAP7_75t_SL g1889 ( 
.A(n_1670),
.Y(n_1889)
);

NAND2xp33_ASAP7_75t_SL g1890 ( 
.A(n_1571),
.B(n_867),
.Y(n_1890)
);

HB1xp67_ASAP7_75t_L g1891 ( 
.A(n_1625),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1553),
.Y(n_1892)
);

NOR3xp33_ASAP7_75t_L g1893 ( 
.A(n_1627),
.B(n_1353),
.C(n_1296),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1618),
.B(n_1008),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1559),
.Y(n_1895)
);

INVx4_ASAP7_75t_L g1896 ( 
.A(n_1484),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1625),
.B(n_1273),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1475),
.A2(n_978),
.B1(n_897),
.B2(n_945),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1622),
.B(n_1365),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1628),
.B(n_1266),
.Y(n_1900)
);

BUFx2_ASAP7_75t_L g1901 ( 
.A(n_1628),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1561),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1527),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1576),
.B(n_1151),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1527),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1562),
.B(n_1340),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1528),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1655),
.B(n_1656),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1570),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1567),
.B(n_1411),
.Y(n_1910)
);

AOI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1684),
.A2(n_1193),
.B1(n_1166),
.B2(n_1035),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1572),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1573),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1654),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1575),
.Y(n_1915)
);

CKINVDCx20_ASAP7_75t_R g1916 ( 
.A(n_1615),
.Y(n_1916)
);

BUFx3_ASAP7_75t_L g1917 ( 
.A(n_1577),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1578),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1528),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1579),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1580),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1475),
.B(n_1010),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1581),
.B(n_1386),
.Y(n_1923)
);

AND2x2_ASAP7_75t_SL g1924 ( 
.A(n_1478),
.B(n_652),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1582),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1533),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1583),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1585),
.B(n_1386),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1533),
.Y(n_1929)
);

AND2x6_ASAP7_75t_SL g1930 ( 
.A(n_1615),
.B(n_656),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1586),
.B(n_1386),
.Y(n_1931)
);

INVxp67_ASAP7_75t_L g1932 ( 
.A(n_1456),
.Y(n_1932)
);

INVx1_ASAP7_75t_SL g1933 ( 
.A(n_1687),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1588),
.B(n_1590),
.Y(n_1934)
);

BUFx3_ASAP7_75t_L g1935 ( 
.A(n_1591),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1480),
.B(n_1190),
.Y(n_1936)
);

INVx4_ASAP7_75t_SL g1937 ( 
.A(n_1556),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1595),
.B(n_1386),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_1463),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1597),
.B(n_1413),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1535),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1602),
.B(n_1647),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1535),
.Y(n_1943)
);

INVx3_ASAP7_75t_L g1944 ( 
.A(n_1536),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1650),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_L g1946 ( 
.A1(n_1478),
.A2(n_1019),
.B1(n_1032),
.B2(n_874),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1664),
.B(n_1190),
.Y(n_1947)
);

INVx2_ASAP7_75t_SL g1948 ( 
.A(n_1671),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1672),
.B(n_1361),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1487),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1675),
.B(n_1275),
.Y(n_1951)
);

OR2x6_ASAP7_75t_L g1952 ( 
.A(n_1481),
.B(n_1141),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1536),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1481),
.B(n_1396),
.Y(n_1954)
);

INVx6_ASAP7_75t_L g1955 ( 
.A(n_1548),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1487),
.Y(n_1956)
);

INVx4_ASAP7_75t_SL g1957 ( 
.A(n_1556),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1691),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1707),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1720),
.B(n_1521),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1720),
.B(n_1709),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1707),
.Y(n_1962)
);

NAND3xp33_ASAP7_75t_L g1963 ( 
.A(n_1704),
.B(n_1345),
.C(n_1354),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1814),
.B(n_1521),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1847),
.B(n_1396),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1704),
.A2(n_1472),
.B1(n_1492),
.B2(n_1556),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1814),
.B(n_1483),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1710),
.Y(n_1968)
);

NOR3xp33_ASAP7_75t_L g1969 ( 
.A(n_1690),
.B(n_1337),
.C(n_1141),
.Y(n_1969)
);

AOI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1690),
.A2(n_1492),
.B1(n_1472),
.B2(n_1556),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1696),
.Y(n_1971)
);

INVxp67_ASAP7_75t_L g1972 ( 
.A(n_1794),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1710),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1694),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1839),
.B(n_1483),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1724),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1724),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1709),
.B(n_1693),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1694),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1802),
.A2(n_1495),
.B1(n_1488),
.B2(n_657),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1842),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1693),
.B(n_1488),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1845),
.Y(n_1983)
);

NAND3xp33_ASAP7_75t_SL g1984 ( 
.A(n_1893),
.B(n_1311),
.C(n_930),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1733),
.Y(n_1985)
);

BUFx2_ASAP7_75t_L g1986 ( 
.A(n_1901),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1742),
.B(n_1746),
.Y(n_1987)
);

BUFx5_ASAP7_75t_L g1988 ( 
.A(n_1698),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1864),
.B(n_1321),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1850),
.Y(n_1990)
);

BUFx6f_ASAP7_75t_L g1991 ( 
.A(n_1691),
.Y(n_1991)
);

OAI22x1_ASAP7_75t_SL g1992 ( 
.A1(n_1767),
.A2(n_944),
.B1(n_946),
.B2(n_875),
.Y(n_1992)
);

AOI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1699),
.A2(n_1492),
.B1(n_1472),
.B2(n_1563),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_L g1994 ( 
.A(n_1703),
.B(n_1321),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1924),
.A2(n_1472),
.B1(n_1492),
.B2(n_1563),
.Y(n_1995)
);

INVx2_ASAP7_75t_SL g1996 ( 
.A(n_1880),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1855),
.Y(n_1997)
);

INVx8_ASAP7_75t_L g1998 ( 
.A(n_1698),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1856),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1871),
.B(n_1472),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1811),
.B(n_1195),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_SL g2002 ( 
.A(n_1742),
.B(n_1345),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1754),
.B(n_1472),
.Y(n_2003)
);

OR2x2_ASAP7_75t_SL g2004 ( 
.A(n_1753),
.B(n_1345),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1880),
.Y(n_2005)
);

AOI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1703),
.A2(n_1492),
.B1(n_1563),
.B2(n_1679),
.Y(n_2006)
);

OAI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1750),
.A2(n_1495),
.B1(n_1208),
.B2(n_1243),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_SL g2008 ( 
.A(n_1722),
.B(n_948),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1857),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1859),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1746),
.B(n_1676),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1730),
.B(n_1492),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1733),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1755),
.B(n_1676),
.Y(n_2014)
);

OAI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1781),
.A2(n_1245),
.B1(n_1248),
.B2(n_1199),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1748),
.B(n_1563),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1751),
.B(n_1563),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1820),
.B(n_1185),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1736),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1755),
.B(n_1484),
.Y(n_2020)
);

OR2x6_ASAP7_75t_L g2021 ( 
.A(n_1806),
.B(n_1019),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_1789),
.B(n_1504),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1811),
.B(n_1186),
.Y(n_2023)
);

A2O1A1Ixp33_ASAP7_75t_L g2024 ( 
.A1(n_1942),
.A2(n_1470),
.B(n_1644),
.C(n_1640),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1861),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1760),
.B(n_1563),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1695),
.Y(n_2027)
);

XOR2xp5_ASAP7_75t_L g2028 ( 
.A(n_1757),
.B(n_994),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1774),
.B(n_1680),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1776),
.B(n_1450),
.Y(n_2030)
);

BUFx6f_ASAP7_75t_L g2031 ( 
.A(n_1691),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1736),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1789),
.B(n_1652),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1777),
.B(n_1450),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_1891),
.Y(n_2035)
);

BUFx3_ASAP7_75t_L g2036 ( 
.A(n_1799),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1689),
.B(n_1002),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1779),
.B(n_1450),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1700),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1788),
.B(n_1455),
.Y(n_2040)
);

OR2x6_ASAP7_75t_L g2041 ( 
.A(n_1806),
.B(n_1889),
.Y(n_2041)
);

NAND2xp33_ASAP7_75t_L g2042 ( 
.A(n_1698),
.B(n_1676),
.Y(n_2042)
);

NOR2xp67_ASAP7_75t_L g2043 ( 
.A(n_1740),
.B(n_1159),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1789),
.B(n_1676),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1708),
.Y(n_2045)
);

INVxp67_ASAP7_75t_L g2046 ( 
.A(n_1876),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1900),
.B(n_1189),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1711),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1897),
.B(n_1191),
.Y(n_2049)
);

INVx1_ASAP7_75t_SL g2050 ( 
.A(n_1764),
.Y(n_2050)
);

NAND2xp33_ASAP7_75t_L g2051 ( 
.A(n_1698),
.B(n_1676),
.Y(n_2051)
);

AOI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1819),
.A2(n_1584),
.B1(n_1548),
.B2(n_1455),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1790),
.B(n_1455),
.Y(n_2053)
);

NAND2xp33_ASAP7_75t_L g2054 ( 
.A(n_1698),
.B(n_1504),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1791),
.B(n_1795),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1798),
.B(n_1474),
.Y(n_2056)
);

OAI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_1717),
.A2(n_1470),
.B(n_1640),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1807),
.B(n_1474),
.Y(n_2058)
);

OR2x2_ASAP7_75t_L g2059 ( 
.A(n_1853),
.B(n_1192),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1691),
.B(n_1504),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1816),
.B(n_1821),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1689),
.B(n_1013),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1723),
.Y(n_2063)
);

NOR2xp33_ASAP7_75t_L g2064 ( 
.A(n_1782),
.B(n_1021),
.Y(n_2064)
);

INVx3_ASAP7_75t_L g2065 ( 
.A(n_1712),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_1712),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1727),
.Y(n_2067)
);

OAI22xp33_ASAP7_75t_L g2068 ( 
.A1(n_1784),
.A2(n_1052),
.B1(n_1056),
.B2(n_1039),
.Y(n_2068)
);

INVxp67_ASAP7_75t_SL g2069 ( 
.A(n_1702),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1737),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_1765),
.B(n_659),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1728),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_1819),
.A2(n_1584),
.B1(n_1548),
.B2(n_1474),
.Y(n_2073)
);

AOI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_1924),
.A2(n_1778),
.B1(n_1843),
.B2(n_1719),
.Y(n_2074)
);

AOI22xp33_ASAP7_75t_L g2075 ( 
.A1(n_1719),
.A2(n_1658),
.B1(n_1660),
.B2(n_1644),
.Y(n_2075)
);

BUFx3_ASAP7_75t_L g2076 ( 
.A(n_1799),
.Y(n_2076)
);

OAI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_1802),
.A2(n_657),
.B1(n_663),
.B2(n_656),
.Y(n_2077)
);

AND2x4_ASAP7_75t_L g2078 ( 
.A(n_1808),
.B(n_1269),
.Y(n_2078)
);

NOR2xp33_ASAP7_75t_L g2079 ( 
.A(n_1783),
.B(n_660),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1702),
.B(n_1681),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_1718),
.B(n_1504),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1714),
.B(n_1681),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1718),
.B(n_1504),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1714),
.B(n_1683),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1737),
.Y(n_2085)
);

INVxp67_ASAP7_75t_L g2086 ( 
.A(n_1891),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_1848),
.B(n_1271),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1729),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1759),
.Y(n_2089)
);

AOI221xp5_ASAP7_75t_L g2090 ( 
.A1(n_1875),
.A2(n_666),
.B1(n_733),
.B2(n_726),
.C(n_673),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1828),
.B(n_1505),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1759),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1713),
.Y(n_2093)
);

OAI21xp33_ASAP7_75t_L g2094 ( 
.A1(n_1734),
.A2(n_791),
.B(n_786),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1858),
.B(n_1830),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1832),
.B(n_1658),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1836),
.B(n_1660),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1713),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1826),
.B(n_1661),
.Y(n_2099)
);

NAND3xp33_ASAP7_75t_L g2100 ( 
.A(n_1734),
.B(n_715),
.C(n_710),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1826),
.B(n_1661),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1844),
.B(n_1666),
.Y(n_2102)
);

INVx4_ASAP7_75t_L g2103 ( 
.A(n_1749),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1749),
.B(n_1652),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1692),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_1815),
.B(n_1652),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1844),
.B(n_1666),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1863),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1906),
.B(n_1923),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_1917),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1928),
.B(n_1673),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1931),
.B(n_1673),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1766),
.Y(n_2113)
);

INVxp67_ASAP7_75t_L g2114 ( 
.A(n_1747),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1873),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1938),
.B(n_1683),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1766),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1882),
.B(n_1505),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1885),
.B(n_1505),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1888),
.B(n_1509),
.Y(n_2120)
);

NAND2xp33_ASAP7_75t_L g2121 ( 
.A(n_1719),
.B(n_1531),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1892),
.Y(n_2122)
);

OAI22xp5_ASAP7_75t_L g2123 ( 
.A1(n_1735),
.A2(n_664),
.B1(n_667),
.B2(n_663),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1895),
.B(n_1509),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1902),
.B(n_1909),
.Y(n_2125)
);

BUFx12f_ASAP7_75t_SL g2126 ( 
.A(n_1806),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_L g2127 ( 
.A(n_1815),
.B(n_870),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_1914),
.B(n_905),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1912),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1913),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1769),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1915),
.B(n_1509),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_1732),
.B(n_1531),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1769),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_1932),
.B(n_934),
.Y(n_2135)
);

NAND3xp33_ASAP7_75t_L g2136 ( 
.A(n_1747),
.B(n_719),
.C(n_718),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1773),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_1917),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1918),
.B(n_1520),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1920),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1921),
.Y(n_2141)
);

NOR3xp33_ASAP7_75t_L g2142 ( 
.A(n_1743),
.B(n_1211),
.C(n_1198),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1925),
.B(n_1927),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_1952),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_1935),
.Y(n_2145)
);

AND2x6_ASAP7_75t_L g2146 ( 
.A(n_1717),
.B(n_1688),
.Y(n_2146)
);

O2A1O1Ixp33_ASAP7_75t_L g2147 ( 
.A1(n_1768),
.A2(n_1032),
.B(n_1686),
.C(n_1688),
.Y(n_2147)
);

INVxp67_ASAP7_75t_L g2148 ( 
.A(n_1904),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1773),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1775),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1934),
.B(n_1520),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_SL g2152 ( 
.A(n_1756),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_SL g2153 ( 
.A(n_1745),
.B(n_1633),
.Y(n_2153)
);

AOI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_1942),
.A2(n_1910),
.B1(n_1922),
.B2(n_1772),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1775),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1793),
.Y(n_2156)
);

NAND2xp33_ASAP7_75t_L g2157 ( 
.A(n_1719),
.B(n_1633),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_1701),
.B(n_1633),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1951),
.B(n_1520),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_1954),
.B(n_1215),
.Y(n_2160)
);

AOI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_1910),
.A2(n_1584),
.B1(n_1599),
.B2(n_1547),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1951),
.B(n_1547),
.Y(n_2162)
);

OR2x2_ASAP7_75t_L g2163 ( 
.A(n_1933),
.B(n_1216),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_1770),
.B(n_960),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1793),
.Y(n_2165)
);

OR2x6_ASAP7_75t_L g2166 ( 
.A(n_1952),
.B(n_1219),
.Y(n_2166)
);

NOR2xp67_ASAP7_75t_L g2167 ( 
.A(n_1945),
.B(n_1270),
.Y(n_2167)
);

INVxp67_ASAP7_75t_L g2168 ( 
.A(n_1817),
.Y(n_2168)
);

OAI22xp33_ASAP7_75t_L g2169 ( 
.A1(n_1939),
.A2(n_1935),
.B1(n_1948),
.B2(n_1952),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1870),
.B(n_1949),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_1812),
.B(n_1531),
.Y(n_2171)
);

BUFx8_ASAP7_75t_L g2172 ( 
.A(n_1936),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1870),
.B(n_1547),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_SL g2174 ( 
.A(n_1812),
.B(n_1531),
.Y(n_2174)
);

BUFx6f_ASAP7_75t_SL g2175 ( 
.A(n_1756),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1870),
.B(n_1599),
.Y(n_2176)
);

INVx2_ASAP7_75t_SL g2177 ( 
.A(n_1833),
.Y(n_2177)
);

INVxp67_ASAP7_75t_L g2178 ( 
.A(n_1890),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1949),
.B(n_1599),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_1770),
.B(n_1220),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_1735),
.B(n_1614),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1801),
.Y(n_2182)
);

BUFx6f_ASAP7_75t_L g2183 ( 
.A(n_1725),
.Y(n_2183)
);

NAND3xp33_ASAP7_75t_L g2184 ( 
.A(n_1768),
.B(n_724),
.C(n_720),
.Y(n_2184)
);

BUFx6f_ASAP7_75t_L g2185 ( 
.A(n_1725),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_L g2186 ( 
.A(n_1780),
.B(n_1024),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1719),
.B(n_1614),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1778),
.B(n_1614),
.Y(n_2188)
);

A2O1A1Ixp33_ASAP7_75t_L g2189 ( 
.A1(n_1780),
.A2(n_1079),
.B(n_1081),
.C(n_1078),
.Y(n_2189)
);

NAND2xp33_ASAP7_75t_L g2190 ( 
.A(n_1778),
.B(n_1633),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_SL g2191 ( 
.A(n_1872),
.B(n_1633),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_1872),
.B(n_1648),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_1947),
.B(n_1715),
.Y(n_2193)
);

OAI22xp5_ASAP7_75t_SL g2194 ( 
.A1(n_1786),
.A2(n_1027),
.B1(n_1025),
.B2(n_754),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1706),
.B(n_1721),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1706),
.B(n_1558),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1801),
.Y(n_2197)
);

INVx8_ASAP7_75t_L g2198 ( 
.A(n_1778),
.Y(n_2198)
);

NAND2x1p5_ASAP7_75t_L g2199 ( 
.A(n_1872),
.B(n_1616),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1706),
.B(n_1558),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_1872),
.B(n_1652),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1706),
.B(n_1560),
.Y(n_2202)
);

NOR2xp67_ASAP7_75t_L g2203 ( 
.A(n_1911),
.B(n_1277),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1721),
.B(n_1560),
.Y(n_2204)
);

INVxp67_ASAP7_75t_L g2205 ( 
.A(n_1890),
.Y(n_2205)
);

INVxp67_ASAP7_75t_L g2206 ( 
.A(n_1716),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1810),
.Y(n_2207)
);

INVx3_ASAP7_75t_L g2208 ( 
.A(n_1833),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_1875),
.B(n_1531),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_1772),
.B(n_734),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1721),
.B(n_1565),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1810),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_1739),
.B(n_1608),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1721),
.B(n_1565),
.Y(n_2214)
);

NAND2xp33_ASAP7_75t_L g2215 ( 
.A(n_1778),
.B(n_1621),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1950),
.B(n_1574),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_SL g2217 ( 
.A(n_1739),
.B(n_1621),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1829),
.Y(n_2218)
);

INVxp33_ASAP7_75t_L g2219 ( 
.A(n_1716),
.Y(n_2219)
);

OAI22xp33_ASAP7_75t_L g2220 ( 
.A1(n_1726),
.A2(n_667),
.B1(n_676),
.B2(n_664),
.Y(n_2220)
);

NAND2xp33_ASAP7_75t_L g2221 ( 
.A(n_1843),
.B(n_1621),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1829),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1956),
.B(n_1574),
.Y(n_2223)
);

INVx1_ASAP7_75t_SL g2224 ( 
.A(n_2050),
.Y(n_2224)
);

OAI22xp5_ASAP7_75t_SL g2225 ( 
.A1(n_2028),
.A2(n_1916),
.B1(n_1835),
.B2(n_1869),
.Y(n_2225)
);

AOI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_2109),
.A2(n_1697),
.B(n_1800),
.Y(n_2226)
);

CKINVDCx5p33_ASAP7_75t_R g2227 ( 
.A(n_1971),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2027),
.Y(n_2228)
);

BUFx6f_ASAP7_75t_L g2229 ( 
.A(n_1958),
.Y(n_2229)
);

BUFx6f_ASAP7_75t_L g2230 ( 
.A(n_1958),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_1958),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_SL g2232 ( 
.A(n_1961),
.B(n_1715),
.Y(n_2232)
);

INVx3_ASAP7_75t_L g2233 ( 
.A(n_2103),
.Y(n_2233)
);

OR2x6_ASAP7_75t_L g2234 ( 
.A(n_1998),
.B(n_1743),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2039),
.Y(n_2235)
);

INVxp67_ASAP7_75t_L g2236 ( 
.A(n_1986),
.Y(n_2236)
);

AOI22xp33_ASAP7_75t_L g2237 ( 
.A1(n_2164),
.A2(n_1899),
.B1(n_1922),
.B2(n_1843),
.Y(n_2237)
);

INVx3_ASAP7_75t_L g2238 ( 
.A(n_2103),
.Y(n_2238)
);

INVx6_ASAP7_75t_L g2239 ( 
.A(n_2172),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1978),
.B(n_1843),
.Y(n_2240)
);

AOI21xp5_ASAP7_75t_L g2241 ( 
.A1(n_2109),
.A2(n_1813),
.B(n_1800),
.Y(n_2241)
);

INVx5_ASAP7_75t_L g2242 ( 
.A(n_1998),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_1991),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1978),
.B(n_2170),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_2110),
.B(n_1738),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1976),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2045),
.Y(n_2247)
);

INVx5_ASAP7_75t_L g2248 ( 
.A(n_1998),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1977),
.Y(n_2249)
);

AOI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_2037),
.A2(n_1738),
.B1(n_1744),
.B2(n_1899),
.Y(n_2250)
);

NAND3xp33_ASAP7_75t_L g2251 ( 
.A(n_2186),
.B(n_1744),
.C(n_1946),
.Y(n_2251)
);

BUFx3_ASAP7_75t_L g2252 ( 
.A(n_2005),
.Y(n_2252)
);

INVx2_ASAP7_75t_SL g2253 ( 
.A(n_2035),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2048),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_1985),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2063),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_1991),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_2110),
.B(n_1752),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_SL g2259 ( 
.A(n_2138),
.B(n_1752),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2067),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2071),
.B(n_1705),
.Y(n_2261)
);

INVx5_ASAP7_75t_L g2262 ( 
.A(n_2198),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2072),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2013),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2088),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2079),
.B(n_1705),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2023),
.B(n_1705),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_2138),
.B(n_1763),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2108),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2001),
.B(n_1898),
.Y(n_2270)
);

INVx2_ASAP7_75t_SL g2271 ( 
.A(n_1996),
.Y(n_2271)
);

INVxp67_ASAP7_75t_SL g2272 ( 
.A(n_2195),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_1991),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2115),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2180),
.B(n_1898),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2019),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2114),
.B(n_1946),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_2031),
.Y(n_2278)
);

NOR2xp33_ASAP7_75t_L g2279 ( 
.A(n_2062),
.B(n_1787),
.Y(n_2279)
);

AND2x4_ASAP7_75t_L g2280 ( 
.A(n_2177),
.B(n_2208),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2145),
.B(n_1867),
.Y(n_2281)
);

AOI22x1_ASAP7_75t_L g2282 ( 
.A1(n_2032),
.A2(n_1833),
.B1(n_1834),
.B2(n_1831),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2070),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2122),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2145),
.B(n_1867),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2154),
.B(n_1763),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_2208),
.B(n_1962),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2085),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2129),
.Y(n_2289)
);

BUFx6f_ASAP7_75t_L g2290 ( 
.A(n_2031),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2127),
.B(n_1792),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2130),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2193),
.B(n_1792),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2140),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2141),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2069),
.B(n_1843),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2096),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2096),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_2064),
.B(n_1787),
.Y(n_2299)
);

OAI22xp5_ASAP7_75t_SL g2300 ( 
.A1(n_2194),
.A2(n_1916),
.B1(n_760),
.B2(n_788),
.Y(n_2300)
);

NOR3xp33_ASAP7_75t_SL g2301 ( 
.A(n_1984),
.B(n_738),
.C(n_736),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1967),
.B(n_1804),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1967),
.B(n_1887),
.Y(n_2303)
);

INVxp67_ASAP7_75t_L g2304 ( 
.A(n_2128),
.Y(n_2304)
);

INVx2_ASAP7_75t_SL g2305 ( 
.A(n_2163),
.Y(n_2305)
);

OR2x2_ASAP7_75t_L g2306 ( 
.A(n_2018),
.B(n_1823),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_SL g2307 ( 
.A(n_1965),
.B(n_1823),
.Y(n_2307)
);

HB1xp67_ASAP7_75t_L g2308 ( 
.A(n_2086),
.Y(n_2308)
);

BUFx6f_ASAP7_75t_L g2309 ( 
.A(n_2031),
.Y(n_2309)
);

NOR2xp33_ASAP7_75t_L g2310 ( 
.A(n_1972),
.B(n_1878),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2097),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2095),
.B(n_1887),
.Y(n_2312)
);

INVx4_ASAP7_75t_L g2313 ( 
.A(n_2183),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2089),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2092),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2097),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1981),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2095),
.B(n_1831),
.Y(n_2318)
);

O2A1O1Ixp33_ASAP7_75t_L g2319 ( 
.A1(n_2178),
.A2(n_1803),
.B(n_1818),
.C(n_1854),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2049),
.B(n_1726),
.Y(n_2320)
);

AOI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_2210),
.A2(n_1803),
.B1(n_1818),
.B2(n_1851),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2195),
.B(n_1834),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1983),
.Y(n_2323)
);

BUFx6f_ASAP7_75t_L g2324 ( 
.A(n_2183),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2046),
.B(n_1878),
.Y(n_2325)
);

NOR2xp33_ASAP7_75t_L g2326 ( 
.A(n_2219),
.B(n_1851),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1990),
.Y(n_2327)
);

OR2x6_ASAP7_75t_L g2328 ( 
.A(n_2198),
.B(n_2041),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2179),
.B(n_1838),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1997),
.Y(n_2330)
);

BUFx3_ASAP7_75t_L g2331 ( 
.A(n_2036),
.Y(n_2331)
);

OAI22xp33_ASAP7_75t_L g2332 ( 
.A1(n_2008),
.A2(n_1866),
.B1(n_1862),
.B2(n_1846),
.Y(n_2332)
);

AOI22xp33_ASAP7_75t_SL g2333 ( 
.A1(n_1994),
.A2(n_1805),
.B1(n_1862),
.B2(n_873),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_2169),
.B(n_1725),
.Y(n_2334)
);

INVx2_ASAP7_75t_SL g2335 ( 
.A(n_2059),
.Y(n_2335)
);

INVx1_ASAP7_75t_SL g2336 ( 
.A(n_2047),
.Y(n_2336)
);

HB1xp67_ASAP7_75t_L g2337 ( 
.A(n_2168),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2055),
.B(n_1838),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1999),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2135),
.B(n_1762),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2009),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2061),
.B(n_2125),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2010),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2025),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2150),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2155),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_1960),
.B(n_1841),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2113),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_1968),
.B(n_1973),
.Y(n_2349)
);

OR2x2_ASAP7_75t_L g2350 ( 
.A(n_2160),
.B(n_1796),
.Y(n_2350)
);

HB1xp67_ASAP7_75t_L g2351 ( 
.A(n_2148),
.Y(n_2351)
);

AOI22xp33_ASAP7_75t_L g2352 ( 
.A1(n_2209),
.A2(n_1908),
.B1(n_1894),
.B2(n_1825),
.Y(n_2352)
);

BUFx6f_ASAP7_75t_L g2353 ( 
.A(n_2183),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2165),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2182),
.Y(n_2355)
);

AOI22xp33_ASAP7_75t_L g2356 ( 
.A1(n_2206),
.A2(n_1908),
.B1(n_1894),
.B2(n_1825),
.Y(n_2356)
);

AOI22xp33_ASAP7_75t_L g2357 ( 
.A1(n_2184),
.A2(n_1877),
.B1(n_1881),
.B2(n_1796),
.Y(n_2357)
);

BUFx3_ASAP7_75t_L g2358 ( 
.A(n_2076),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_1960),
.B(n_1841),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_1964),
.B(n_1852),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2212),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2218),
.Y(n_2362)
);

OAI22xp5_ASAP7_75t_L g2363 ( 
.A1(n_2074),
.A2(n_1881),
.B1(n_1884),
.B2(n_1877),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_2144),
.Y(n_2364)
);

BUFx3_ASAP7_75t_L g2365 ( 
.A(n_2172),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_1964),
.B(n_1852),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_1975),
.B(n_1860),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_1989),
.B(n_1725),
.Y(n_2368)
);

OAI22xp5_ASAP7_75t_L g2369 ( 
.A1(n_1975),
.A2(n_1884),
.B1(n_1955),
.B2(n_1865),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2117),
.Y(n_2370)
);

INVx2_ASAP7_75t_SL g2371 ( 
.A(n_2078),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2131),
.Y(n_2372)
);

AOI22xp33_ASAP7_75t_L g2373 ( 
.A1(n_2205),
.A2(n_1854),
.B1(n_1940),
.B2(n_1944),
.Y(n_2373)
);

OR2x2_ASAP7_75t_L g2374 ( 
.A(n_2078),
.B(n_1860),
.Y(n_2374)
);

INVx1_ASAP7_75t_SL g2375 ( 
.A(n_2087),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2222),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2143),
.B(n_1865),
.Y(n_2377)
);

BUFx2_ASAP7_75t_L g2378 ( 
.A(n_2166),
.Y(n_2378)
);

NOR2xp33_ASAP7_75t_L g2379 ( 
.A(n_2068),
.B(n_1758),
.Y(n_2379)
);

HB1xp67_ASAP7_75t_L g2380 ( 
.A(n_1959),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2007),
.B(n_1868),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2087),
.B(n_1868),
.Y(n_2382)
);

O2A1O1Ixp5_ASAP7_75t_L g2383 ( 
.A1(n_2106),
.A2(n_1879),
.B(n_1903),
.C(n_1874),
.Y(n_2383)
);

AND2x6_ASAP7_75t_SL g2384 ( 
.A(n_2021),
.B(n_676),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_SL g2385 ( 
.A(n_2015),
.B(n_1731),
.Y(n_2385)
);

INVx1_ASAP7_75t_SL g2386 ( 
.A(n_2105),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_1982),
.B(n_1874),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_1982),
.B(n_1879),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2134),
.Y(n_2389)
);

AND2x4_ASAP7_75t_L g2390 ( 
.A(n_2065),
.B(n_2066),
.Y(n_2390)
);

INVxp67_ASAP7_75t_L g2391 ( 
.A(n_2043),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2111),
.B(n_1903),
.Y(n_2392)
);

BUFx2_ASAP7_75t_L g2393 ( 
.A(n_2166),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2137),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2111),
.B(n_1905),
.Y(n_2395)
);

HB1xp67_ASAP7_75t_L g2396 ( 
.A(n_2166),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2112),
.B(n_1905),
.Y(n_2397)
);

OAI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_2024),
.A2(n_1919),
.B(n_1907),
.Y(n_2398)
);

BUFx6f_ASAP7_75t_L g2399 ( 
.A(n_2185),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2149),
.Y(n_2400)
);

BUFx2_ASAP7_75t_L g2401 ( 
.A(n_2126),
.Y(n_2401)
);

INVx3_ASAP7_75t_L g2402 ( 
.A(n_2185),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2167),
.B(n_1222),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2156),
.Y(n_2404)
);

AOI22xp33_ASAP7_75t_L g2405 ( 
.A1(n_2100),
.A2(n_1758),
.B1(n_1824),
.B2(n_1771),
.Y(n_2405)
);

BUFx3_ASAP7_75t_L g2406 ( 
.A(n_2041),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2094),
.B(n_1840),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2112),
.B(n_1907),
.Y(n_2408)
);

INVx3_ASAP7_75t_L g2409 ( 
.A(n_2185),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_SL g2410 ( 
.A(n_2203),
.B(n_1731),
.Y(n_2410)
);

NOR2xp33_ASAP7_75t_L g2411 ( 
.A(n_2136),
.B(n_1840),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2197),
.Y(n_2412)
);

BUFx2_ASAP7_75t_L g2413 ( 
.A(n_2041),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2207),
.Y(n_2414)
);

BUFx3_ASAP7_75t_L g2415 ( 
.A(n_2004),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2116),
.B(n_1919),
.Y(n_2416)
);

AOI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_2065),
.A2(n_1955),
.B1(n_1824),
.B2(n_1827),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2116),
.B(n_1926),
.Y(n_2418)
);

NAND2x1p5_ASAP7_75t_L g2419 ( 
.A(n_2066),
.B(n_1883),
.Y(n_2419)
);

INVx3_ASAP7_75t_L g2420 ( 
.A(n_2198),
.Y(n_2420)
);

NOR2xp67_ASAP7_75t_L g2421 ( 
.A(n_1963),
.B(n_1926),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2090),
.B(n_1223),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2093),
.B(n_1741),
.Y(n_2423)
);

INVx3_ASAP7_75t_L g2424 ( 
.A(n_2199),
.Y(n_2424)
);

INVx3_ASAP7_75t_L g2425 ( 
.A(n_2199),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2159),
.B(n_1929),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_L g2427 ( 
.A(n_2002),
.B(n_1771),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_SL g2428 ( 
.A(n_2098),
.B(n_1731),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_1974),
.Y(n_2429)
);

INVxp67_ASAP7_75t_L g2430 ( 
.A(n_2142),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2216),
.Y(n_2431)
);

AOI22xp33_ASAP7_75t_L g2432 ( 
.A1(n_1979),
.A2(n_2176),
.B1(n_2173),
.B2(n_2123),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_1987),
.B(n_1741),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2216),
.Y(n_2434)
);

INVx5_ASAP7_75t_L g2435 ( 
.A(n_2146),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_SL g2436 ( 
.A(n_1988),
.B(n_1731),
.Y(n_2436)
);

NAND2x1p5_ASAP7_75t_L g2437 ( 
.A(n_2022),
.B(n_1813),
.Y(n_2437)
);

INVx3_ASAP7_75t_L g2438 ( 
.A(n_2146),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2080),
.B(n_1929),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2223),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2223),
.Y(n_2441)
);

OAI22xp5_ASAP7_75t_L g2442 ( 
.A1(n_1980),
.A2(n_1955),
.B1(n_1941),
.B2(n_1953),
.Y(n_2442)
);

AND2x4_ASAP7_75t_L g2443 ( 
.A(n_2171),
.B(n_2174),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2029),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2118),
.Y(n_2445)
);

INVx2_ASAP7_75t_SL g2446 ( 
.A(n_2021),
.Y(n_2446)
);

AND2x4_ASAP7_75t_L g2447 ( 
.A(n_2033),
.B(n_1741),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_1969),
.B(n_1224),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2119),
.Y(n_2449)
);

OAI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_2057),
.A2(n_1943),
.B(n_1941),
.Y(n_2450)
);

NOR2xp33_ASAP7_75t_L g2451 ( 
.A(n_2220),
.B(n_1944),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2021),
.B(n_1234),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2080),
.B(n_2082),
.Y(n_2453)
);

INVx5_ASAP7_75t_L g2454 ( 
.A(n_2146),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2120),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2124),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2132),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2342),
.B(n_2151),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_SL g2459 ( 
.A(n_2250),
.B(n_1988),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_SL g2460 ( 
.A(n_2237),
.B(n_1988),
.Y(n_2460)
);

NAND2xp33_ASAP7_75t_SL g2461 ( 
.A(n_2227),
.B(n_2152),
.Y(n_2461)
);

NAND2xp33_ASAP7_75t_SL g2462 ( 
.A(n_2301),
.B(n_2152),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_SL g2463 ( 
.A(n_2286),
.B(n_2291),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_SL g2464 ( 
.A(n_2244),
.B(n_1988),
.Y(n_2464)
);

AND2x4_ASAP7_75t_L g2465 ( 
.A(n_2234),
.B(n_2044),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2444),
.B(n_2261),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2244),
.B(n_1988),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_SL g2468 ( 
.A(n_2266),
.B(n_1988),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_SL g2469 ( 
.A(n_2304),
.B(n_2003),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_SL g2470 ( 
.A(n_2336),
.B(n_2000),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_SL g2471 ( 
.A(n_2336),
.B(n_2052),
.Y(n_2471)
);

NAND2xp33_ASAP7_75t_SL g2472 ( 
.A(n_2340),
.B(n_2175),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_SL g2473 ( 
.A(n_2305),
.B(n_2073),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_SL g2474 ( 
.A(n_2224),
.B(n_1970),
.Y(n_2474)
);

AND2x2_ASAP7_75t_SL g2475 ( 
.A(n_2299),
.B(n_2042),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2267),
.B(n_2162),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2297),
.B(n_2196),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_SL g2478 ( 
.A(n_2224),
.B(n_1966),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2234),
.B(n_2158),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2298),
.B(n_2196),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2375),
.B(n_1995),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_SL g2482 ( 
.A(n_2375),
.B(n_2332),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_SL g2483 ( 
.A(n_2306),
.B(n_2335),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_2279),
.B(n_2006),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_SL g2485 ( 
.A(n_2326),
.B(n_2371),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_2251),
.B(n_1993),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_SL g2487 ( 
.A(n_2325),
.B(n_2253),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_SL g2488 ( 
.A(n_2333),
.B(n_2147),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2311),
.B(n_2200),
.Y(n_2489)
);

AND2x4_ASAP7_75t_L g2490 ( 
.A(n_2234),
.B(n_2213),
.Y(n_2490)
);

NAND2xp33_ASAP7_75t_SL g2491 ( 
.A(n_2277),
.B(n_2175),
.Y(n_2491)
);

NAND2xp33_ASAP7_75t_SL g2492 ( 
.A(n_2270),
.B(n_2217),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_SL g2493 ( 
.A(n_2293),
.B(n_2139),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2316),
.B(n_2202),
.Y(n_2494)
);

NAND2xp33_ASAP7_75t_SL g2495 ( 
.A(n_2275),
.B(n_2350),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_SL g2496 ( 
.A(n_2386),
.B(n_2016),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2431),
.B(n_2202),
.Y(n_2497)
);

AND2x4_ASAP7_75t_L g2498 ( 
.A(n_2328),
.B(n_2081),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_SL g2499 ( 
.A(n_2386),
.B(n_2017),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_SL g2500 ( 
.A(n_2310),
.B(n_2026),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_2349),
.B(n_2161),
.Y(n_2501)
);

NAND2xp33_ASAP7_75t_SL g2502 ( 
.A(n_2368),
.B(n_2181),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_SL g2503 ( 
.A(n_2349),
.B(n_2430),
.Y(n_2503)
);

NAND2xp33_ASAP7_75t_SL g2504 ( 
.A(n_2320),
.B(n_2232),
.Y(n_2504)
);

NAND2xp33_ASAP7_75t_SL g2505 ( 
.A(n_2307),
.B(n_2374),
.Y(n_2505)
);

NOR2xp33_ASAP7_75t_L g2506 ( 
.A(n_2236),
.B(n_1992),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_SL g2507 ( 
.A(n_2287),
.B(n_2187),
.Y(n_2507)
);

AND2x4_ASAP7_75t_L g2508 ( 
.A(n_2328),
.B(n_2083),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_SL g2509 ( 
.A(n_2287),
.B(n_2188),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_SL g2510 ( 
.A(n_2391),
.B(n_2012),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_2308),
.B(n_2133),
.Y(n_2511)
);

AND2x2_ASAP7_75t_SL g2512 ( 
.A(n_2443),
.B(n_2190),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_SL g2513 ( 
.A(n_2280),
.B(n_2153),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_2280),
.B(n_2075),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_SL g2515 ( 
.A(n_2351),
.B(n_2030),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_SL g2516 ( 
.A(n_2337),
.B(n_2034),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_SL g2517 ( 
.A(n_2390),
.B(n_2038),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_SL g2518 ( 
.A(n_2390),
.B(n_2040),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_SL g2519 ( 
.A(n_2321),
.B(n_2053),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_SL g2520 ( 
.A(n_2271),
.B(n_2056),
.Y(n_2520)
);

AND2x4_ASAP7_75t_L g2521 ( 
.A(n_2328),
.B(n_2104),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_SL g2522 ( 
.A(n_2382),
.B(n_2379),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_SL g2523 ( 
.A(n_2403),
.B(n_2058),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2434),
.B(n_2200),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2364),
.B(n_2448),
.Y(n_2525)
);

AND3x1_ASAP7_75t_L g2526 ( 
.A(n_2446),
.B(n_692),
.C(n_681),
.Y(n_2526)
);

NAND2xp33_ASAP7_75t_SL g2527 ( 
.A(n_2228),
.B(n_2107),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_L g2528 ( 
.A(n_2380),
.B(n_2091),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_2378),
.B(n_2204),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2440),
.B(n_2204),
.Y(n_2530)
);

NAND2xp33_ASAP7_75t_SL g2531 ( 
.A(n_2235),
.B(n_2099),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_SL g2532 ( 
.A(n_2393),
.B(n_2211),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_SL g2533 ( 
.A(n_2247),
.B(n_2211),
.Y(n_2533)
);

AND2x4_ASAP7_75t_L g2534 ( 
.A(n_2242),
.B(n_2248),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2441),
.B(n_2214),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_SL g2536 ( 
.A(n_2254),
.B(n_2214),
.Y(n_2536)
);

NAND2xp33_ASAP7_75t_SL g2537 ( 
.A(n_2256),
.B(n_2099),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_2260),
.B(n_2263),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_SL g2539 ( 
.A(n_2265),
.B(n_2101),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_2269),
.B(n_2101),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_SL g2541 ( 
.A(n_2274),
.B(n_2102),
.Y(n_2541)
);

NAND2xp33_ASAP7_75t_SL g2542 ( 
.A(n_2284),
.B(n_2289),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_SL g2543 ( 
.A(n_2292),
.B(n_2102),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_SL g2544 ( 
.A(n_2294),
.B(n_2107),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_SL g2545 ( 
.A(n_2295),
.B(n_1761),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2272),
.B(n_2082),
.Y(n_2546)
);

AND2x2_ASAP7_75t_L g2547 ( 
.A(n_2422),
.B(n_2123),
.Y(n_2547)
);

NAND2xp33_ASAP7_75t_SL g2548 ( 
.A(n_2317),
.B(n_2011),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_SL g2549 ( 
.A(n_2331),
.B(n_1761),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_SL g2550 ( 
.A(n_2358),
.B(n_1761),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_SL g2551 ( 
.A(n_2443),
.B(n_1761),
.Y(n_2551)
);

NAND2xp33_ASAP7_75t_L g2552 ( 
.A(n_2242),
.B(n_2146),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2312),
.B(n_2084),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2312),
.B(n_2084),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_SL g2555 ( 
.A(n_2323),
.B(n_1785),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_SL g2556 ( 
.A(n_2327),
.B(n_1785),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2445),
.B(n_2189),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2449),
.B(n_2077),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_SL g2559 ( 
.A(n_2330),
.B(n_1785),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_SL g2560 ( 
.A(n_2339),
.B(n_1785),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_SL g2561 ( 
.A(n_2341),
.B(n_1797),
.Y(n_2561)
);

AND2x4_ASAP7_75t_L g2562 ( 
.A(n_2242),
.B(n_2060),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2455),
.B(n_2077),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_SL g2564 ( 
.A(n_2343),
.B(n_1797),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_SL g2565 ( 
.A(n_2344),
.B(n_1797),
.Y(n_2565)
);

AND2x4_ASAP7_75t_L g2566 ( 
.A(n_2242),
.B(n_2014),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2456),
.B(n_1980),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2457),
.B(n_1943),
.Y(n_2568)
);

NAND2xp33_ASAP7_75t_SL g2569 ( 
.A(n_2324),
.B(n_2020),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_SL g2570 ( 
.A(n_2245),
.B(n_1797),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_SL g2571 ( 
.A(n_2252),
.B(n_1809),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_SL g2572 ( 
.A(n_2427),
.B(n_1809),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_SL g2573 ( 
.A(n_2300),
.B(n_1809),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_SL g2574 ( 
.A(n_2225),
.B(n_1809),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_SL g2575 ( 
.A(n_2396),
.B(n_1837),
.Y(n_2575)
);

NAND2xp33_ASAP7_75t_SL g2576 ( 
.A(n_2324),
.B(n_2191),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2377),
.B(n_1953),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_SL g2578 ( 
.A(n_2435),
.B(n_1837),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_SL g2579 ( 
.A(n_2435),
.B(n_1837),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_SL g2580 ( 
.A(n_2435),
.B(n_1837),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_SL g2581 ( 
.A(n_2435),
.B(n_1827),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2452),
.B(n_1272),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_SL g2583 ( 
.A(n_2454),
.B(n_1937),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2454),
.B(n_1937),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2338),
.B(n_2146),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2454),
.B(n_1937),
.Y(n_2586)
);

AND2x4_ASAP7_75t_L g2587 ( 
.A(n_2248),
.B(n_2192),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_SL g2588 ( 
.A(n_2454),
.B(n_1957),
.Y(n_2588)
);

AND2x4_ASAP7_75t_L g2589 ( 
.A(n_2248),
.B(n_2201),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_SL g2590 ( 
.A(n_2411),
.B(n_2281),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_SL g2591 ( 
.A(n_2285),
.B(n_1957),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_SL g2592 ( 
.A(n_2401),
.B(n_1957),
.Y(n_2592)
);

NAND2xp33_ASAP7_75t_SL g2593 ( 
.A(n_2324),
.B(n_1822),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_SL g2594 ( 
.A(n_2413),
.B(n_1849),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_SL g2595 ( 
.A(n_2407),
.B(n_2429),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_SL g2596 ( 
.A(n_2421),
.B(n_1849),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_SL g2597 ( 
.A(n_2451),
.B(n_2258),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_2259),
.B(n_1883),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_SL g2599 ( 
.A(n_2268),
.B(n_1886),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2338),
.B(n_2057),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2406),
.B(n_705),
.Y(n_2601)
);

NAND2xp33_ASAP7_75t_SL g2602 ( 
.A(n_2353),
.B(n_2399),
.Y(n_2602)
);

NAND2xp33_ASAP7_75t_SL g2603 ( 
.A(n_2353),
.B(n_1886),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_SL g2604 ( 
.A(n_2233),
.B(n_2238),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_SL g2605 ( 
.A(n_2233),
.B(n_1822),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_SL g2606 ( 
.A(n_2238),
.B(n_1896),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_SL g2607 ( 
.A(n_2229),
.B(n_1896),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_SL g2608 ( 
.A(n_2229),
.B(n_729),
.Y(n_2608)
);

NAND2xp33_ASAP7_75t_SL g2609 ( 
.A(n_2353),
.B(n_2051),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_SL g2610 ( 
.A(n_2229),
.B(n_729),
.Y(n_2610)
);

NAND2xp33_ASAP7_75t_SL g2611 ( 
.A(n_2399),
.B(n_2054),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_SL g2612 ( 
.A(n_2230),
.B(n_2231),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_SL g2613 ( 
.A(n_2230),
.B(n_729),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_2230),
.B(n_729),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_2231),
.B(n_783),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2246),
.B(n_783),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_SL g2617 ( 
.A(n_2231),
.B(n_783),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2303),
.B(n_2121),
.Y(n_2618)
);

NAND2xp33_ASAP7_75t_SL g2619 ( 
.A(n_2399),
.B(n_2157),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_SL g2620 ( 
.A(n_2243),
.B(n_783),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_SL g2621 ( 
.A(n_2243),
.B(n_818),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_SL g2622 ( 
.A(n_2243),
.B(n_818),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_SL g2623 ( 
.A(n_2257),
.B(n_818),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_SL g2624 ( 
.A(n_2257),
.B(n_818),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_SL g2625 ( 
.A(n_2257),
.B(n_2273),
.Y(n_2625)
);

NAND2xp33_ASAP7_75t_SL g2626 ( 
.A(n_2273),
.B(n_2215),
.Y(n_2626)
);

NAND2xp33_ASAP7_75t_SL g2627 ( 
.A(n_2273),
.B(n_2221),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_SL g2628 ( 
.A(n_2278),
.B(n_999),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_SL g2629 ( 
.A(n_2278),
.B(n_999),
.Y(n_2629)
);

NAND2xp33_ASAP7_75t_SL g2630 ( 
.A(n_2278),
.B(n_739),
.Y(n_2630)
);

NAND2xp33_ASAP7_75t_SL g2631 ( 
.A(n_2290),
.B(n_740),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_SL g2632 ( 
.A(n_2290),
.B(n_999),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2303),
.B(n_1538),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2302),
.B(n_1538),
.Y(n_2634)
);

NAND2xp33_ASAP7_75t_SL g2635 ( 
.A(n_2290),
.B(n_741),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_2309),
.B(n_999),
.Y(n_2636)
);

NAND2xp33_ASAP7_75t_SL g2637 ( 
.A(n_2309),
.B(n_742),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2249),
.B(n_1026),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_2309),
.B(n_1026),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_SL g2640 ( 
.A(n_2356),
.B(n_1026),
.Y(n_2640)
);

AND2x4_ASAP7_75t_L g2641 ( 
.A(n_2248),
.B(n_1616),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2302),
.B(n_2318),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_SL g2643 ( 
.A(n_2262),
.B(n_1026),
.Y(n_2643)
);

NAND2xp33_ASAP7_75t_SL g2644 ( 
.A(n_2420),
.B(n_2313),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_SL g2645 ( 
.A(n_2262),
.B(n_743),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_SL g2646 ( 
.A(n_2262),
.B(n_745),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_SL g2647 ( 
.A(n_2262),
.B(n_746),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2318),
.B(n_2322),
.Y(n_2648)
);

NAND2xp33_ASAP7_75t_SL g2649 ( 
.A(n_2420),
.B(n_748),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_SL g2650 ( 
.A(n_2432),
.B(n_750),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_SL g2651 ( 
.A(n_2319),
.B(n_751),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_SL g2652 ( 
.A(n_2423),
.B(n_753),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_SL g2653 ( 
.A(n_2423),
.B(n_755),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_SL g2654 ( 
.A(n_2357),
.B(n_757),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_SL g2655 ( 
.A(n_2345),
.B(n_758),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_SL g2656 ( 
.A(n_2346),
.B(n_761),
.Y(n_2656)
);

NAND2xp33_ASAP7_75t_SL g2657 ( 
.A(n_2313),
.B(n_763),
.Y(n_2657)
);

AND2x2_ASAP7_75t_SL g2658 ( 
.A(n_2381),
.B(n_681),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_SL g2659 ( 
.A(n_2354),
.B(n_764),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_SL g2660 ( 
.A(n_2355),
.B(n_2361),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_SL g2661 ( 
.A(n_2362),
.B(n_765),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_SL g2662 ( 
.A(n_2376),
.B(n_2385),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_SL g2663 ( 
.A(n_2296),
.B(n_767),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_SL g2664 ( 
.A(n_2240),
.B(n_1674),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_SL g2665 ( 
.A(n_2240),
.B(n_1564),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2322),
.B(n_1546),
.Y(n_2666)
);

NAND2xp33_ASAP7_75t_SL g2667 ( 
.A(n_2410),
.B(n_775),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_SL g2668 ( 
.A(n_2296),
.B(n_778),
.Y(n_2668)
);

NAND2xp33_ASAP7_75t_SL g2669 ( 
.A(n_2334),
.B(n_779),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_SL g2670 ( 
.A(n_2415),
.B(n_785),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_SL g2671 ( 
.A(n_2405),
.B(n_2255),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_SL g2672 ( 
.A(n_2264),
.B(n_787),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_SL g2673 ( 
.A(n_2276),
.B(n_790),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_SL g2674 ( 
.A(n_2283),
.B(n_792),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_2288),
.B(n_797),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_SL g2676 ( 
.A(n_2314),
.B(n_798),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_SL g2677 ( 
.A(n_2315),
.B(n_799),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2348),
.B(n_1267),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_SL g2679 ( 
.A(n_2370),
.B(n_800),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2372),
.B(n_1267),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_SL g2681 ( 
.A(n_2404),
.B(n_2412),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_SL g2682 ( 
.A(n_2389),
.B(n_801),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2367),
.B(n_1546),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_SL g2684 ( 
.A(n_2394),
.B(n_802),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_SL g2685 ( 
.A(n_2400),
.B(n_804),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_SL g2686 ( 
.A(n_2414),
.B(n_807),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_SL g2687 ( 
.A(n_2373),
.B(n_810),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_SL g2688 ( 
.A(n_2352),
.B(n_811),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2367),
.B(n_1550),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_SL g2690 ( 
.A(n_2417),
.B(n_816),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_SL g2691 ( 
.A(n_2363),
.B(n_817),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_SL g2692 ( 
.A(n_2363),
.B(n_819),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_SL g2693 ( 
.A(n_2453),
.B(n_820),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_SL g2694 ( 
.A(n_2453),
.B(n_822),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_SL g2695 ( 
.A(n_2433),
.B(n_824),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_SL g2696 ( 
.A(n_2433),
.B(n_825),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_SL g2697 ( 
.A(n_2447),
.B(n_2402),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_SL g2698 ( 
.A(n_2447),
.B(n_826),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2329),
.B(n_1550),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_SL g2700 ( 
.A(n_2402),
.B(n_829),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_SL g2701 ( 
.A(n_2409),
.B(n_832),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_SL g2702 ( 
.A(n_2409),
.B(n_833),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2365),
.B(n_692),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_SL g2704 ( 
.A(n_2438),
.B(n_2369),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2239),
.B(n_698),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_SL g2706 ( 
.A(n_2438),
.B(n_834),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_SL g2707 ( 
.A(n_2369),
.B(n_836),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2241),
.B(n_1564),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_SL g2709 ( 
.A(n_2392),
.B(n_1564),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2329),
.B(n_1555),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_SL g2711 ( 
.A(n_2392),
.B(n_2395),
.Y(n_2711)
);

AOI22xp5_ASAP7_75t_L g2712 ( 
.A1(n_2491),
.A2(n_2239),
.B1(n_2442),
.B2(n_838),
.Y(n_2712)
);

OAI22xp5_ASAP7_75t_L g2713 ( 
.A1(n_2475),
.A2(n_2437),
.B1(n_2419),
.B2(n_2442),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2568),
.Y(n_2714)
);

AND2x4_ASAP7_75t_L g2715 ( 
.A(n_2498),
.B(n_2424),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2538),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2477),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2466),
.B(n_2387),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2547),
.B(n_2387),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2678),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_2461),
.Y(n_2721)
);

AND2x4_ASAP7_75t_L g2722 ( 
.A(n_2498),
.B(n_2508),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2658),
.B(n_2388),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2680),
.Y(n_2724)
);

OR2x2_ASAP7_75t_L g2725 ( 
.A(n_2503),
.B(n_2360),
.Y(n_2725)
);

NAND2xp33_ASAP7_75t_L g2726 ( 
.A(n_2558),
.B(n_2419),
.Y(n_2726)
);

AND3x1_ASAP7_75t_SL g2727 ( 
.A(n_2658),
.B(n_699),
.C(n_698),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2582),
.B(n_699),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2660),
.Y(n_2729)
);

HB1xp67_ASAP7_75t_L g2730 ( 
.A(n_2464),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2480),
.Y(n_2731)
);

NOR2xp33_ASAP7_75t_L g2732 ( 
.A(n_2482),
.B(n_2384),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2463),
.B(n_2458),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2681),
.Y(n_2734)
);

INVx6_ASAP7_75t_L g2735 ( 
.A(n_2534),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2616),
.B(n_707),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2463),
.B(n_2528),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2595),
.Y(n_2738)
);

INVx8_ASAP7_75t_L g2739 ( 
.A(n_2534),
.Y(n_2739)
);

INVx4_ASAP7_75t_L g2740 ( 
.A(n_2534),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2638),
.B(n_707),
.Y(n_2741)
);

AND2x4_ASAP7_75t_L g2742 ( 
.A(n_2498),
.B(n_2424),
.Y(n_2742)
);

INVx3_ASAP7_75t_L g2743 ( 
.A(n_2641),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2533),
.Y(n_2744)
);

CKINVDCx5p33_ASAP7_75t_R g2745 ( 
.A(n_2472),
.Y(n_2745)
);

BUFx12f_ASAP7_75t_L g2746 ( 
.A(n_2703),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2590),
.B(n_2388),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2483),
.B(n_2522),
.Y(n_2748)
);

AND2x4_ASAP7_75t_SL g2749 ( 
.A(n_2508),
.B(n_2425),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2705),
.B(n_2601),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2489),
.B(n_2395),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2494),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2536),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_SL g2754 ( 
.A(n_2475),
.B(n_2226),
.Y(n_2754)
);

NOR2xp33_ASAP7_75t_R g2755 ( 
.A(n_2504),
.B(n_2425),
.Y(n_2755)
);

CKINVDCx11_ASAP7_75t_R g2756 ( 
.A(n_2508),
.Y(n_2756)
);

CKINVDCx20_ASAP7_75t_R g2757 ( 
.A(n_2462),
.Y(n_2757)
);

AOI22xp5_ASAP7_75t_L g2758 ( 
.A1(n_2505),
.A2(n_844),
.B1(n_847),
.B2(n_837),
.Y(n_2758)
);

BUFx8_ASAP7_75t_L g2759 ( 
.A(n_2521),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2497),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2485),
.B(n_2525),
.Y(n_2761)
);

BUFx2_ASAP7_75t_L g2762 ( 
.A(n_2630),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2524),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_SL g2764 ( 
.A(n_2495),
.B(n_2397),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_SL g2765 ( 
.A(n_2484),
.B(n_2512),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_2512),
.B(n_2397),
.Y(n_2766)
);

BUFx4f_ASAP7_75t_L g2767 ( 
.A(n_2521),
.Y(n_2767)
);

AOI21xp33_ASAP7_75t_L g2768 ( 
.A1(n_2691),
.A2(n_2426),
.B(n_2282),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2530),
.B(n_2408),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2516),
.B(n_708),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2539),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2535),
.B(n_2408),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2540),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2541),
.Y(n_2774)
);

HB1xp67_ASAP7_75t_L g2775 ( 
.A(n_2464),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_2506),
.Y(n_2776)
);

BUFx3_ASAP7_75t_L g2777 ( 
.A(n_2521),
.Y(n_2777)
);

BUFx2_ASAP7_75t_L g2778 ( 
.A(n_2631),
.Y(n_2778)
);

O2A1O1Ixp33_ASAP7_75t_L g2779 ( 
.A1(n_2488),
.A2(n_711),
.B(n_714),
.C(n_708),
.Y(n_2779)
);

BUFx2_ASAP7_75t_L g2780 ( 
.A(n_2635),
.Y(n_2780)
);

AOI22xp33_ASAP7_75t_L g2781 ( 
.A1(n_2692),
.A2(n_2640),
.B1(n_2650),
.B2(n_2669),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2543),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_SL g2783 ( 
.A(n_2476),
.B(n_2416),
.Y(n_2783)
);

INVx4_ASAP7_75t_L g2784 ( 
.A(n_2641),
.Y(n_2784)
);

OR2x2_ASAP7_75t_L g2785 ( 
.A(n_2515),
.B(n_2360),
.Y(n_2785)
);

CKINVDCx5p33_ASAP7_75t_R g2786 ( 
.A(n_2487),
.Y(n_2786)
);

BUFx4f_ASAP7_75t_L g2787 ( 
.A(n_2465),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2544),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2642),
.B(n_2416),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2563),
.B(n_2693),
.Y(n_2790)
);

BUFx3_ASAP7_75t_L g2791 ( 
.A(n_2465),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2694),
.B(n_711),
.Y(n_2792)
);

OAI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_2567),
.A2(n_2437),
.B1(n_2418),
.B2(n_2428),
.Y(n_2793)
);

OAI22xp5_ASAP7_75t_L g2794 ( 
.A1(n_2546),
.A2(n_2418),
.B1(n_2439),
.B2(n_2366),
.Y(n_2794)
);

OR2x6_ASAP7_75t_L g2795 ( 
.A(n_2465),
.B(n_2398),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2542),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2633),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_SL g2798 ( 
.A(n_2618),
.B(n_2366),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2511),
.Y(n_2799)
);

OAI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2574),
.A2(n_2439),
.B1(n_2359),
.B2(n_2347),
.Y(n_2800)
);

BUFx6f_ASAP7_75t_L g2801 ( 
.A(n_2490),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2529),
.B(n_714),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2597),
.B(n_2347),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2648),
.B(n_2359),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2532),
.B(n_721),
.Y(n_2805)
);

AND2x4_ASAP7_75t_L g2806 ( 
.A(n_2490),
.B(n_2436),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2470),
.B(n_848),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2698),
.B(n_721),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2695),
.B(n_723),
.Y(n_2809)
);

INVxp67_ASAP7_75t_L g2810 ( 
.A(n_2612),
.Y(n_2810)
);

OAI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2473),
.A2(n_2398),
.B1(n_2450),
.B2(n_851),
.Y(n_2811)
);

NAND2x1p5_ASAP7_75t_L g2812 ( 
.A(n_2551),
.B(n_1616),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2696),
.B(n_723),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2526),
.B(n_2652),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2666),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_L g2816 ( 
.A(n_2471),
.B(n_2450),
.Y(n_2816)
);

CKINVDCx20_ASAP7_75t_R g2817 ( 
.A(n_2637),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2653),
.B(n_727),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2520),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2662),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2699),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_SL g2822 ( 
.A(n_2492),
.B(n_2383),
.Y(n_2822)
);

BUFx3_ASAP7_75t_L g2823 ( 
.A(n_2479),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2469),
.B(n_849),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2553),
.B(n_854),
.Y(n_2825)
);

AND2x2_ASAP7_75t_L g2826 ( 
.A(n_2474),
.B(n_727),
.Y(n_2826)
);

INVxp67_ASAP7_75t_SL g2827 ( 
.A(n_2554),
.Y(n_2827)
);

BUFx4f_ASAP7_75t_L g2828 ( 
.A(n_2479),
.Y(n_2828)
);

BUFx6f_ASAP7_75t_L g2829 ( 
.A(n_2490),
.Y(n_2829)
);

BUFx2_ASAP7_75t_L g2830 ( 
.A(n_2602),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2655),
.B(n_731),
.Y(n_2831)
);

CKINVDCx20_ASAP7_75t_R g2832 ( 
.A(n_2657),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2711),
.B(n_855),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2710),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2683),
.Y(n_2835)
);

BUFx6f_ASAP7_75t_L g2836 ( 
.A(n_2479),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2656),
.B(n_731),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2689),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2711),
.B(n_856),
.Y(n_2839)
);

INVx1_ASAP7_75t_SL g2840 ( 
.A(n_2670),
.Y(n_2840)
);

BUFx3_ASAP7_75t_L g2841 ( 
.A(n_2587),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2523),
.B(n_857),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2478),
.B(n_861),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2577),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2625),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2659),
.B(n_2661),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2557),
.Y(n_2847)
);

BUFx3_ASAP7_75t_L g2848 ( 
.A(n_2587),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2575),
.Y(n_2849)
);

OAI21xp5_ASAP7_75t_L g2850 ( 
.A1(n_2486),
.A2(n_1557),
.B(n_1555),
.Y(n_2850)
);

NOR2xp33_ASAP7_75t_L g2851 ( 
.A(n_2688),
.B(n_2481),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2545),
.Y(n_2852)
);

NAND2x1p5_ASAP7_75t_L g2853 ( 
.A(n_2501),
.B(n_2566),
.Y(n_2853)
);

INVx2_ASAP7_75t_SL g2854 ( 
.A(n_2549),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2608),
.B(n_862),
.Y(n_2855)
);

A2O1A1Ixp33_ASAP7_75t_L g2856 ( 
.A1(n_2527),
.A2(n_2531),
.B(n_2537),
.C(n_2459),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2610),
.B(n_2613),
.Y(n_2857)
);

AND2x4_ASAP7_75t_L g2858 ( 
.A(n_2697),
.B(n_1620),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2555),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2634),
.Y(n_2860)
);

NOR2xp33_ASAP7_75t_L g2861 ( 
.A(n_2514),
.B(n_2663),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2556),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_L g2863 ( 
.A1(n_2707),
.A2(n_744),
.B1(n_747),
.B2(n_732),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2614),
.B(n_732),
.Y(n_2864)
);

A2O1A1Ixp33_ASAP7_75t_L g2865 ( 
.A1(n_2459),
.A2(n_808),
.B(n_839),
.C(n_768),
.Y(n_2865)
);

CKINVDCx5p33_ASAP7_75t_R g2866 ( 
.A(n_2649),
.Y(n_2866)
);

BUFx6f_ASAP7_75t_L g2867 ( 
.A(n_2641),
.Y(n_2867)
);

O2A1O1Ixp33_ASAP7_75t_SL g2868 ( 
.A1(n_2704),
.A2(n_747),
.B(n_768),
.C(n_744),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2585),
.Y(n_2869)
);

AND3x1_ASAP7_75t_SL g2870 ( 
.A(n_2615),
.B(n_774),
.C(n_769),
.Y(n_2870)
);

OAI22xp5_ASAP7_75t_SL g2871 ( 
.A1(n_2566),
.A2(n_878),
.B1(n_880),
.B2(n_863),
.Y(n_2871)
);

HB1xp67_ASAP7_75t_L g2872 ( 
.A(n_2467),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2617),
.B(n_769),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_SL g2874 ( 
.A(n_2548),
.B(n_1557),
.Y(n_2874)
);

AND2x2_ASAP7_75t_L g2875 ( 
.A(n_2620),
.B(n_774),
.Y(n_2875)
);

BUFx6f_ASAP7_75t_L g2876 ( 
.A(n_2587),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2559),
.Y(n_2877)
);

OAI221xp5_ASAP7_75t_L g2878 ( 
.A1(n_2682),
.A2(n_795),
.B1(n_910),
.B2(n_858),
.C(n_827),
.Y(n_2878)
);

OAI22xp5_ASAP7_75t_L g2879 ( 
.A1(n_2573),
.A2(n_882),
.B1(n_884),
.B2(n_881),
.Y(n_2879)
);

CKINVDCx5p33_ASAP7_75t_R g2880 ( 
.A(n_2667),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2621),
.B(n_2622),
.Y(n_2881)
);

BUFx2_ASAP7_75t_L g2882 ( 
.A(n_2576),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_L g2883 ( 
.A(n_2668),
.B(n_888),
.Y(n_2883)
);

CKINVDCx5p33_ASAP7_75t_R g2884 ( 
.A(n_2700),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2623),
.B(n_889),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2560),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2624),
.B(n_891),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2628),
.B(n_781),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_SL g2889 ( 
.A(n_2519),
.B(n_781),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2561),
.Y(n_2890)
);

CKINVDCx16_ASAP7_75t_R g2891 ( 
.A(n_2589),
.Y(n_2891)
);

BUFx2_ASAP7_75t_L g2892 ( 
.A(n_2569),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2467),
.Y(n_2893)
);

NOR2xp33_ASAP7_75t_L g2894 ( 
.A(n_2654),
.B(n_892),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2629),
.B(n_894),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2600),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2632),
.B(n_896),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2709),
.Y(n_2898)
);

INVx2_ASAP7_75t_L g2899 ( 
.A(n_2709),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2636),
.B(n_898),
.Y(n_2900)
);

AND2x2_ASAP7_75t_L g2901 ( 
.A(n_2639),
.B(n_789),
.Y(n_2901)
);

NAND2x1p5_ASAP7_75t_L g2902 ( 
.A(n_2566),
.B(n_1620),
.Y(n_2902)
);

OAI22xp5_ASAP7_75t_SL g2903 ( 
.A1(n_2562),
.A2(n_916),
.B1(n_917),
.B2(n_915),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2671),
.Y(n_2904)
);

CKINVDCx5p33_ASAP7_75t_R g2905 ( 
.A(n_2701),
.Y(n_2905)
);

CKINVDCx5p33_ASAP7_75t_R g2906 ( 
.A(n_2702),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2493),
.B(n_919),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2564),
.Y(n_2908)
);

AND2x2_ASAP7_75t_L g2909 ( 
.A(n_2643),
.B(n_789),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2562),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2565),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2570),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2562),
.Y(n_2913)
);

OAI22xp5_ASAP7_75t_SL g2914 ( 
.A1(n_2589),
.A2(n_925),
.B1(n_927),
.B2(n_921),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2500),
.B(n_929),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_SL g2916 ( 
.A(n_2589),
.B(n_931),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2684),
.B(n_795),
.Y(n_2917)
);

AND2x2_ASAP7_75t_L g2918 ( 
.A(n_2685),
.B(n_803),
.Y(n_2918)
);

NAND2x1_ASAP7_75t_L g2919 ( 
.A(n_2644),
.B(n_1620),
.Y(n_2919)
);

CKINVDCx11_ASAP7_75t_R g2920 ( 
.A(n_2645),
.Y(n_2920)
);

AND2x2_ASAP7_75t_L g2921 ( 
.A(n_2686),
.B(n_803),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2517),
.B(n_937),
.Y(n_2922)
);

AND2x2_ASAP7_75t_L g2923 ( 
.A(n_2690),
.B(n_805),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_SL g2924 ( 
.A(n_2502),
.B(n_805),
.Y(n_2924)
);

INVxp67_ASAP7_75t_L g2925 ( 
.A(n_2550),
.Y(n_2925)
);

OAI22xp5_ASAP7_75t_L g2926 ( 
.A1(n_2672),
.A2(n_939),
.B1(n_949),
.B2(n_938),
.Y(n_2926)
);

CKINVDCx16_ASAP7_75t_R g2927 ( 
.A(n_2609),
.Y(n_2927)
);

AND2x2_ASAP7_75t_L g2928 ( 
.A(n_2673),
.B(n_808),
.Y(n_2928)
);

BUFx2_ASAP7_75t_SL g2929 ( 
.A(n_2571),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2513),
.Y(n_2930)
);

NOR2x1_ASAP7_75t_L g2931 ( 
.A(n_2646),
.B(n_813),
.Y(n_2931)
);

AND2x2_ASAP7_75t_L g2932 ( 
.A(n_2674),
.B(n_813),
.Y(n_2932)
);

INVxp67_ASAP7_75t_L g2933 ( 
.A(n_2675),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2518),
.B(n_2687),
.Y(n_2934)
);

AND2x2_ASAP7_75t_L g2935 ( 
.A(n_2676),
.B(n_815),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2664),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2496),
.B(n_950),
.Y(n_2937)
);

OR2x2_ASAP7_75t_L g2938 ( 
.A(n_2677),
.B(n_815),
.Y(n_2938)
);

BUFx2_ASAP7_75t_L g2939 ( 
.A(n_2611),
.Y(n_2939)
);

INVx4_ASAP7_75t_L g2940 ( 
.A(n_2619),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2499),
.B(n_2679),
.Y(n_2941)
);

OAI22xp5_ASAP7_75t_SL g2942 ( 
.A1(n_2647),
.A2(n_954),
.B1(n_956),
.B2(n_953),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2507),
.B(n_957),
.Y(n_2943)
);

INVx8_ASAP7_75t_L g2944 ( 
.A(n_2626),
.Y(n_2944)
);

O2A1O1Ixp33_ASAP7_75t_L g2945 ( 
.A1(n_2651),
.A2(n_823),
.B(n_827),
.C(n_821),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2509),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2592),
.B(n_821),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2510),
.B(n_961),
.Y(n_2948)
);

BUFx2_ASAP7_75t_L g2949 ( 
.A(n_2627),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2604),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2591),
.Y(n_2951)
);

AND2x2_ASAP7_75t_L g2952 ( 
.A(n_2594),
.B(n_823),
.Y(n_2952)
);

BUFx3_ASAP7_75t_L g2953 ( 
.A(n_2593),
.Y(n_2953)
);

INVx6_ASAP7_75t_L g2954 ( 
.A(n_2603),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2572),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2468),
.B(n_962),
.Y(n_2956)
);

NAND2xp33_ASAP7_75t_L g2957 ( 
.A(n_2706),
.B(n_965),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2607),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2664),
.Y(n_2959)
);

NOR2xp33_ASAP7_75t_L g2960 ( 
.A(n_2468),
.B(n_966),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2665),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2581),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2665),
.B(n_968),
.Y(n_2963)
);

NOR2xp67_ASAP7_75t_L g2964 ( 
.A(n_2596),
.B(n_568),
.Y(n_2964)
);

AOI22xp33_ASAP7_75t_L g2965 ( 
.A1(n_2460),
.A2(n_835),
.B1(n_839),
.B2(n_831),
.Y(n_2965)
);

AOI22xp33_ASAP7_75t_L g2966 ( 
.A1(n_2460),
.A2(n_835),
.B1(n_841),
.B2(n_831),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2598),
.B(n_969),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2599),
.B(n_841),
.Y(n_2968)
);

CKINVDCx5p33_ASAP7_75t_R g2969 ( 
.A(n_2605),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2606),
.B(n_970),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2578),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2579),
.Y(n_2972)
);

CKINVDCx5p33_ASAP7_75t_R g2973 ( 
.A(n_2583),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2580),
.B(n_973),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2708),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2584),
.B(n_843),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2586),
.B(n_974),
.Y(n_2977)
);

CKINVDCx20_ASAP7_75t_R g2978 ( 
.A(n_2588),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2708),
.Y(n_2979)
);

AND2x4_ASAP7_75t_L g2980 ( 
.A(n_2552),
.B(n_1631),
.Y(n_2980)
);

AND2x2_ASAP7_75t_L g2981 ( 
.A(n_2582),
.B(n_843),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2568),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2466),
.B(n_976),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2466),
.B(n_979),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2568),
.Y(n_2985)
);

OAI22xp5_ASAP7_75t_SL g2986 ( 
.A1(n_2526),
.A2(n_987),
.B1(n_988),
.B2(n_980),
.Y(n_2986)
);

NAND2x1p5_ASAP7_75t_L g2987 ( 
.A(n_2534),
.B(n_1631),
.Y(n_2987)
);

NOR2xp33_ASAP7_75t_R g2988 ( 
.A(n_2461),
.B(n_1930),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2568),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2466),
.B(n_990),
.Y(n_2990)
);

NAND2xp33_ASAP7_75t_SL g2991 ( 
.A(n_2642),
.B(n_846),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2466),
.B(n_992),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2466),
.B(n_996),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2893),
.Y(n_2994)
);

BUFx12f_ASAP7_75t_L g2995 ( 
.A(n_2920),
.Y(n_2995)
);

AND2x4_ASAP7_75t_L g2996 ( 
.A(n_2722),
.B(n_2910),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2730),
.Y(n_2997)
);

BUFx3_ASAP7_75t_L g2998 ( 
.A(n_2759),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2730),
.Y(n_2999)
);

OAI21x1_ASAP7_75t_L g3000 ( 
.A1(n_2822),
.A2(n_1601),
.B(n_1587),
.Y(n_3000)
);

OAI21x1_ASAP7_75t_L g3001 ( 
.A1(n_2822),
.A2(n_1601),
.B(n_1587),
.Y(n_3001)
);

AOI22x1_ASAP7_75t_L g3002 ( 
.A1(n_2927),
.A2(n_1005),
.B1(n_1011),
.B2(n_1004),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_L g3003 ( 
.A(n_2765),
.B(n_846),
.Y(n_3003)
);

OAI21x1_ASAP7_75t_L g3004 ( 
.A1(n_2754),
.A2(n_1611),
.B(n_1603),
.Y(n_3004)
);

OAI21x1_ASAP7_75t_L g3005 ( 
.A1(n_2754),
.A2(n_1611),
.B(n_1603),
.Y(n_3005)
);

NAND2x1p5_ASAP7_75t_L g3006 ( 
.A(n_2940),
.B(n_1631),
.Y(n_3006)
);

BUFx2_ASAP7_75t_L g3007 ( 
.A(n_2759),
.Y(n_3007)
);

OAI21xp5_ASAP7_75t_L g3008 ( 
.A1(n_2894),
.A2(n_858),
.B(n_850),
.Y(n_3008)
);

AND2x4_ASAP7_75t_L g3009 ( 
.A(n_2722),
.B(n_571),
.Y(n_3009)
);

BUFx4_ASAP7_75t_SL g3010 ( 
.A(n_2817),
.Y(n_3010)
);

AND2x2_ASAP7_75t_L g3011 ( 
.A(n_2891),
.B(n_850),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2775),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2775),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2872),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2872),
.Y(n_3015)
);

BUFx6f_ASAP7_75t_L g3016 ( 
.A(n_2739),
.Y(n_3016)
);

BUFx10_ASAP7_75t_L g3017 ( 
.A(n_2732),
.Y(n_3017)
);

OAI21x1_ASAP7_75t_L g3018 ( 
.A1(n_2975),
.A2(n_1619),
.B(n_1612),
.Y(n_3018)
);

BUFx8_ASAP7_75t_L g3019 ( 
.A(n_2746),
.Y(n_3019)
);

AO21x2_ASAP7_75t_L g3020 ( 
.A1(n_2856),
.A2(n_864),
.B(n_859),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2771),
.Y(n_3021)
);

INVx3_ASAP7_75t_L g3022 ( 
.A(n_2735),
.Y(n_3022)
);

BUFx3_ASAP7_75t_L g3023 ( 
.A(n_2739),
.Y(n_3023)
);

OAI21x1_ASAP7_75t_L g3024 ( 
.A1(n_2975),
.A2(n_1619),
.B(n_1612),
.Y(n_3024)
);

AOI22x1_ASAP7_75t_L g3025 ( 
.A1(n_2939),
.A2(n_1014),
.B1(n_1016),
.B2(n_1012),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2893),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2773),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2717),
.B(n_1017),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2717),
.B(n_2731),
.Y(n_3029)
);

BUFx3_ASAP7_75t_L g3030 ( 
.A(n_2739),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2774),
.Y(n_3031)
);

INVx1_ASAP7_75t_SL g3032 ( 
.A(n_2786),
.Y(n_3032)
);

BUFx3_ASAP7_75t_L g3033 ( 
.A(n_2735),
.Y(n_3033)
);

BUFx6f_ASAP7_75t_L g3034 ( 
.A(n_2867),
.Y(n_3034)
);

OAI21x1_ASAP7_75t_L g3035 ( 
.A1(n_2979),
.A2(n_1639),
.B(n_1636),
.Y(n_3035)
);

BUFx6f_ASAP7_75t_L g3036 ( 
.A(n_2867),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2782),
.Y(n_3037)
);

HB1xp67_ASAP7_75t_L g3038 ( 
.A(n_2936),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2788),
.Y(n_3039)
);

OAI21xp5_ASAP7_75t_L g3040 ( 
.A1(n_2894),
.A2(n_864),
.B(n_859),
.Y(n_3040)
);

BUFx6f_ASAP7_75t_L g3041 ( 
.A(n_2867),
.Y(n_3041)
);

OAI21xp5_ASAP7_75t_L g3042 ( 
.A1(n_2781),
.A2(n_872),
.B(n_869),
.Y(n_3042)
);

OR2x6_ASAP7_75t_L g3043 ( 
.A(n_2795),
.B(n_1439),
.Y(n_3043)
);

OA21x2_ASAP7_75t_L g3044 ( 
.A1(n_2856),
.A2(n_1258),
.B(n_1257),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2936),
.Y(n_3045)
);

OAI21x1_ASAP7_75t_L g3046 ( 
.A1(n_2979),
.A2(n_1639),
.B(n_1636),
.Y(n_3046)
);

NAND2x1p5_ASAP7_75t_L g3047 ( 
.A(n_2940),
.B(n_1635),
.Y(n_3047)
);

BUFx8_ASAP7_75t_L g3048 ( 
.A(n_2762),
.Y(n_3048)
);

BUFx6f_ASAP7_75t_L g3049 ( 
.A(n_2867),
.Y(n_3049)
);

INVx2_ASAP7_75t_SL g3050 ( 
.A(n_2735),
.Y(n_3050)
);

BUFx3_ASAP7_75t_L g3051 ( 
.A(n_2830),
.Y(n_3051)
);

INVx3_ASAP7_75t_SL g3052 ( 
.A(n_2721),
.Y(n_3052)
);

BUFx12f_ASAP7_75t_L g3053 ( 
.A(n_2920),
.Y(n_3053)
);

OR2x6_ASAP7_75t_L g3054 ( 
.A(n_2795),
.B(n_1439),
.Y(n_3054)
);

BUFx3_ASAP7_75t_L g3055 ( 
.A(n_2756),
.Y(n_3055)
);

INVx1_ASAP7_75t_SL g3056 ( 
.A(n_2750),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2959),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2731),
.B(n_1018),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2959),
.Y(n_3059)
);

OAI21xp5_ASAP7_75t_L g3060 ( 
.A1(n_2781),
.A2(n_872),
.B(n_869),
.Y(n_3060)
);

OAI21x1_ASAP7_75t_L g3061 ( 
.A1(n_2713),
.A2(n_1635),
.B(n_1385),
.Y(n_3061)
);

INVx2_ASAP7_75t_SL g3062 ( 
.A(n_2767),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2820),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2869),
.Y(n_3064)
);

BUFx3_ASAP7_75t_L g3065 ( 
.A(n_2756),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2738),
.Y(n_3066)
);

INVx4_ASAP7_75t_L g3067 ( 
.A(n_2944),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2869),
.Y(n_3068)
);

BUFx2_ASAP7_75t_SL g3069 ( 
.A(n_2832),
.Y(n_3069)
);

NOR2xp33_ASAP7_75t_SL g3070 ( 
.A(n_2776),
.B(n_1022),
.Y(n_3070)
);

INVx3_ASAP7_75t_L g3071 ( 
.A(n_2944),
.Y(n_3071)
);

CKINVDCx14_ASAP7_75t_R g3072 ( 
.A(n_2988),
.Y(n_3072)
);

BUFx3_ASAP7_75t_L g3073 ( 
.A(n_2715),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2827),
.Y(n_3074)
);

NAND2x1p5_ASAP7_75t_L g3075 ( 
.A(n_2796),
.B(n_2892),
.Y(n_3075)
);

BUFx2_ASAP7_75t_SL g3076 ( 
.A(n_2757),
.Y(n_3076)
);

BUFx8_ASAP7_75t_L g3077 ( 
.A(n_2778),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2961),
.Y(n_3078)
);

BUFx3_ASAP7_75t_L g3079 ( 
.A(n_2715),
.Y(n_3079)
);

OAI21x1_ASAP7_75t_L g3080 ( 
.A1(n_2898),
.A2(n_1635),
.B(n_1389),
.Y(n_3080)
);

BUFx6f_ASAP7_75t_L g3081 ( 
.A(n_2876),
.Y(n_3081)
);

INVx1_ASAP7_75t_SL g3082 ( 
.A(n_2840),
.Y(n_3082)
);

INVx5_ASAP7_75t_L g3083 ( 
.A(n_2944),
.Y(n_3083)
);

OR2x2_ASAP7_75t_L g3084 ( 
.A(n_2737),
.B(n_877),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2827),
.Y(n_3085)
);

CKINVDCx5p33_ASAP7_75t_R g3086 ( 
.A(n_2988),
.Y(n_3086)
);

OA21x2_ASAP7_75t_L g3087 ( 
.A1(n_2764),
.A2(n_1258),
.B(n_1257),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2716),
.Y(n_3088)
);

AO21x2_ASAP7_75t_L g3089 ( 
.A1(n_2764),
.A2(n_879),
.B(n_877),
.Y(n_3089)
);

INVx5_ASAP7_75t_L g3090 ( 
.A(n_2954),
.Y(n_3090)
);

BUFx12f_ASAP7_75t_L g3091 ( 
.A(n_2866),
.Y(n_3091)
);

OR3x4_ASAP7_75t_SL g3092 ( 
.A(n_2732),
.B(n_885),
.C(n_1023),
.Y(n_3092)
);

OR2x6_ASAP7_75t_L g3093 ( 
.A(n_2795),
.B(n_879),
.Y(n_3093)
);

AOI21xp5_ASAP7_75t_L g3094 ( 
.A1(n_2726),
.A2(n_2718),
.B(n_2789),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_2761),
.B(n_883),
.Y(n_3095)
);

INVx5_ASAP7_75t_L g3096 ( 
.A(n_2954),
.Y(n_3096)
);

BUFx2_ASAP7_75t_L g3097 ( 
.A(n_2742),
.Y(n_3097)
);

AOI22x1_ASAP7_75t_L g3098 ( 
.A1(n_2949),
.A2(n_2882),
.B1(n_2780),
.B2(n_2826),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2729),
.Y(n_3099)
);

BUFx3_ASAP7_75t_L g3100 ( 
.A(n_2742),
.Y(n_3100)
);

BUFx6f_ASAP7_75t_L g3101 ( 
.A(n_2876),
.Y(n_3101)
);

CKINVDCx5p33_ASAP7_75t_R g3102 ( 
.A(n_2745),
.Y(n_3102)
);

NAND2x1p5_ASAP7_75t_L g3103 ( 
.A(n_2766),
.B(n_1564),
.Y(n_3103)
);

BUFx12f_ASAP7_75t_L g3104 ( 
.A(n_2884),
.Y(n_3104)
);

BUFx6f_ASAP7_75t_L g3105 ( 
.A(n_2876),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2961),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2898),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2744),
.Y(n_3108)
);

AOI22x1_ASAP7_75t_L g3109 ( 
.A1(n_2969),
.A2(n_1033),
.B1(n_1034),
.B2(n_1029),
.Y(n_3109)
);

CKINVDCx6p67_ASAP7_75t_R g3110 ( 
.A(n_2814),
.Y(n_3110)
);

AOI21x1_ASAP7_75t_L g3111 ( 
.A1(n_2889),
.A2(n_1261),
.B(n_1260),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2753),
.Y(n_3112)
);

AO21x2_ASAP7_75t_L g3113 ( 
.A1(n_2924),
.A2(n_2889),
.B(n_2768),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2799),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2912),
.Y(n_3115)
);

INVx2_ASAP7_75t_SL g3116 ( 
.A(n_2767),
.Y(n_3116)
);

BUFx3_ASAP7_75t_L g3117 ( 
.A(n_2876),
.Y(n_3117)
);

OR2x2_ASAP7_75t_L g3118 ( 
.A(n_2896),
.B(n_883),
.Y(n_3118)
);

BUFx2_ASAP7_75t_SL g3119 ( 
.A(n_2728),
.Y(n_3119)
);

BUFx2_ASAP7_75t_R g3120 ( 
.A(n_2880),
.Y(n_3120)
);

BUFx3_ASAP7_75t_L g3121 ( 
.A(n_2841),
.Y(n_3121)
);

BUFx6f_ASAP7_75t_L g3122 ( 
.A(n_2836),
.Y(n_3122)
);

CKINVDCx11_ASAP7_75t_R g3123 ( 
.A(n_2978),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2752),
.B(n_1036),
.Y(n_3124)
);

AND2x2_ASAP7_75t_L g3125 ( 
.A(n_2720),
.B(n_895),
.Y(n_3125)
);

OAI21x1_ASAP7_75t_L g3126 ( 
.A1(n_2899),
.A2(n_1399),
.B(n_1373),
.Y(n_3126)
);

OA21x2_ASAP7_75t_L g3127 ( 
.A1(n_2765),
.A2(n_1261),
.B(n_1260),
.Y(n_3127)
);

INVx1_ASAP7_75t_SL g3128 ( 
.A(n_2905),
.Y(n_3128)
);

HB1xp67_ASAP7_75t_L g3129 ( 
.A(n_2899),
.Y(n_3129)
);

BUFx6f_ASAP7_75t_L g3130 ( 
.A(n_2836),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2896),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2955),
.Y(n_3132)
);

AO21x2_ASAP7_75t_L g3133 ( 
.A1(n_2924),
.A2(n_901),
.B(n_895),
.Y(n_3133)
);

BUFx4_ASAP7_75t_SL g3134 ( 
.A(n_2906),
.Y(n_3134)
);

AND2x4_ASAP7_75t_L g3135 ( 
.A(n_2910),
.B(n_572),
.Y(n_3135)
);

AND2x4_ASAP7_75t_L g3136 ( 
.A(n_2913),
.B(n_573),
.Y(n_3136)
);

INVx4_ASAP7_75t_L g3137 ( 
.A(n_2954),
.Y(n_3137)
);

AOI22x1_ASAP7_75t_L g3138 ( 
.A1(n_2857),
.A2(n_1040),
.B1(n_1041),
.B2(n_1038),
.Y(n_3138)
);

AOI22x1_ASAP7_75t_L g3139 ( 
.A1(n_2881),
.A2(n_1050),
.B1(n_1054),
.B2(n_1044),
.Y(n_3139)
);

OAI21x1_ASAP7_75t_L g3140 ( 
.A1(n_2874),
.A2(n_1399),
.B(n_1308),
.Y(n_3140)
);

AO21x2_ASAP7_75t_L g3141 ( 
.A1(n_2874),
.A2(n_906),
.B(n_901),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2752),
.B(n_2760),
.Y(n_3142)
);

INVx1_ASAP7_75t_SL g3143 ( 
.A(n_2981),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_2847),
.Y(n_3144)
);

OA21x2_ASAP7_75t_L g3145 ( 
.A1(n_2816),
.A2(n_2766),
.B(n_2904),
.Y(n_3145)
);

INVx3_ASAP7_75t_L g3146 ( 
.A(n_2740),
.Y(n_3146)
);

OAI21x1_ASAP7_75t_L g3147 ( 
.A1(n_2798),
.A2(n_1308),
.B(n_1325),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2760),
.B(n_1057),
.Y(n_3148)
);

OAI21xp5_ASAP7_75t_L g3149 ( 
.A1(n_2851),
.A2(n_908),
.B(n_906),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2819),
.Y(n_3150)
);

BUFx2_ASAP7_75t_SL g3151 ( 
.A(n_2736),
.Y(n_3151)
);

BUFx3_ASAP7_75t_L g3152 ( 
.A(n_2841),
.Y(n_3152)
);

BUFx12f_ASAP7_75t_L g3153 ( 
.A(n_2938),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_2847),
.Y(n_3154)
);

OAI21x1_ASAP7_75t_L g3155 ( 
.A1(n_2798),
.A2(n_1357),
.B(n_1325),
.Y(n_3155)
);

BUFx8_ASAP7_75t_L g3156 ( 
.A(n_2846),
.Y(n_3156)
);

BUFx3_ASAP7_75t_L g3157 ( 
.A(n_2848),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2724),
.Y(n_3158)
);

HB1xp67_ASAP7_75t_L g3159 ( 
.A(n_2853),
.Y(n_3159)
);

BUFx3_ASAP7_75t_L g3160 ( 
.A(n_2848),
.Y(n_3160)
);

OAI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_2851),
.A2(n_909),
.B(n_908),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2845),
.Y(n_3162)
);

OAI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2883),
.A2(n_910),
.B(n_909),
.Y(n_3163)
);

NAND2x1p5_ASAP7_75t_L g3164 ( 
.A(n_2953),
.B(n_1564),
.Y(n_3164)
);

OAI21x1_ASAP7_75t_L g3165 ( 
.A1(n_2853),
.A2(n_1357),
.B(n_1325),
.Y(n_3165)
);

BUFx2_ASAP7_75t_SL g3166 ( 
.A(n_2741),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2763),
.Y(n_3167)
);

BUFx6f_ASAP7_75t_L g3168 ( 
.A(n_2836),
.Y(n_3168)
);

BUFx3_ASAP7_75t_L g3169 ( 
.A(n_2749),
.Y(n_3169)
);

CKINVDCx6p67_ASAP7_75t_R g3170 ( 
.A(n_2953),
.Y(n_3170)
);

INVx1_ASAP7_75t_SL g3171 ( 
.A(n_2748),
.Y(n_3171)
);

BUFx3_ASAP7_75t_L g3172 ( 
.A(n_2749),
.Y(n_3172)
);

INVx4_ASAP7_75t_L g3173 ( 
.A(n_2740),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2763),
.Y(n_3174)
);

OAI21x1_ASAP7_75t_L g3175 ( 
.A1(n_2793),
.A2(n_2850),
.B(n_2797),
.Y(n_3175)
);

INVx1_ASAP7_75t_SL g3176 ( 
.A(n_2770),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_2913),
.Y(n_3177)
);

AO21x2_ASAP7_75t_L g3178 ( 
.A1(n_2755),
.A2(n_913),
.B(n_911),
.Y(n_3178)
);

AO21x2_ASAP7_75t_L g3179 ( 
.A1(n_2755),
.A2(n_2865),
.B(n_2811),
.Y(n_3179)
);

BUFx3_ASAP7_75t_L g3180 ( 
.A(n_2836),
.Y(n_3180)
);

BUFx6f_ASAP7_75t_L g3181 ( 
.A(n_2801),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2797),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2849),
.Y(n_3183)
);

OAI21x1_ASAP7_75t_L g3184 ( 
.A1(n_2904),
.A2(n_2800),
.B(n_2815),
.Y(n_3184)
);

OAI21xp5_ASAP7_75t_L g3185 ( 
.A1(n_2883),
.A2(n_913),
.B(n_911),
.Y(n_3185)
);

BUFx2_ASAP7_75t_L g3186 ( 
.A(n_2777),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2733),
.B(n_1058),
.Y(n_3187)
);

INVx1_ASAP7_75t_SL g3188 ( 
.A(n_2823),
.Y(n_3188)
);

NOR2xp33_ASAP7_75t_L g3189 ( 
.A(n_2861),
.B(n_914),
.Y(n_3189)
);

AO21x2_ASAP7_75t_L g3190 ( 
.A1(n_2865),
.A2(n_918),
.B(n_914),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_2861),
.B(n_2790),
.Y(n_3191)
);

CKINVDCx6p67_ASAP7_75t_R g3192 ( 
.A(n_2808),
.Y(n_3192)
);

BUFx2_ASAP7_75t_R g3193 ( 
.A(n_2973),
.Y(n_3193)
);

AOI22xp33_ASAP7_75t_L g3194 ( 
.A1(n_2991),
.A2(n_918),
.B1(n_924),
.B2(n_923),
.Y(n_3194)
);

AND2x2_ASAP7_75t_L g3195 ( 
.A(n_2802),
.B(n_923),
.Y(n_3195)
);

OAI21xp5_ASAP7_75t_L g3196 ( 
.A1(n_2960),
.A2(n_2863),
.B(n_2983),
.Y(n_3196)
);

OAI21x1_ASAP7_75t_L g3197 ( 
.A1(n_2815),
.A2(n_1357),
.B(n_1085),
.Y(n_3197)
);

AOI22x1_ASAP7_75t_L g3198 ( 
.A1(n_2930),
.A2(n_924),
.B1(n_936),
.B2(n_933),
.Y(n_3198)
);

OAI21xp5_ASAP7_75t_L g3199 ( 
.A1(n_2960),
.A2(n_936),
.B(n_933),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2785),
.B(n_942),
.Y(n_3200)
);

OR2x6_ASAP7_75t_L g3201 ( 
.A(n_2801),
.B(n_942),
.Y(n_3201)
);

OR2x6_ASAP7_75t_L g3202 ( 
.A(n_2801),
.B(n_959),
.Y(n_3202)
);

BUFx8_ASAP7_75t_L g3203 ( 
.A(n_2809),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2951),
.Y(n_3204)
);

INVx4_ASAP7_75t_L g3205 ( 
.A(n_2784),
.Y(n_3205)
);

INVx2_ASAP7_75t_SL g3206 ( 
.A(n_2828),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2946),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2852),
.Y(n_3208)
);

OAI21x1_ASAP7_75t_L g3209 ( 
.A1(n_2835),
.A2(n_1085),
.B(n_1081),
.Y(n_3209)
);

INVx3_ASAP7_75t_L g3210 ( 
.A(n_2801),
.Y(n_3210)
);

OAI21x1_ASAP7_75t_L g3211 ( 
.A1(n_2835),
.A2(n_1087),
.B(n_1086),
.Y(n_3211)
);

AOI22x1_ASAP7_75t_L g3212 ( 
.A1(n_2950),
.A2(n_959),
.B1(n_971),
.B2(n_963),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_2844),
.Y(n_3213)
);

BUFx4f_ASAP7_75t_SL g3214 ( 
.A(n_2784),
.Y(n_3214)
);

BUFx12f_ASAP7_75t_L g3215 ( 
.A(n_2813),
.Y(n_3215)
);

AO21x2_ASAP7_75t_L g3216 ( 
.A1(n_2868),
.A2(n_971),
.B(n_963),
.Y(n_3216)
);

AND2x2_ASAP7_75t_L g3217 ( 
.A(n_2805),
.B(n_2947),
.Y(n_3217)
);

AOI22x1_ASAP7_75t_L g3218 ( 
.A1(n_2929),
.A2(n_972),
.B1(n_981),
.B2(n_977),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2859),
.Y(n_3219)
);

OAI21x1_ASAP7_75t_L g3220 ( 
.A1(n_2838),
.A2(n_1087),
.B(n_1086),
.Y(n_3220)
);

OAI21x1_ASAP7_75t_L g3221 ( 
.A1(n_2838),
.A2(n_1095),
.B(n_1091),
.Y(n_3221)
);

AND2x4_ASAP7_75t_L g3222 ( 
.A(n_2791),
.B(n_576),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2862),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2877),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2886),
.Y(n_3225)
);

OAI21x1_ASAP7_75t_L g3226 ( 
.A1(n_2794),
.A2(n_2834),
.B(n_2821),
.Y(n_3226)
);

HB1xp67_ASAP7_75t_L g3227 ( 
.A(n_2816),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2890),
.Y(n_3228)
);

AND2x2_ASAP7_75t_L g3229 ( 
.A(n_2923),
.B(n_972),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_2844),
.Y(n_3230)
);

AO21x2_ASAP7_75t_L g3231 ( 
.A1(n_2868),
.A2(n_981),
.B(n_977),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2860),
.Y(n_3232)
);

CKINVDCx5p33_ASAP7_75t_R g3233 ( 
.A(n_2933),
.Y(n_3233)
);

INVxp67_ASAP7_75t_SL g3234 ( 
.A(n_2860),
.Y(n_3234)
);

BUFx6f_ASAP7_75t_L g3235 ( 
.A(n_2829),
.Y(n_3235)
);

AO21x2_ASAP7_75t_L g3236 ( 
.A1(n_2783),
.A2(n_983),
.B(n_982),
.Y(n_3236)
);

BUFx6f_ASAP7_75t_L g3237 ( 
.A(n_2829),
.Y(n_3237)
);

BUFx2_ASAP7_75t_L g3238 ( 
.A(n_2777),
.Y(n_3238)
);

BUFx6f_ASAP7_75t_L g3239 ( 
.A(n_2829),
.Y(n_3239)
);

BUFx2_ASAP7_75t_SL g3240 ( 
.A(n_2854),
.Y(n_3240)
);

NAND2x1p5_ASAP7_75t_L g3241 ( 
.A(n_2787),
.B(n_1569),
.Y(n_3241)
);

BUFx4f_ASAP7_75t_L g3242 ( 
.A(n_2829),
.Y(n_3242)
);

BUFx6f_ASAP7_75t_L g3243 ( 
.A(n_2828),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2908),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2911),
.Y(n_3245)
);

INVx1_ASAP7_75t_SL g3246 ( 
.A(n_2823),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2725),
.Y(n_3247)
);

BUFx6f_ASAP7_75t_L g3248 ( 
.A(n_2787),
.Y(n_3248)
);

INVx4_ASAP7_75t_SL g3249 ( 
.A(n_2791),
.Y(n_3249)
);

OAI21x1_ASAP7_75t_L g3250 ( 
.A1(n_2821),
.A2(n_1095),
.B(n_1091),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_2714),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_SL g3252 ( 
.A(n_2723),
.B(n_982),
.Y(n_3252)
);

BUFx3_ASAP7_75t_L g3253 ( 
.A(n_2743),
.Y(n_3253)
);

BUFx12f_ASAP7_75t_L g3254 ( 
.A(n_2818),
.Y(n_3254)
);

OAI21x1_ASAP7_75t_L g3255 ( 
.A1(n_2834),
.A2(n_1097),
.B(n_1096),
.Y(n_3255)
);

AOI22xp5_ASAP7_75t_L g3256 ( 
.A1(n_2916),
.A2(n_2712),
.B1(n_2933),
.B2(n_2991),
.Y(n_3256)
);

INVx2_ASAP7_75t_SL g3257 ( 
.A(n_2743),
.Y(n_3257)
);

INVx1_ASAP7_75t_SL g3258 ( 
.A(n_2941),
.Y(n_3258)
);

OAI21xp5_ASAP7_75t_L g3259 ( 
.A1(n_2863),
.A2(n_984),
.B(n_983),
.Y(n_3259)
);

INVx1_ASAP7_75t_SL g3260 ( 
.A(n_2928),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_2719),
.B(n_984),
.Y(n_3261)
);

BUFx3_ASAP7_75t_L g3262 ( 
.A(n_2806),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_2714),
.Y(n_3263)
);

BUFx4f_ASAP7_75t_L g3264 ( 
.A(n_2806),
.Y(n_3264)
);

BUFx3_ASAP7_75t_L g3265 ( 
.A(n_2987),
.Y(n_3265)
);

BUFx4f_ASAP7_75t_L g3266 ( 
.A(n_2987),
.Y(n_3266)
);

OA21x2_ASAP7_75t_L g3267 ( 
.A1(n_2965),
.A2(n_2966),
.B(n_2803),
.Y(n_3267)
);

OAI21x1_ASAP7_75t_L g3268 ( 
.A1(n_2919),
.A2(n_1097),
.B(n_1096),
.Y(n_3268)
);

OAI21x1_ASAP7_75t_L g3269 ( 
.A1(n_2783),
.A2(n_993),
.B(n_991),
.Y(n_3269)
);

AOI22xp33_ASAP7_75t_L g3270 ( 
.A1(n_2878),
.A2(n_991),
.B1(n_995),
.B2(n_993),
.Y(n_3270)
);

AND2x4_ASAP7_75t_L g3271 ( 
.A(n_2734),
.B(n_579),
.Y(n_3271)
);

OA21x2_ASAP7_75t_L g3272 ( 
.A1(n_2965),
.A2(n_997),
.B(n_995),
.Y(n_3272)
);

OAI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_2984),
.A2(n_1001),
.B(n_997),
.Y(n_3273)
);

AOI22x1_ASAP7_75t_L g3274 ( 
.A1(n_2792),
.A2(n_1001),
.B1(n_1015),
.B2(n_1007),
.Y(n_3274)
);

BUFx3_ASAP7_75t_L g3275 ( 
.A(n_2902),
.Y(n_3275)
);

OAI21xp5_ASAP7_75t_L g3276 ( 
.A1(n_2990),
.A2(n_1015),
.B(n_1007),
.Y(n_3276)
);

BUFx2_ASAP7_75t_SL g3277 ( 
.A(n_2952),
.Y(n_3277)
);

CKINVDCx20_ASAP7_75t_R g3278 ( 
.A(n_3123),
.Y(n_3278)
);

AOI22xp33_ASAP7_75t_SL g3279 ( 
.A1(n_3196),
.A2(n_2909),
.B1(n_2864),
.B2(n_2875),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_3114),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3038),
.Y(n_3281)
);

INVx6_ASAP7_75t_L g3282 ( 
.A(n_3090),
.Y(n_3282)
);

AOI22xp5_ASAP7_75t_L g3283 ( 
.A1(n_3256),
.A2(n_2727),
.B1(n_2870),
.B2(n_2957),
.Y(n_3283)
);

AOI22xp33_ASAP7_75t_L g3284 ( 
.A1(n_3199),
.A2(n_2871),
.B1(n_2931),
.B2(n_2903),
.Y(n_3284)
);

OAI22xp5_ASAP7_75t_L g3285 ( 
.A1(n_3163),
.A2(n_2966),
.B1(n_2804),
.B2(n_2769),
.Y(n_3285)
);

INVx2_ASAP7_75t_SL g3286 ( 
.A(n_3134),
.Y(n_3286)
);

BUFx6f_ASAP7_75t_L g3287 ( 
.A(n_3090),
.Y(n_3287)
);

INVx11_ASAP7_75t_L g3288 ( 
.A(n_3019),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3038),
.Y(n_3289)
);

CKINVDCx11_ASAP7_75t_R g3290 ( 
.A(n_3123),
.Y(n_3290)
);

BUFx12f_ASAP7_75t_L g3291 ( 
.A(n_3086),
.Y(n_3291)
);

OAI22xp33_ASAP7_75t_L g3292 ( 
.A1(n_3192),
.A2(n_2758),
.B1(n_2934),
.B2(n_2843),
.Y(n_3292)
);

NAND2x1p5_ASAP7_75t_L g3293 ( 
.A(n_3090),
.B(n_2971),
.Y(n_3293)
);

AOI22xp33_ASAP7_75t_SL g3294 ( 
.A1(n_3185),
.A2(n_3189),
.B1(n_3040),
.B2(n_3008),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_2997),
.Y(n_3295)
);

AOI22xp33_ASAP7_75t_L g3296 ( 
.A1(n_3189),
.A2(n_2914),
.B1(n_2888),
.B2(n_2901),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2999),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3012),
.Y(n_3298)
);

INVx6_ASAP7_75t_L g3299 ( 
.A(n_3019),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3013),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3014),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3015),
.Y(n_3302)
);

BUFx6f_ASAP7_75t_L g3303 ( 
.A(n_3090),
.Y(n_3303)
);

AOI22xp33_ASAP7_75t_L g3304 ( 
.A1(n_3149),
.A2(n_2873),
.B1(n_2831),
.B2(n_2837),
.Y(n_3304)
);

AOI22xp33_ASAP7_75t_L g3305 ( 
.A1(n_3161),
.A2(n_2917),
.B1(n_2921),
.B2(n_2918),
.Y(n_3305)
);

AOI22xp33_ASAP7_75t_L g3306 ( 
.A1(n_3153),
.A2(n_2932),
.B1(n_2935),
.B2(n_2942),
.Y(n_3306)
);

INVx3_ASAP7_75t_L g3307 ( 
.A(n_3122),
.Y(n_3307)
);

CKINVDCx11_ASAP7_75t_R g3308 ( 
.A(n_3052),
.Y(n_3308)
);

INVx6_ASAP7_75t_L g3309 ( 
.A(n_3096),
.Y(n_3309)
);

INVx6_ASAP7_75t_L g3310 ( 
.A(n_3096),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3074),
.Y(n_3311)
);

AOI22xp33_ASAP7_75t_L g3312 ( 
.A1(n_3153),
.A2(n_2956),
.B1(n_2968),
.B2(n_2879),
.Y(n_3312)
);

AOI22xp33_ASAP7_75t_L g3313 ( 
.A1(n_3098),
.A2(n_2915),
.B1(n_2833),
.B2(n_2839),
.Y(n_3313)
);

AOI22xp33_ASAP7_75t_L g3314 ( 
.A1(n_3093),
.A2(n_2855),
.B1(n_2887),
.B2(n_2885),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3162),
.Y(n_3315)
);

CKINVDCx5p33_ASAP7_75t_R g3316 ( 
.A(n_3134),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_3063),
.Y(n_3317)
);

INVx6_ASAP7_75t_L g3318 ( 
.A(n_3019),
.Y(n_3318)
);

AOI22xp33_ASAP7_75t_L g3319 ( 
.A1(n_3093),
.A2(n_2895),
.B1(n_2900),
.B2(n_2897),
.Y(n_3319)
);

AOI22xp33_ASAP7_75t_L g3320 ( 
.A1(n_3093),
.A2(n_2963),
.B1(n_2907),
.B2(n_2824),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3085),
.Y(n_3321)
);

INVx1_ASAP7_75t_SL g3322 ( 
.A(n_3258),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_3066),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_3115),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3129),
.Y(n_3325)
);

INVx1_ASAP7_75t_SL g3326 ( 
.A(n_3171),
.Y(n_3326)
);

OAI22xp5_ASAP7_75t_L g3327 ( 
.A1(n_3194),
.A2(n_2772),
.B1(n_2751),
.B2(n_2810),
.Y(n_3327)
);

AOI22xp33_ASAP7_75t_L g3328 ( 
.A1(n_3191),
.A2(n_3215),
.B1(n_3254),
.B2(n_3119),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3129),
.Y(n_3329)
);

CKINVDCx20_ASAP7_75t_R g3330 ( 
.A(n_3072),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3088),
.Y(n_3331)
);

INVx6_ASAP7_75t_L g3332 ( 
.A(n_3096),
.Y(n_3332)
);

AOI22xp33_ASAP7_75t_L g3333 ( 
.A1(n_3191),
.A2(n_2948),
.B1(n_1020),
.B2(n_1031),
.Y(n_3333)
);

BUFx12f_ASAP7_75t_L g3334 ( 
.A(n_3086),
.Y(n_3334)
);

AOI22xp33_ASAP7_75t_SL g3335 ( 
.A1(n_3003),
.A2(n_2986),
.B1(n_2727),
.B2(n_2825),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_3183),
.Y(n_3336)
);

AOI22xp33_ASAP7_75t_L g3337 ( 
.A1(n_3215),
.A2(n_1020),
.B1(n_1031),
.B2(n_1028),
.Y(n_3337)
);

INVx4_ASAP7_75t_L g3338 ( 
.A(n_3096),
.Y(n_3338)
);

BUFx3_ASAP7_75t_L g3339 ( 
.A(n_2998),
.Y(n_3339)
);

OAI22xp5_ASAP7_75t_L g3340 ( 
.A1(n_3194),
.A2(n_2810),
.B1(n_2747),
.B2(n_2992),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3099),
.Y(n_3341)
);

AOI22xp33_ASAP7_75t_SL g3342 ( 
.A1(n_3003),
.A2(n_2807),
.B1(n_2937),
.B2(n_2842),
.Y(n_3342)
);

INVx4_ASAP7_75t_L g3343 ( 
.A(n_3083),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_2994),
.Y(n_3344)
);

AOI22xp5_ASAP7_75t_L g3345 ( 
.A1(n_3254),
.A2(n_2870),
.B1(n_2964),
.B2(n_2993),
.Y(n_3345)
);

INVx4_ASAP7_75t_L g3346 ( 
.A(n_3083),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_L g3347 ( 
.A1(n_3151),
.A2(n_1028),
.B1(n_1045),
.B2(n_1042),
.Y(n_3347)
);

INVx1_ASAP7_75t_SL g3348 ( 
.A(n_3227),
.Y(n_3348)
);

CKINVDCx11_ASAP7_75t_R g3349 ( 
.A(n_3052),
.Y(n_3349)
);

BUFx8_ASAP7_75t_L g3350 ( 
.A(n_2995),
.Y(n_3350)
);

INVx2_ASAP7_75t_SL g3351 ( 
.A(n_2998),
.Y(n_3351)
);

BUFx6f_ASAP7_75t_L g3352 ( 
.A(n_3137),
.Y(n_3352)
);

AOI22xp33_ASAP7_75t_L g3353 ( 
.A1(n_3166),
.A2(n_3276),
.B1(n_3273),
.B2(n_3277),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2994),
.Y(n_3354)
);

INVx6_ASAP7_75t_L g3355 ( 
.A(n_3137),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3026),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3026),
.Y(n_3357)
);

INVx6_ASAP7_75t_L g3358 ( 
.A(n_3048),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_SL g3359 ( 
.A1(n_3203),
.A2(n_1042),
.B1(n_1047),
.B2(n_1046),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3208),
.Y(n_3360)
);

CKINVDCx5p33_ASAP7_75t_R g3361 ( 
.A(n_3010),
.Y(n_3361)
);

CKINVDCx11_ASAP7_75t_R g3362 ( 
.A(n_2995),
.Y(n_3362)
);

OAI22xp5_ASAP7_75t_L g3363 ( 
.A1(n_3143),
.A2(n_2925),
.B1(n_2985),
.B2(n_2982),
.Y(n_3363)
);

AOI22xp33_ASAP7_75t_SL g3364 ( 
.A1(n_3203),
.A2(n_1047),
.B1(n_2943),
.B2(n_2922),
.Y(n_3364)
);

INVx3_ASAP7_75t_L g3365 ( 
.A(n_3122),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_3150),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_3132),
.Y(n_3367)
);

AOI22xp33_ASAP7_75t_L g3368 ( 
.A1(n_3043),
.A2(n_2976),
.B1(n_2967),
.B2(n_2958),
.Y(n_3368)
);

BUFx3_ASAP7_75t_L g3369 ( 
.A(n_3091),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3219),
.Y(n_3370)
);

CKINVDCx5p33_ASAP7_75t_R g3371 ( 
.A(n_3010),
.Y(n_3371)
);

BUFx3_ASAP7_75t_L g3372 ( 
.A(n_3091),
.Y(n_3372)
);

BUFx2_ASAP7_75t_L g3373 ( 
.A(n_3051),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_3021),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_SL g3375 ( 
.A1(n_3203),
.A2(n_2982),
.B1(n_2989),
.B2(n_2985),
.Y(n_3375)
);

BUFx2_ASAP7_75t_L g3376 ( 
.A(n_3051),
.Y(n_3376)
);

CKINVDCx20_ASAP7_75t_R g3377 ( 
.A(n_3072),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3223),
.Y(n_3378)
);

AOI22xp33_ASAP7_75t_SL g3379 ( 
.A1(n_3020),
.A2(n_2989),
.B1(n_2926),
.B2(n_2972),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3224),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3225),
.Y(n_3381)
);

AOI22xp5_ASAP7_75t_SL g3382 ( 
.A1(n_3055),
.A2(n_2925),
.B1(n_2962),
.B2(n_2974),
.Y(n_3382)
);

BUFx3_ASAP7_75t_L g3383 ( 
.A(n_3055),
.Y(n_3383)
);

AOI22xp33_ASAP7_75t_SL g3384 ( 
.A1(n_3020),
.A2(n_3042),
.B1(n_3060),
.B2(n_3274),
.Y(n_3384)
);

OAI22xp5_ASAP7_75t_L g3385 ( 
.A1(n_3176),
.A2(n_2779),
.B1(n_2945),
.B2(n_2977),
.Y(n_3385)
);

CKINVDCx11_ASAP7_75t_R g3386 ( 
.A(n_3053),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3228),
.Y(n_3387)
);

AOI22xp33_ASAP7_75t_L g3388 ( 
.A1(n_3043),
.A2(n_2858),
.B1(n_2970),
.B2(n_2980),
.Y(n_3388)
);

BUFx2_ASAP7_75t_L g3389 ( 
.A(n_3156),
.Y(n_3389)
);

BUFx8_ASAP7_75t_SL g3390 ( 
.A(n_3007),
.Y(n_3390)
);

AOI22xp33_ASAP7_75t_L g3391 ( 
.A1(n_3043),
.A2(n_2858),
.B1(n_2980),
.B2(n_2902),
.Y(n_3391)
);

INVxp67_ASAP7_75t_SL g3392 ( 
.A(n_3234),
.Y(n_3392)
);

AOI22xp33_ASAP7_75t_L g3393 ( 
.A1(n_3054),
.A2(n_2812),
.B1(n_1382),
.B2(n_1415),
.Y(n_3393)
);

AOI22xp33_ASAP7_75t_L g3394 ( 
.A1(n_3054),
.A2(n_2812),
.B1(n_1382),
.B2(n_1415),
.Y(n_3394)
);

BUFx4_ASAP7_75t_SL g3395 ( 
.A(n_3065),
.Y(n_3395)
);

INVx1_ASAP7_75t_SL g3396 ( 
.A(n_3227),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3244),
.Y(n_3397)
);

INVx2_ASAP7_75t_L g3398 ( 
.A(n_3027),
.Y(n_3398)
);

CKINVDCx11_ASAP7_75t_R g3399 ( 
.A(n_3053),
.Y(n_3399)
);

INVx8_ASAP7_75t_L g3400 ( 
.A(n_3083),
.Y(n_3400)
);

OAI22xp5_ASAP7_75t_L g3401 ( 
.A1(n_3233),
.A2(n_885),
.B1(n_3),
.B2(n_1),
.Y(n_3401)
);

BUFx10_ASAP7_75t_L g3402 ( 
.A(n_3102),
.Y(n_3402)
);

BUFx2_ASAP7_75t_SL g3403 ( 
.A(n_3065),
.Y(n_3403)
);

BUFx6f_ASAP7_75t_L g3404 ( 
.A(n_3034),
.Y(n_3404)
);

BUFx4f_ASAP7_75t_SL g3405 ( 
.A(n_3104),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3245),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3234),
.B(n_3094),
.Y(n_3407)
);

AOI22xp33_ASAP7_75t_SL g3408 ( 
.A1(n_3156),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_3408)
);

CKINVDCx11_ASAP7_75t_R g3409 ( 
.A(n_3104),
.Y(n_3409)
);

NAND2x1p5_ASAP7_75t_L g3410 ( 
.A(n_3083),
.B(n_1330),
.Y(n_3410)
);

CKINVDCx5p33_ASAP7_75t_R g3411 ( 
.A(n_3102),
.Y(n_3411)
);

OAI21xp33_ASAP7_75t_L g3412 ( 
.A1(n_3270),
.A2(n_1413),
.B(n_1382),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3078),
.Y(n_3413)
);

OAI21xp5_ASAP7_75t_SL g3414 ( 
.A1(n_3270),
.A2(n_2),
.B(n_6),
.Y(n_3414)
);

CKINVDCx11_ASAP7_75t_R g3415 ( 
.A(n_3017),
.Y(n_3415)
);

CKINVDCx11_ASAP7_75t_R g3416 ( 
.A(n_3017),
.Y(n_3416)
);

AOI22xp33_ASAP7_75t_L g3417 ( 
.A1(n_3054),
.A2(n_1413),
.B1(n_1415),
.B2(n_1382),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3078),
.Y(n_3418)
);

CKINVDCx5p33_ASAP7_75t_R g3419 ( 
.A(n_3076),
.Y(n_3419)
);

BUFx2_ASAP7_75t_SL g3420 ( 
.A(n_3082),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3106),
.Y(n_3421)
);

INVx4_ASAP7_75t_L g3422 ( 
.A(n_3170),
.Y(n_3422)
);

AOI22xp33_ASAP7_75t_L g3423 ( 
.A1(n_3011),
.A2(n_1415),
.B1(n_1422),
.B2(n_1413),
.Y(n_3423)
);

AOI22xp5_ASAP7_75t_L g3424 ( 
.A1(n_3260),
.A2(n_1415),
.B1(n_1422),
.B2(n_1413),
.Y(n_3424)
);

AOI22xp33_ASAP7_75t_L g3425 ( 
.A1(n_3233),
.A2(n_1426),
.B1(n_1429),
.B2(n_1422),
.Y(n_3425)
);

OAI21xp5_ASAP7_75t_SL g3426 ( 
.A1(n_3259),
.A2(n_7),
.B(n_8),
.Y(n_3426)
);

AND2x2_ASAP7_75t_L g3427 ( 
.A(n_2996),
.B(n_3247),
.Y(n_3427)
);

BUFx2_ASAP7_75t_L g3428 ( 
.A(n_3156),
.Y(n_3428)
);

CKINVDCx11_ASAP7_75t_R g3429 ( 
.A(n_3110),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3106),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3031),
.Y(n_3431)
);

AOI22xp33_ASAP7_75t_L g3432 ( 
.A1(n_2996),
.A2(n_1426),
.B1(n_1429),
.B2(n_1422),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3107),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3107),
.Y(n_3434)
);

CKINVDCx11_ASAP7_75t_R g3435 ( 
.A(n_3128),
.Y(n_3435)
);

HB1xp67_ASAP7_75t_L g3436 ( 
.A(n_3075),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_3037),
.Y(n_3437)
);

BUFx3_ASAP7_75t_L g3438 ( 
.A(n_3048),
.Y(n_3438)
);

OAI22xp33_ASAP7_75t_L g3439 ( 
.A1(n_3070),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_3439)
);

AOI22xp33_ASAP7_75t_L g3440 ( 
.A1(n_2996),
.A2(n_1426),
.B1(n_1429),
.B2(n_1422),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3045),
.Y(n_3441)
);

INVx2_ASAP7_75t_L g3442 ( 
.A(n_3039),
.Y(n_3442)
);

BUFx2_ASAP7_75t_L g3443 ( 
.A(n_3121),
.Y(n_3443)
);

AOI22xp33_ASAP7_75t_L g3444 ( 
.A1(n_3217),
.A2(n_1429),
.B1(n_1438),
.B2(n_1426),
.Y(n_3444)
);

INVx2_ASAP7_75t_SL g3445 ( 
.A(n_3048),
.Y(n_3445)
);

BUFx6f_ASAP7_75t_SL g3446 ( 
.A(n_3009),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3057),
.Y(n_3447)
);

BUFx6f_ASAP7_75t_L g3448 ( 
.A(n_3034),
.Y(n_3448)
);

INVx3_ASAP7_75t_L g3449 ( 
.A(n_3122),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3108),
.Y(n_3450)
);

CKINVDCx20_ASAP7_75t_R g3451 ( 
.A(n_3077),
.Y(n_3451)
);

CKINVDCx5p33_ASAP7_75t_R g3452 ( 
.A(n_3069),
.Y(n_3452)
);

OAI22xp33_ASAP7_75t_L g3453 ( 
.A1(n_3201),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_3453)
);

OAI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_3056),
.A2(n_15),
.B1(n_11),
.B2(n_14),
.Y(n_3454)
);

CKINVDCx11_ASAP7_75t_R g3455 ( 
.A(n_3032),
.Y(n_3455)
);

INVx6_ASAP7_75t_L g3456 ( 
.A(n_3077),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3059),
.Y(n_3457)
);

CKINVDCx11_ASAP7_75t_R g3458 ( 
.A(n_3092),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3112),
.Y(n_3459)
);

AOI22xp33_ASAP7_75t_L g3460 ( 
.A1(n_3179),
.A2(n_1429),
.B1(n_1438),
.B2(n_1426),
.Y(n_3460)
);

AOI22xp33_ASAP7_75t_SL g3461 ( 
.A1(n_3218),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_3461)
);

AOI22xp33_ASAP7_75t_L g3462 ( 
.A1(n_3179),
.A2(n_3138),
.B1(n_3139),
.B2(n_3271),
.Y(n_3462)
);

OAI22xp5_ASAP7_75t_L g3463 ( 
.A1(n_3193),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_3463)
);

AOI22xp33_ASAP7_75t_L g3464 ( 
.A1(n_3271),
.A2(n_1438),
.B1(n_1330),
.B2(n_1350),
.Y(n_3464)
);

BUFx2_ASAP7_75t_L g3465 ( 
.A(n_3121),
.Y(n_3465)
);

INVx6_ASAP7_75t_L g3466 ( 
.A(n_3077),
.Y(n_3466)
);

OAI22xp5_ASAP7_75t_L g3467 ( 
.A1(n_3272),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3207),
.Y(n_3468)
);

BUFx2_ASAP7_75t_L g3469 ( 
.A(n_3152),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3204),
.Y(n_3470)
);

AOI22xp33_ASAP7_75t_L g3471 ( 
.A1(n_3271),
.A2(n_1438),
.B1(n_1330),
.B2(n_1350),
.Y(n_3471)
);

INVx3_ASAP7_75t_L g3472 ( 
.A(n_3122),
.Y(n_3472)
);

BUFx2_ASAP7_75t_L g3473 ( 
.A(n_3152),
.Y(n_3473)
);

BUFx12f_ASAP7_75t_L g3474 ( 
.A(n_3067),
.Y(n_3474)
);

CKINVDCx5p33_ASAP7_75t_R g3475 ( 
.A(n_3120),
.Y(n_3475)
);

BUFx2_ASAP7_75t_L g3476 ( 
.A(n_3157),
.Y(n_3476)
);

OAI22xp5_ASAP7_75t_SL g3477 ( 
.A1(n_3092),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3167),
.Y(n_3478)
);

CKINVDCx5p33_ASAP7_75t_R g3479 ( 
.A(n_3033),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3174),
.Y(n_3480)
);

AOI22xp33_ASAP7_75t_L g3481 ( 
.A1(n_3262),
.A2(n_1438),
.B1(n_1330),
.B2(n_1350),
.Y(n_3481)
);

BUFx6f_ASAP7_75t_L g3482 ( 
.A(n_3034),
.Y(n_3482)
);

AOI22xp33_ASAP7_75t_L g3483 ( 
.A1(n_3262),
.A2(n_1330),
.B1(n_1350),
.B2(n_1347),
.Y(n_3483)
);

AOI22xp33_ASAP7_75t_L g3484 ( 
.A1(n_3229),
.A2(n_1347),
.B1(n_1352),
.B2(n_1350),
.Y(n_3484)
);

AOI22xp33_ASAP7_75t_L g3485 ( 
.A1(n_3198),
.A2(n_1347),
.B1(n_1356),
.B2(n_1352),
.Y(n_3485)
);

OAI22xp5_ASAP7_75t_L g3486 ( 
.A1(n_3272),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_3486)
);

CKINVDCx5p33_ASAP7_75t_R g3487 ( 
.A(n_3033),
.Y(n_3487)
);

INVx6_ASAP7_75t_L g3488 ( 
.A(n_3067),
.Y(n_3488)
);

OAI22xp33_ASAP7_75t_L g3489 ( 
.A1(n_3201),
.A2(n_29),
.B1(n_24),
.B2(n_28),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3158),
.Y(n_3490)
);

OAI22xp33_ASAP7_75t_L g3491 ( 
.A1(n_3201),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_3491)
);

OAI22xp33_ASAP7_75t_L g3492 ( 
.A1(n_3202),
.A2(n_34),
.B1(n_30),
.B2(n_32),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3131),
.Y(n_3493)
);

OAI22xp5_ASAP7_75t_L g3494 ( 
.A1(n_3272),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_3494)
);

AOI22xp5_ASAP7_75t_L g3495 ( 
.A1(n_3009),
.A2(n_3178),
.B1(n_3252),
.B2(n_3195),
.Y(n_3495)
);

CKINVDCx6p67_ASAP7_75t_R g3496 ( 
.A(n_3240),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3226),
.Y(n_3497)
);

BUFx6f_ASAP7_75t_L g3498 ( 
.A(n_3034),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3226),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3213),
.Y(n_3500)
);

BUFx4_ASAP7_75t_SL g3501 ( 
.A(n_3023),
.Y(n_3501)
);

AOI22xp33_ASAP7_75t_SL g3502 ( 
.A1(n_3178),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_3131),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_L g3504 ( 
.A1(n_3009),
.A2(n_1347),
.B1(n_1356),
.B2(n_1352),
.Y(n_3504)
);

BUFx3_ASAP7_75t_L g3505 ( 
.A(n_3117),
.Y(n_3505)
);

CKINVDCx11_ASAP7_75t_R g3506 ( 
.A(n_3016),
.Y(n_3506)
);

BUFx12f_ASAP7_75t_L g3507 ( 
.A(n_3095),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3213),
.Y(n_3508)
);

BUFx3_ASAP7_75t_L g3509 ( 
.A(n_3117),
.Y(n_3509)
);

AOI22xp33_ASAP7_75t_L g3510 ( 
.A1(n_3212),
.A2(n_1347),
.B1(n_1356),
.B2(n_1352),
.Y(n_3510)
);

CKINVDCx11_ASAP7_75t_R g3511 ( 
.A(n_3016),
.Y(n_3511)
);

INVx6_ASAP7_75t_L g3512 ( 
.A(n_3243),
.Y(n_3512)
);

AOI22xp33_ASAP7_75t_SL g3513 ( 
.A1(n_3267),
.A2(n_3190),
.B1(n_3113),
.B2(n_3089),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3230),
.Y(n_3514)
);

INVx6_ASAP7_75t_L g3515 ( 
.A(n_3016),
.Y(n_3515)
);

BUFx8_ASAP7_75t_L g3516 ( 
.A(n_3125),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3230),
.Y(n_3517)
);

BUFx12f_ASAP7_75t_L g3518 ( 
.A(n_3202),
.Y(n_3518)
);

CKINVDCx5p33_ASAP7_75t_R g3519 ( 
.A(n_3180),
.Y(n_3519)
);

AOI22xp33_ASAP7_75t_L g3520 ( 
.A1(n_3252),
.A2(n_1352),
.B1(n_1358),
.B2(n_1356),
.Y(n_3520)
);

AND2x4_ASAP7_75t_L g3521 ( 
.A(n_3157),
.B(n_585),
.Y(n_3521)
);

CKINVDCx20_ASAP7_75t_R g3522 ( 
.A(n_3097),
.Y(n_3522)
);

OAI22xp33_ASAP7_75t_L g3523 ( 
.A1(n_3202),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_3523)
);

BUFx2_ASAP7_75t_L g3524 ( 
.A(n_3160),
.Y(n_3524)
);

BUFx2_ASAP7_75t_SL g3525 ( 
.A(n_3071),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_3348),
.B(n_3145),
.Y(n_3526)
);

AND2x4_ASAP7_75t_L g3527 ( 
.A(n_3348),
.B(n_3159),
.Y(n_3527)
);

AOI21x1_ASAP7_75t_L g3528 ( 
.A1(n_3389),
.A2(n_3200),
.B(n_3261),
.Y(n_3528)
);

AOI21x1_ASAP7_75t_L g3529 ( 
.A1(n_3428),
.A2(n_3187),
.B(n_3269),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3396),
.B(n_3145),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_3294),
.A2(n_3113),
.B(n_3264),
.Y(n_3531)
);

AND2x2_ASAP7_75t_L g3532 ( 
.A(n_3373),
.B(n_3145),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3396),
.B(n_3322),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3331),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3341),
.Y(n_3535)
);

OAI21x1_ASAP7_75t_L g3536 ( 
.A1(n_3497),
.A2(n_3147),
.B(n_3155),
.Y(n_3536)
);

AND2x4_ASAP7_75t_L g3537 ( 
.A(n_3436),
.B(n_3159),
.Y(n_3537)
);

AND2x4_ASAP7_75t_L g3538 ( 
.A(n_3376),
.B(n_3249),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_3490),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3360),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3370),
.Y(n_3541)
);

AOI21x1_ASAP7_75t_L g3542 ( 
.A1(n_3467),
.A2(n_3269),
.B(n_3127),
.Y(n_3542)
);

OA21x2_ASAP7_75t_L g3543 ( 
.A1(n_3407),
.A2(n_3184),
.B(n_3147),
.Y(n_3543)
);

AOI22xp33_ASAP7_75t_L g3544 ( 
.A1(n_3294),
.A2(n_3264),
.B1(n_3136),
.B2(n_3135),
.Y(n_3544)
);

OAI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3335),
.A2(n_3075),
.B(n_3058),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3378),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3322),
.B(n_3068),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3326),
.B(n_3251),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3380),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3326),
.B(n_3263),
.Y(n_3550)
);

INVx6_ASAP7_75t_L g3551 ( 
.A(n_3402),
.Y(n_3551)
);

AND2x4_ASAP7_75t_L g3552 ( 
.A(n_3443),
.B(n_3249),
.Y(n_3552)
);

AOI22xp33_ASAP7_75t_L g3553 ( 
.A1(n_3458),
.A2(n_3136),
.B1(n_3135),
.B2(n_3222),
.Y(n_3553)
);

BUFx6f_ASAP7_75t_L g3554 ( 
.A(n_3352),
.Y(n_3554)
);

AOI21x1_ASAP7_75t_L g3555 ( 
.A1(n_3467),
.A2(n_3127),
.B(n_3124),
.Y(n_3555)
);

OA21x2_ASAP7_75t_L g3556 ( 
.A1(n_3407),
.A2(n_3184),
.B(n_3175),
.Y(n_3556)
);

OR2x2_ASAP7_75t_L g3557 ( 
.A(n_3281),
.B(n_3289),
.Y(n_3557)
);

INVx2_ASAP7_75t_L g3558 ( 
.A(n_3280),
.Y(n_3558)
);

OA21x2_ASAP7_75t_L g3559 ( 
.A1(n_3499),
.A2(n_3001),
.B(n_3000),
.Y(n_3559)
);

OA21x2_ASAP7_75t_L g3560 ( 
.A1(n_3460),
.A2(n_3001),
.B(n_3000),
.Y(n_3560)
);

HB1xp67_ASAP7_75t_L g3561 ( 
.A(n_3325),
.Y(n_3561)
);

OAI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_3335),
.A2(n_3148),
.B(n_3028),
.Y(n_3562)
);

AO31x2_ASAP7_75t_L g3563 ( 
.A1(n_3486),
.A2(n_3177),
.A3(n_3154),
.B(n_3144),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3315),
.Y(n_3564)
);

BUFx3_ASAP7_75t_L g3565 ( 
.A(n_3390),
.Y(n_3565)
);

OAI21x1_ASAP7_75t_L g3566 ( 
.A1(n_3293),
.A2(n_3155),
.B(n_3061),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3381),
.Y(n_3567)
);

AO21x2_ASAP7_75t_L g3568 ( 
.A1(n_3292),
.A2(n_3089),
.B(n_3080),
.Y(n_3568)
);

AOI22xp33_ASAP7_75t_L g3569 ( 
.A1(n_3477),
.A2(n_3136),
.B1(n_3135),
.B2(n_3222),
.Y(n_3569)
);

A2O1A1Ixp33_ASAP7_75t_L g3570 ( 
.A1(n_3426),
.A2(n_3266),
.B(n_3084),
.C(n_3071),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3387),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3397),
.Y(n_3572)
);

NAND2xp33_ASAP7_75t_R g3573 ( 
.A(n_3316),
.B(n_3022),
.Y(n_3573)
);

AOI221xp5_ASAP7_75t_L g3574 ( 
.A1(n_3401),
.A2(n_3142),
.B1(n_3029),
.B2(n_3118),
.C(n_3188),
.Y(n_3574)
);

AOI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_3285),
.A2(n_3267),
.B(n_3242),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3406),
.Y(n_3576)
);

AND2x2_ASAP7_75t_L g3577 ( 
.A(n_3427),
.B(n_3186),
.Y(n_3577)
);

INVx3_ASAP7_75t_L g3578 ( 
.A(n_3505),
.Y(n_3578)
);

NOR2xp33_ASAP7_75t_L g3579 ( 
.A(n_3507),
.B(n_3419),
.Y(n_3579)
);

AO21x2_ASAP7_75t_L g3580 ( 
.A1(n_3486),
.A2(n_3080),
.B(n_3236),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3317),
.B(n_3182),
.Y(n_3581)
);

AOI21xp5_ASAP7_75t_SL g3582 ( 
.A1(n_3446),
.A2(n_3222),
.B(n_3243),
.Y(n_3582)
);

XOR2x2_ASAP7_75t_L g3583 ( 
.A(n_3286),
.B(n_3062),
.Y(n_3583)
);

OAI21xp5_ASAP7_75t_L g3584 ( 
.A1(n_3426),
.A2(n_3109),
.B(n_3002),
.Y(n_3584)
);

AOI222xp33_ASAP7_75t_L g3585 ( 
.A1(n_3414),
.A2(n_3246),
.B1(n_3249),
.B2(n_3177),
.C1(n_3248),
.C2(n_3243),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3459),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3468),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3465),
.B(n_3238),
.Y(n_3588)
);

AO31x2_ASAP7_75t_L g3589 ( 
.A1(n_3494),
.A2(n_3346),
.A3(n_3343),
.B(n_3338),
.Y(n_3589)
);

OAI21x1_ASAP7_75t_SL g3590 ( 
.A1(n_3345),
.A2(n_3232),
.B(n_3182),
.Y(n_3590)
);

AOI21x1_ASAP7_75t_L g3591 ( 
.A1(n_3494),
.A2(n_3363),
.B(n_3401),
.Y(n_3591)
);

OAI21x1_ASAP7_75t_L g3592 ( 
.A1(n_3293),
.A2(n_3126),
.B(n_3005),
.Y(n_3592)
);

INVxp67_ASAP7_75t_L g3593 ( 
.A(n_3420),
.Y(n_3593)
);

AOI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_3285),
.A2(n_3267),
.B(n_3242),
.Y(n_3594)
);

OAI22xp5_ASAP7_75t_L g3595 ( 
.A1(n_3284),
.A2(n_3206),
.B1(n_3116),
.B2(n_3266),
.Y(n_3595)
);

INVx4_ASAP7_75t_SL g3596 ( 
.A(n_3299),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3412),
.A2(n_3384),
.B(n_3392),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3470),
.Y(n_3598)
);

OA21x2_ASAP7_75t_L g3599 ( 
.A1(n_3462),
.A2(n_3126),
.B(n_3165),
.Y(n_3599)
);

AOI21xp33_ASAP7_75t_L g3600 ( 
.A1(n_3313),
.A2(n_3257),
.B(n_3236),
.Y(n_3600)
);

AOI21xp5_ASAP7_75t_L g3601 ( 
.A1(n_3384),
.A2(n_3044),
.B(n_3087),
.Y(n_3601)
);

OAI21xp5_ASAP7_75t_L g3602 ( 
.A1(n_3342),
.A2(n_3025),
.B(n_3050),
.Y(n_3602)
);

AND2x2_ASAP7_75t_L g3603 ( 
.A(n_3469),
.B(n_3160),
.Y(n_3603)
);

AO31x2_ASAP7_75t_L g3604 ( 
.A1(n_3343),
.A2(n_3154),
.A3(n_3144),
.B(n_3232),
.Y(n_3604)
);

OAI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_3342),
.A2(n_3103),
.B(n_3210),
.Y(n_3605)
);

AOI21xp5_ASAP7_75t_L g3606 ( 
.A1(n_3414),
.A2(n_3044),
.B(n_3087),
.Y(n_3606)
);

AND2x2_ASAP7_75t_L g3607 ( 
.A(n_3473),
.B(n_3073),
.Y(n_3607)
);

OR2x2_ASAP7_75t_L g3608 ( 
.A(n_3329),
.B(n_3064),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3323),
.Y(n_3609)
);

OAI21x1_ASAP7_75t_L g3610 ( 
.A1(n_3363),
.A2(n_3005),
.B(n_3004),
.Y(n_3610)
);

OAI21x1_ASAP7_75t_L g3611 ( 
.A1(n_3410),
.A2(n_3004),
.B(n_3140),
.Y(n_3611)
);

OR2x6_ASAP7_75t_L g3612 ( 
.A(n_3400),
.B(n_3243),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3324),
.Y(n_3613)
);

AOI22xp33_ASAP7_75t_L g3614 ( 
.A1(n_3279),
.A2(n_3073),
.B1(n_3100),
.B2(n_3079),
.Y(n_3614)
);

OR2x6_ASAP7_75t_L g3615 ( 
.A(n_3400),
.B(n_3282),
.Y(n_3615)
);

A2O1A1Ixp33_ASAP7_75t_L g3616 ( 
.A1(n_3283),
.A2(n_3248),
.B(n_3172),
.C(n_3169),
.Y(n_3616)
);

OR2x6_ASAP7_75t_L g3617 ( 
.A(n_3400),
.B(n_3248),
.Y(n_3617)
);

OAI22xp33_ASAP7_75t_L g3618 ( 
.A1(n_3495),
.A2(n_3248),
.B1(n_3079),
.B2(n_3100),
.Y(n_3618)
);

OA21x2_ASAP7_75t_L g3619 ( 
.A1(n_3311),
.A2(n_3165),
.B(n_3024),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_3336),
.Y(n_3620)
);

INVx2_ASAP7_75t_L g3621 ( 
.A(n_3366),
.Y(n_3621)
);

AOI22xp33_ASAP7_75t_L g3622 ( 
.A1(n_3279),
.A2(n_3190),
.B1(n_3133),
.B2(n_3022),
.Y(n_3622)
);

AOI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_3385),
.A2(n_3044),
.B(n_3087),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3367),
.B(n_3064),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3374),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3398),
.B(n_3210),
.Y(n_3626)
);

OR2x2_ASAP7_75t_L g3627 ( 
.A(n_3295),
.B(n_3103),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3431),
.B(n_3180),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_3437),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3442),
.B(n_3450),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3297),
.Y(n_3631)
);

OA21x2_ASAP7_75t_L g3632 ( 
.A1(n_3321),
.A2(n_3024),
.B(n_3018),
.Y(n_3632)
);

AND2x4_ASAP7_75t_L g3633 ( 
.A(n_3476),
.B(n_3130),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3298),
.B(n_3130),
.Y(n_3634)
);

INVx2_ASAP7_75t_SL g3635 ( 
.A(n_3395),
.Y(n_3635)
);

OAI211xp5_ASAP7_75t_L g3636 ( 
.A1(n_3408),
.A2(n_3253),
.B(n_3127),
.C(n_3275),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3300),
.B(n_3130),
.Y(n_3637)
);

AO31x2_ASAP7_75t_L g3638 ( 
.A1(n_3346),
.A2(n_3173),
.A3(n_3205),
.B(n_3216),
.Y(n_3638)
);

OAI22xp5_ASAP7_75t_L g3639 ( 
.A1(n_3296),
.A2(n_3241),
.B1(n_3214),
.B2(n_3169),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_SL g3640 ( 
.A(n_3382),
.B(n_3016),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_3524),
.B(n_3383),
.Y(n_3641)
);

BUFx6f_ASAP7_75t_L g3642 ( 
.A(n_3352),
.Y(n_3642)
);

OAI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_3364),
.A2(n_3164),
.B(n_3146),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3301),
.Y(n_3644)
);

AOI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_3385),
.A2(n_3133),
.B(n_3216),
.Y(n_3645)
);

OA21x2_ASAP7_75t_L g3646 ( 
.A1(n_3302),
.A2(n_3035),
.B(n_3018),
.Y(n_3646)
);

OAI21x1_ASAP7_75t_L g3647 ( 
.A1(n_3410),
.A2(n_3140),
.B(n_3046),
.Y(n_3647)
);

AOI22xp33_ASAP7_75t_L g3648 ( 
.A1(n_3408),
.A2(n_3253),
.B1(n_3275),
.B2(n_3172),
.Y(n_3648)
);

INVx4_ASAP7_75t_L g3649 ( 
.A(n_3352),
.Y(n_3649)
);

OAI222xp33_ASAP7_75t_L g3650 ( 
.A1(n_3463),
.A2(n_3353),
.B1(n_3502),
.B2(n_3375),
.C1(n_3359),
.C2(n_3379),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3441),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3447),
.Y(n_3652)
);

AO31x2_ASAP7_75t_L g3653 ( 
.A1(n_3338),
.A2(n_3173),
.A3(n_3205),
.B(n_3231),
.Y(n_3653)
);

HB1xp67_ASAP7_75t_L g3654 ( 
.A(n_3344),
.Y(n_3654)
);

AO21x2_ASAP7_75t_L g3655 ( 
.A1(n_3457),
.A2(n_3356),
.B(n_3354),
.Y(n_3655)
);

OAI22xp5_ASAP7_75t_L g3656 ( 
.A1(n_3359),
.A2(n_3241),
.B1(n_3214),
.B2(n_3164),
.Y(n_3656)
);

INVx4_ASAP7_75t_SL g3657 ( 
.A(n_3299),
.Y(n_3657)
);

BUFx8_ASAP7_75t_L g3658 ( 
.A(n_3291),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3500),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3508),
.Y(n_3660)
);

OA21x2_ASAP7_75t_L g3661 ( 
.A1(n_3357),
.A2(n_3046),
.B(n_3035),
.Y(n_3661)
);

NOR2xp33_ASAP7_75t_L g3662 ( 
.A(n_3452),
.B(n_3023),
.Y(n_3662)
);

OAI22xp33_ASAP7_75t_L g3663 ( 
.A1(n_3463),
.A2(n_3030),
.B1(n_3168),
.B2(n_3130),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3514),
.Y(n_3664)
);

AOI22xp33_ASAP7_75t_L g3665 ( 
.A1(n_3364),
.A2(n_3231),
.B1(n_3181),
.B2(n_3168),
.Y(n_3665)
);

NAND2xp33_ASAP7_75t_R g3666 ( 
.A(n_3361),
.B(n_3146),
.Y(n_3666)
);

AOI22xp5_ASAP7_75t_L g3667 ( 
.A1(n_3446),
.A2(n_3141),
.B1(n_3030),
.B2(n_3265),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3478),
.B(n_3168),
.Y(n_3668)
);

OR2x6_ASAP7_75t_L g3669 ( 
.A(n_3282),
.B(n_3168),
.Y(n_3669)
);

OR2x2_ASAP7_75t_L g3670 ( 
.A(n_3413),
.B(n_3181),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3480),
.Y(n_3671)
);

AND2x4_ASAP7_75t_L g3672 ( 
.A(n_3418),
.B(n_3181),
.Y(n_3672)
);

AOI22xp33_ASAP7_75t_SL g3673 ( 
.A1(n_3518),
.A2(n_3181),
.B1(n_3237),
.B2(n_3235),
.Y(n_3673)
);

INVx2_ASAP7_75t_SL g3674 ( 
.A(n_3501),
.Y(n_3674)
);

AND2x2_ASAP7_75t_L g3675 ( 
.A(n_3403),
.B(n_3235),
.Y(n_3675)
);

OR2x2_ASAP7_75t_L g3676 ( 
.A(n_3421),
.B(n_3235),
.Y(n_3676)
);

AOI22xp33_ASAP7_75t_L g3677 ( 
.A1(n_3461),
.A2(n_3237),
.B1(n_3239),
.B2(n_3235),
.Y(n_3677)
);

AND2x4_ASAP7_75t_L g3678 ( 
.A(n_3430),
.B(n_3237),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3433),
.Y(n_3679)
);

OA21x2_ASAP7_75t_L g3680 ( 
.A1(n_3434),
.A2(n_3197),
.B(n_3268),
.Y(n_3680)
);

BUFx6f_ASAP7_75t_L g3681 ( 
.A(n_3308),
.Y(n_3681)
);

BUFx2_ASAP7_75t_L g3682 ( 
.A(n_3509),
.Y(n_3682)
);

AOI22xp33_ASAP7_75t_L g3683 ( 
.A1(n_3461),
.A2(n_3239),
.B1(n_3237),
.B2(n_3101),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3328),
.B(n_3239),
.Y(n_3684)
);

AOI22xp33_ASAP7_75t_L g3685 ( 
.A1(n_3502),
.A2(n_3239),
.B1(n_3101),
.B2(n_3105),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3493),
.B(n_3081),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3503),
.Y(n_3687)
);

AND2x2_ASAP7_75t_L g3688 ( 
.A(n_3351),
.B(n_3081),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3517),
.Y(n_3689)
);

AND2x2_ASAP7_75t_L g3690 ( 
.A(n_3445),
.B(n_3081),
.Y(n_3690)
);

A2O1A1Ixp33_ASAP7_75t_L g3691 ( 
.A1(n_3305),
.A2(n_3265),
.B(n_3101),
.C(n_3105),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3375),
.B(n_3081),
.Y(n_3692)
);

OA21x2_ASAP7_75t_L g3693 ( 
.A1(n_3368),
.A2(n_3197),
.B(n_3268),
.Y(n_3693)
);

OA21x2_ASAP7_75t_L g3694 ( 
.A1(n_3388),
.A2(n_3211),
.B(n_3209),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3513),
.Y(n_3695)
);

OAI21x1_ASAP7_75t_L g3696 ( 
.A1(n_3307),
.A2(n_3111),
.B(n_3209),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3327),
.B(n_3101),
.Y(n_3697)
);

AND2x4_ASAP7_75t_L g3698 ( 
.A(n_3307),
.B(n_3105),
.Y(n_3698)
);

CKINVDCx11_ASAP7_75t_R g3699 ( 
.A(n_3278),
.Y(n_3699)
);

OAI21xp5_ASAP7_75t_L g3700 ( 
.A1(n_3333),
.A2(n_3047),
.B(n_3006),
.Y(n_3700)
);

AOI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_3340),
.A2(n_3141),
.B(n_3047),
.Y(n_3701)
);

OAI21xp5_ASAP7_75t_L g3702 ( 
.A1(n_3304),
.A2(n_3006),
.B(n_3255),
.Y(n_3702)
);

OAI22xp33_ASAP7_75t_L g3703 ( 
.A1(n_3496),
.A2(n_3105),
.B1(n_3041),
.B2(n_3049),
.Y(n_3703)
);

O2A1O1Ixp5_ASAP7_75t_L g3704 ( 
.A1(n_3439),
.A2(n_3041),
.B(n_3049),
.C(n_3036),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3365),
.Y(n_3705)
);

OAI21xp5_ASAP7_75t_L g3706 ( 
.A1(n_3379),
.A2(n_3220),
.B(n_3211),
.Y(n_3706)
);

AOI21xp5_ASAP7_75t_L g3707 ( 
.A1(n_3340),
.A2(n_3221),
.B(n_3220),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_3327),
.A2(n_3250),
.B(n_3221),
.Y(n_3708)
);

OR2x2_ASAP7_75t_L g3709 ( 
.A(n_3365),
.B(n_3036),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3449),
.B(n_3036),
.Y(n_3710)
);

AOI21xp5_ASAP7_75t_L g3711 ( 
.A1(n_3464),
.A2(n_3250),
.B(n_3041),
.Y(n_3711)
);

AND2x2_ASAP7_75t_L g3712 ( 
.A(n_3339),
.B(n_3036),
.Y(n_3712)
);

AOI21xp5_ASAP7_75t_L g3713 ( 
.A1(n_3471),
.A2(n_3049),
.B(n_3041),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3513),
.Y(n_3714)
);

OAI21x1_ASAP7_75t_L g3715 ( 
.A1(n_3449),
.A2(n_3049),
.B(n_587),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3472),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3472),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3282),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3320),
.B(n_39),
.Y(n_3719)
);

AND2x4_ASAP7_75t_L g3720 ( 
.A(n_3404),
.B(n_39),
.Y(n_3720)
);

AOI22xp33_ASAP7_75t_SL g3721 ( 
.A1(n_3516),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_3721)
);

INVx3_ASAP7_75t_L g3722 ( 
.A(n_3309),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3522),
.B(n_40),
.Y(n_3723)
);

AND2x2_ASAP7_75t_L g3724 ( 
.A(n_3479),
.B(n_41),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3309),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3309),
.Y(n_3726)
);

BUFx2_ASAP7_75t_L g3727 ( 
.A(n_3519),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3404),
.Y(n_3728)
);

AOI21xp5_ASAP7_75t_L g3729 ( 
.A1(n_3504),
.A2(n_1358),
.B(n_1356),
.Y(n_3729)
);

AOI21x1_ASAP7_75t_L g3730 ( 
.A1(n_3454),
.A2(n_42),
.B(n_43),
.Y(n_3730)
);

OAI22xp5_ASAP7_75t_L g3731 ( 
.A1(n_3306),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_SL g3732 ( 
.A(n_3422),
.B(n_1358),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3312),
.B(n_44),
.Y(n_3733)
);

AOI221xp5_ASAP7_75t_L g3734 ( 
.A1(n_3453),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.C(n_48),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3404),
.Y(n_3735)
);

BUFx6f_ASAP7_75t_L g3736 ( 
.A(n_3681),
.Y(n_3736)
);

INVx2_ASAP7_75t_L g3737 ( 
.A(n_3716),
.Y(n_3737)
);

INVx4_ASAP7_75t_SL g3738 ( 
.A(n_3681),
.Y(n_3738)
);

OAI21x1_ASAP7_75t_L g3739 ( 
.A1(n_3575),
.A2(n_3391),
.B(n_3424),
.Y(n_3739)
);

AOI21xp33_ASAP7_75t_L g3740 ( 
.A1(n_3719),
.A2(n_3562),
.B(n_3733),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_SL g3741 ( 
.A(n_3681),
.B(n_3371),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_3641),
.B(n_3415),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3716),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3534),
.Y(n_3744)
);

OAI221xp5_ASAP7_75t_L g3745 ( 
.A1(n_3721),
.A2(n_3337),
.B1(n_3319),
.B2(n_3314),
.C(n_3347),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_3531),
.A2(n_3523),
.B(n_3491),
.Y(n_3746)
);

A2O1A1Ixp33_ASAP7_75t_L g3747 ( 
.A1(n_3545),
.A2(n_3454),
.B(n_3438),
.C(n_3369),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3534),
.Y(n_3748)
);

OAI21x1_ASAP7_75t_L g3749 ( 
.A1(n_3594),
.A2(n_3394),
.B(n_3393),
.Y(n_3749)
);

OAI22xp5_ASAP7_75t_L g3750 ( 
.A1(n_3570),
.A2(n_3492),
.B1(n_3489),
.B2(n_3358),
.Y(n_3750)
);

OAI211xp5_ASAP7_75t_L g3751 ( 
.A1(n_3734),
.A2(n_3290),
.B(n_3416),
.C(n_3429),
.Y(n_3751)
);

AOI22xp33_ASAP7_75t_L g3752 ( 
.A1(n_3584),
.A2(n_3516),
.B1(n_3318),
.B2(n_3405),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3717),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3535),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3535),
.Y(n_3755)
);

AOI22xp33_ASAP7_75t_L g3756 ( 
.A1(n_3544),
.A2(n_3318),
.B1(n_3456),
.B2(n_3358),
.Y(n_3756)
);

AOI31xp33_ASAP7_75t_L g3757 ( 
.A1(n_3640),
.A2(n_3475),
.A3(n_3411),
.B(n_3487),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3588),
.B(n_3372),
.Y(n_3758)
);

AOI221xp5_ASAP7_75t_L g3759 ( 
.A1(n_3650),
.A2(n_3423),
.B1(n_3422),
.B2(n_3444),
.C(n_3425),
.Y(n_3759)
);

OAI22xp5_ASAP7_75t_L g3760 ( 
.A1(n_3569),
.A2(n_3466),
.B1(n_3456),
.B2(n_3451),
.Y(n_3760)
);

AOI21xp5_ASAP7_75t_L g3761 ( 
.A1(n_3645),
.A2(n_3521),
.B(n_3303),
.Y(n_3761)
);

AOI22xp33_ASAP7_75t_L g3762 ( 
.A1(n_3731),
.A2(n_3466),
.B1(n_3362),
.B2(n_3399),
.Y(n_3762)
);

OAI211xp5_ASAP7_75t_SL g3763 ( 
.A1(n_3602),
.A2(n_3386),
.B(n_3349),
.C(n_3409),
.Y(n_3763)
);

OAI22xp5_ASAP7_75t_SL g3764 ( 
.A1(n_3635),
.A2(n_3330),
.B1(n_3377),
.B2(n_3334),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3577),
.B(n_3402),
.Y(n_3765)
);

AOI22xp33_ASAP7_75t_L g3766 ( 
.A1(n_3639),
.A2(n_3350),
.B1(n_3521),
.B2(n_3474),
.Y(n_3766)
);

AOI22xp33_ASAP7_75t_L g3767 ( 
.A1(n_3585),
.A2(n_3350),
.B1(n_3355),
.B2(n_3435),
.Y(n_3767)
);

OAI33xp33_ASAP7_75t_L g3768 ( 
.A1(n_3695),
.A2(n_50),
.A3(n_52),
.B1(n_46),
.B2(n_48),
.B3(n_51),
.Y(n_3768)
);

AOI22xp5_ASAP7_75t_L g3769 ( 
.A1(n_3663),
.A2(n_3355),
.B1(n_3310),
.B2(n_3332),
.Y(n_3769)
);

OAI22xp5_ASAP7_75t_L g3770 ( 
.A1(n_3648),
.A2(n_3310),
.B1(n_3332),
.B2(n_3303),
.Y(n_3770)
);

AOI22xp33_ASAP7_75t_L g3771 ( 
.A1(n_3618),
.A2(n_3595),
.B1(n_3614),
.B2(n_3684),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3717),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3705),
.Y(n_3773)
);

HB1xp67_ASAP7_75t_L g3774 ( 
.A(n_3532),
.Y(n_3774)
);

OAI22xp5_ASAP7_75t_L g3775 ( 
.A1(n_3665),
.A2(n_3310),
.B1(n_3303),
.B2(n_3287),
.Y(n_3775)
);

AND2x4_ASAP7_75t_L g3776 ( 
.A(n_3718),
.B(n_3448),
.Y(n_3776)
);

AOI22xp5_ASAP7_75t_L g3777 ( 
.A1(n_3656),
.A2(n_3488),
.B1(n_3512),
.B2(n_3515),
.Y(n_3777)
);

NOR2xp33_ASAP7_75t_L g3778 ( 
.A(n_3551),
.B(n_3455),
.Y(n_3778)
);

AOI22xp33_ASAP7_75t_SL g3779 ( 
.A1(n_3636),
.A2(n_3287),
.B1(n_3512),
.B2(n_3488),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3654),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3526),
.B(n_3448),
.Y(n_3781)
);

OAI21x1_ASAP7_75t_L g3782 ( 
.A1(n_3529),
.A2(n_3417),
.B(n_3481),
.Y(n_3782)
);

OAI211xp5_ASAP7_75t_SL g3783 ( 
.A1(n_3574),
.A2(n_3506),
.B(n_3511),
.C(n_3484),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3557),
.Y(n_3784)
);

AOI221xp5_ASAP7_75t_L g3785 ( 
.A1(n_3695),
.A2(n_3520),
.B1(n_3525),
.B2(n_3498),
.C(n_3482),
.Y(n_3785)
);

OAI221xp5_ASAP7_75t_L g3786 ( 
.A1(n_3685),
.A2(n_3512),
.B1(n_3287),
.B2(n_3432),
.C(n_3440),
.Y(n_3786)
);

AOI22xp33_ASAP7_75t_L g3787 ( 
.A1(n_3590),
.A2(n_3600),
.B1(n_3714),
.B2(n_3697),
.Y(n_3787)
);

BUFx3_ASAP7_75t_L g3788 ( 
.A(n_3565),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3655),
.Y(n_3789)
);

A2O1A1Ixp33_ASAP7_75t_L g3790 ( 
.A1(n_3704),
.A2(n_3510),
.B(n_3485),
.C(n_3448),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3631),
.Y(n_3791)
);

AOI21x1_ASAP7_75t_L g3792 ( 
.A1(n_3528),
.A2(n_3288),
.B(n_3515),
.Y(n_3792)
);

AOI222xp33_ASAP7_75t_L g3793 ( 
.A1(n_3622),
.A2(n_52),
.B1(n_54),
.B2(n_50),
.C1(n_51),
.C2(n_53),
.Y(n_3793)
);

AOI21xp5_ASAP7_75t_L g3794 ( 
.A1(n_3582),
.A2(n_3483),
.B(n_3482),
.Y(n_3794)
);

AND2x2_ASAP7_75t_L g3795 ( 
.A(n_3682),
.B(n_3498),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3631),
.Y(n_3796)
);

AOI22xp33_ASAP7_75t_L g3797 ( 
.A1(n_3714),
.A2(n_3498),
.B1(n_3482),
.B2(n_1358),
.Y(n_3797)
);

OAI221xp5_ASAP7_75t_L g3798 ( 
.A1(n_3591),
.A2(n_56),
.B1(n_53),
.B2(n_54),
.C(n_57),
.Y(n_3798)
);

AOI22xp33_ASAP7_75t_SL g3799 ( 
.A1(n_3597),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_3799)
);

NOR2x1p5_ASAP7_75t_L g3800 ( 
.A(n_3722),
.B(n_58),
.Y(n_3800)
);

OAI22xp33_ASAP7_75t_L g3801 ( 
.A1(n_3667),
.A2(n_62),
.B1(n_59),
.B2(n_60),
.Y(n_3801)
);

BUFx3_ASAP7_75t_L g3802 ( 
.A(n_3658),
.Y(n_3802)
);

OR2x2_ASAP7_75t_L g3803 ( 
.A(n_3530),
.B(n_3533),
.Y(n_3803)
);

AND2x2_ASAP7_75t_L g3804 ( 
.A(n_3603),
.B(n_63),
.Y(n_3804)
);

AOI22xp33_ASAP7_75t_L g3805 ( 
.A1(n_3553),
.A2(n_1358),
.B1(n_1372),
.B2(n_1430),
.Y(n_3805)
);

AOI22xp33_ASAP7_75t_L g3806 ( 
.A1(n_3702),
.A2(n_3605),
.B1(n_3683),
.B2(n_3677),
.Y(n_3806)
);

OAI221xp5_ASAP7_75t_L g3807 ( 
.A1(n_3616),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.C(n_67),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3540),
.Y(n_3808)
);

OR2x2_ASAP7_75t_L g3809 ( 
.A(n_3561),
.B(n_64),
.Y(n_3809)
);

AOI22xp33_ASAP7_75t_L g3810 ( 
.A1(n_3723),
.A2(n_1372),
.B1(n_1430),
.B2(n_1283),
.Y(n_3810)
);

OAI22xp5_ASAP7_75t_L g3811 ( 
.A1(n_3730),
.A2(n_68),
.B1(n_65),
.B2(n_67),
.Y(n_3811)
);

AOI22xp33_ASAP7_75t_L g3812 ( 
.A1(n_3551),
.A2(n_3700),
.B1(n_3720),
.B2(n_3692),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3609),
.B(n_70),
.Y(n_3813)
);

OAI21x1_ASAP7_75t_L g3814 ( 
.A1(n_3623),
.A2(n_3555),
.B(n_3601),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3541),
.Y(n_3815)
);

O2A1O1Ixp33_ASAP7_75t_SL g3816 ( 
.A1(n_3674),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_3816)
);

OAI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3701),
.A2(n_71),
.B(n_73),
.Y(n_3817)
);

OAI22xp5_ASAP7_75t_SL g3818 ( 
.A1(n_3579),
.A2(n_76),
.B1(n_73),
.B2(n_75),
.Y(n_3818)
);

AOI22xp33_ASAP7_75t_L g3819 ( 
.A1(n_3720),
.A2(n_1372),
.B1(n_1430),
.B2(n_1283),
.Y(n_3819)
);

HB1xp67_ASAP7_75t_L g3820 ( 
.A(n_3527),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3546),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3549),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3567),
.Y(n_3823)
);

OR2x2_ASAP7_75t_L g3824 ( 
.A(n_3608),
.B(n_77),
.Y(n_3824)
);

CKINVDCx5p33_ASAP7_75t_R g3825 ( 
.A(n_3699),
.Y(n_3825)
);

OAI211xp5_ASAP7_75t_L g3826 ( 
.A1(n_3691),
.A2(n_80),
.B(n_78),
.C(n_79),
.Y(n_3826)
);

OAI22xp5_ASAP7_75t_L g3827 ( 
.A1(n_3606),
.A2(n_81),
.B1(n_78),
.B2(n_79),
.Y(n_3827)
);

OAI22xp5_ASAP7_75t_L g3828 ( 
.A1(n_3593),
.A2(n_84),
.B1(n_81),
.B2(n_82),
.Y(n_3828)
);

BUFx12f_ASAP7_75t_L g3829 ( 
.A(n_3658),
.Y(n_3829)
);

AOI22xp33_ASAP7_75t_SL g3830 ( 
.A1(n_3643),
.A2(n_86),
.B1(n_82),
.B2(n_84),
.Y(n_3830)
);

BUFx3_ASAP7_75t_L g3831 ( 
.A(n_3727),
.Y(n_3831)
);

OAI21x1_ASAP7_75t_L g3832 ( 
.A1(n_3542),
.A2(n_86),
.B(n_87),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3571),
.Y(n_3833)
);

BUFx6f_ASAP7_75t_L g3834 ( 
.A(n_3554),
.Y(n_3834)
);

AO21x1_ASAP7_75t_SL g3835 ( 
.A1(n_3718),
.A2(n_3726),
.B(n_3725),
.Y(n_3835)
);

OAI222xp33_ASAP7_75t_L g3836 ( 
.A1(n_3673),
.A2(n_90),
.B1(n_92),
.B2(n_88),
.C1(n_89),
.C2(n_91),
.Y(n_3836)
);

OAI21xp33_ASAP7_75t_L g3837 ( 
.A1(n_3628),
.A2(n_89),
.B(n_91),
.Y(n_3837)
);

OAI22xp5_ASAP7_75t_L g3838 ( 
.A1(n_3547),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_3838)
);

NOR2xp33_ASAP7_75t_L g3839 ( 
.A(n_3662),
.B(n_93),
.Y(n_3839)
);

CKINVDCx20_ASAP7_75t_R g3840 ( 
.A(n_3596),
.Y(n_3840)
);

OAI211xp5_ASAP7_75t_SL g3841 ( 
.A1(n_3548),
.A2(n_98),
.B(n_94),
.C(n_95),
.Y(n_3841)
);

AOI22xp33_ASAP7_75t_L g3842 ( 
.A1(n_3568),
.A2(n_3537),
.B1(n_3607),
.B2(n_3724),
.Y(n_3842)
);

INVx4_ASAP7_75t_L g3843 ( 
.A(n_3596),
.Y(n_3843)
);

OAI22xp33_ASAP7_75t_L g3844 ( 
.A1(n_3615),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_3844)
);

OA21x2_ASAP7_75t_L g3845 ( 
.A1(n_3725),
.A2(n_99),
.B(n_100),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3572),
.Y(n_3846)
);

AOI22xp33_ASAP7_75t_L g3847 ( 
.A1(n_3537),
.A2(n_1372),
.B1(n_1430),
.B2(n_1283),
.Y(n_3847)
);

OAI221xp5_ASAP7_75t_L g3848 ( 
.A1(n_3706),
.A2(n_104),
.B1(n_101),
.B2(n_102),
.C(n_106),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3576),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_3613),
.B(n_102),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_3625),
.B(n_104),
.Y(n_3851)
);

OAI21xp33_ASAP7_75t_L g3852 ( 
.A1(n_3550),
.A2(n_107),
.B(n_108),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3578),
.B(n_3527),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3586),
.Y(n_3854)
);

AOI21xp33_ASAP7_75t_L g3855 ( 
.A1(n_3556),
.A2(n_110),
.B(n_111),
.Y(n_3855)
);

AOI22xp33_ASAP7_75t_L g3856 ( 
.A1(n_3726),
.A2(n_1372),
.B1(n_1430),
.B2(n_1283),
.Y(n_3856)
);

INVx2_ASAP7_75t_SL g3857 ( 
.A(n_3578),
.Y(n_3857)
);

AOI22xp33_ASAP7_75t_L g3858 ( 
.A1(n_3690),
.A2(n_1430),
.B1(n_115),
.B2(n_112),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3587),
.Y(n_3859)
);

AND2x2_ASAP7_75t_L g3860 ( 
.A(n_3712),
.B(n_112),
.Y(n_3860)
);

BUFx4f_ASAP7_75t_SL g3861 ( 
.A(n_3554),
.Y(n_3861)
);

AOI22xp33_ASAP7_75t_L g3862 ( 
.A1(n_3694),
.A2(n_116),
.B1(n_113),
.B2(n_115),
.Y(n_3862)
);

OAI221xp5_ASAP7_75t_L g3863 ( 
.A1(n_3573),
.A2(n_118),
.B1(n_113),
.B2(n_117),
.C(n_120),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3598),
.Y(n_3864)
);

AOI221xp5_ASAP7_75t_L g3865 ( 
.A1(n_3644),
.A2(n_125),
.B1(n_122),
.B2(n_123),
.C(n_126),
.Y(n_3865)
);

OAI22xp5_ASAP7_75t_L g3866 ( 
.A1(n_3627),
.A2(n_3713),
.B1(n_3626),
.B2(n_3637),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3651),
.Y(n_3867)
);

AOI22xp33_ASAP7_75t_L g3868 ( 
.A1(n_3694),
.A2(n_130),
.B1(n_127),
.B2(n_128),
.Y(n_3868)
);

AOI22xp33_ASAP7_75t_SL g3869 ( 
.A1(n_3538),
.A2(n_133),
.B1(n_127),
.B2(n_131),
.Y(n_3869)
);

OAI21x1_ASAP7_75t_L g3870 ( 
.A1(n_3707),
.A2(n_131),
.B(n_134),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3687),
.Y(n_3871)
);

HB1xp67_ASAP7_75t_L g3872 ( 
.A(n_3670),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3687),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3652),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3659),
.Y(n_3875)
);

HB1xp67_ASAP7_75t_L g3876 ( 
.A(n_3676),
.Y(n_3876)
);

OAI21x1_ASAP7_75t_L g3877 ( 
.A1(n_3536),
.A2(n_135),
.B(n_136),
.Y(n_3877)
);

OA21x2_ASAP7_75t_L g3878 ( 
.A1(n_3689),
.A2(n_135),
.B(n_136),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3689),
.B(n_137),
.Y(n_3879)
);

AOI222xp33_ASAP7_75t_L g3880 ( 
.A1(n_3657),
.A2(n_140),
.B1(n_142),
.B2(n_138),
.C1(n_139),
.C2(n_141),
.Y(n_3880)
);

INVx2_ASAP7_75t_L g3881 ( 
.A(n_3539),
.Y(n_3881)
);

AOI221xp5_ASAP7_75t_L g3882 ( 
.A1(n_3630),
.A2(n_141),
.B1(n_138),
.B2(n_140),
.C(n_142),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3660),
.Y(n_3883)
);

AOI221xp5_ASAP7_75t_L g3884 ( 
.A1(n_3664),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.C(n_148),
.Y(n_3884)
);

AOI22xp33_ASAP7_75t_L g3885 ( 
.A1(n_3732),
.A2(n_150),
.B1(n_144),
.B2(n_145),
.Y(n_3885)
);

OA21x2_ASAP7_75t_L g3886 ( 
.A1(n_3679),
.A2(n_150),
.B(n_151),
.Y(n_3886)
);

HB1xp67_ASAP7_75t_L g3887 ( 
.A(n_3604),
.Y(n_3887)
);

INVx3_ASAP7_75t_L g3888 ( 
.A(n_3722),
.Y(n_3888)
);

AOI221xp5_ASAP7_75t_L g3889 ( 
.A1(n_3703),
.A2(n_156),
.B1(n_152),
.B2(n_154),
.C(n_158),
.Y(n_3889)
);

AOI22xp33_ASAP7_75t_L g3890 ( 
.A1(n_3538),
.A2(n_159),
.B1(n_154),
.B2(n_158),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3558),
.B(n_159),
.Y(n_3891)
);

AOI221xp5_ASAP7_75t_L g3892 ( 
.A1(n_3634),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.C(n_165),
.Y(n_3892)
);

NOR2xp33_ASAP7_75t_L g3893 ( 
.A(n_3657),
.B(n_161),
.Y(n_3893)
);

BUFx6f_ASAP7_75t_L g3894 ( 
.A(n_3554),
.Y(n_3894)
);

AOI22xp33_ASAP7_75t_L g3895 ( 
.A1(n_3688),
.A2(n_167),
.B1(n_162),
.B2(n_166),
.Y(n_3895)
);

O2A1O1Ixp33_ASAP7_75t_L g3896 ( 
.A1(n_3708),
.A2(n_170),
.B(n_168),
.C(n_169),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3564),
.Y(n_3897)
);

OAI21xp5_ASAP7_75t_SL g3898 ( 
.A1(n_3552),
.A2(n_169),
.B(n_170),
.Y(n_3898)
);

AND2x2_ASAP7_75t_L g3899 ( 
.A(n_3675),
.B(n_171),
.Y(n_3899)
);

NOR2xp33_ASAP7_75t_L g3900 ( 
.A(n_3649),
.B(n_171),
.Y(n_3900)
);

AOI222xp33_ASAP7_75t_L g3901 ( 
.A1(n_3583),
.A2(n_176),
.B1(n_178),
.B2(n_173),
.C1(n_174),
.C2(n_177),
.Y(n_3901)
);

AOI22xp5_ASAP7_75t_L g3902 ( 
.A1(n_3666),
.A2(n_177),
.B1(n_173),
.B2(n_176),
.Y(n_3902)
);

AOI22xp33_ASAP7_75t_L g3903 ( 
.A1(n_3693),
.A2(n_181),
.B1(n_178),
.B2(n_180),
.Y(n_3903)
);

OAI211xp5_ASAP7_75t_L g3904 ( 
.A1(n_3668),
.A2(n_185),
.B(n_182),
.C(n_183),
.Y(n_3904)
);

HB1xp67_ASAP7_75t_L g3905 ( 
.A(n_3604),
.Y(n_3905)
);

OAI22xp5_ASAP7_75t_L g3906 ( 
.A1(n_3552),
.A2(n_186),
.B1(n_183),
.B2(n_185),
.Y(n_3906)
);

AND2x2_ASAP7_75t_L g3907 ( 
.A(n_3835),
.B(n_3633),
.Y(n_3907)
);

OR2x2_ASAP7_75t_L g3908 ( 
.A(n_3803),
.B(n_3563),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3744),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3748),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3866),
.B(n_3620),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3754),
.Y(n_3912)
);

AND2x2_ASAP7_75t_L g3913 ( 
.A(n_3774),
.B(n_3633),
.Y(n_3913)
);

AND2x4_ASAP7_75t_SL g3914 ( 
.A(n_3843),
.B(n_3615),
.Y(n_3914)
);

OAI21x1_ASAP7_75t_SL g3915 ( 
.A1(n_3843),
.A2(n_3629),
.B(n_3621),
.Y(n_3915)
);

HB1xp67_ASAP7_75t_L g3916 ( 
.A(n_3872),
.Y(n_3916)
);

OR2x2_ASAP7_75t_L g3917 ( 
.A(n_3781),
.B(n_3563),
.Y(n_3917)
);

NOR2x1_ASAP7_75t_SL g3918 ( 
.A(n_3866),
.B(n_3792),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3887),
.Y(n_3919)
);

BUFx2_ASAP7_75t_L g3920 ( 
.A(n_3845),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3755),
.Y(n_3921)
);

OR2x2_ASAP7_75t_L g3922 ( 
.A(n_3781),
.B(n_3563),
.Y(n_3922)
);

INVx2_ASAP7_75t_SL g3923 ( 
.A(n_3820),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3905),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3853),
.B(n_3589),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3789),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_3787),
.B(n_3671),
.Y(n_3927)
);

BUFx3_ASAP7_75t_L g3928 ( 
.A(n_3829),
.Y(n_3928)
);

INVx1_ASAP7_75t_SL g3929 ( 
.A(n_3825),
.Y(n_3929)
);

INVx3_ASAP7_75t_L g3930 ( 
.A(n_3888),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3888),
.B(n_3589),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3780),
.B(n_3735),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3791),
.Y(n_3933)
);

AND2x2_ASAP7_75t_L g3934 ( 
.A(n_3876),
.B(n_3589),
.Y(n_3934)
);

AND2x2_ASAP7_75t_L g3935 ( 
.A(n_3795),
.B(n_3728),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3796),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3875),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3883),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3737),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_3743),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3808),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3815),
.Y(n_3942)
);

HB1xp67_ASAP7_75t_L g3943 ( 
.A(n_3753),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3821),
.Y(n_3944)
);

BUFx6f_ASAP7_75t_L g3945 ( 
.A(n_3736),
.Y(n_3945)
);

INVx2_ASAP7_75t_L g3946 ( 
.A(n_3772),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3822),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3871),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3823),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3833),
.Y(n_3950)
);

HB1xp67_ASAP7_75t_L g3951 ( 
.A(n_3881),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3873),
.Y(n_3952)
);

AND2x2_ASAP7_75t_L g3953 ( 
.A(n_3857),
.B(n_3672),
.Y(n_3953)
);

AND2x4_ASAP7_75t_SL g3954 ( 
.A(n_3840),
.B(n_3612),
.Y(n_3954)
);

AO21x2_ASAP7_75t_L g3955 ( 
.A1(n_3855),
.A2(n_3696),
.B(n_3710),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3784),
.B(n_3672),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_3842),
.B(n_3776),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3776),
.B(n_3758),
.Y(n_3958)
);

AOI221xp5_ASAP7_75t_L g3959 ( 
.A1(n_3740),
.A2(n_3624),
.B1(n_3581),
.B2(n_3686),
.C(n_3678),
.Y(n_3959)
);

OR2x2_ASAP7_75t_L g3960 ( 
.A(n_3897),
.B(n_3556),
.Y(n_3960)
);

BUFx3_ASAP7_75t_L g3961 ( 
.A(n_3802),
.Y(n_3961)
);

INVx3_ASAP7_75t_L g3962 ( 
.A(n_3845),
.Y(n_3962)
);

HB1xp67_ASAP7_75t_L g3963 ( 
.A(n_3846),
.Y(n_3963)
);

INVx2_ASAP7_75t_L g3964 ( 
.A(n_3878),
.Y(n_3964)
);

INVx2_ASAP7_75t_L g3965 ( 
.A(n_3878),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_3765),
.B(n_3773),
.Y(n_3966)
);

OR2x2_ASAP7_75t_L g3967 ( 
.A(n_3849),
.B(n_3604),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3854),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_3859),
.B(n_3678),
.Y(n_3969)
);

INVx3_ASAP7_75t_L g3970 ( 
.A(n_3834),
.Y(n_3970)
);

INVx3_ASAP7_75t_L g3971 ( 
.A(n_3834),
.Y(n_3971)
);

AND2x2_ASAP7_75t_L g3972 ( 
.A(n_3831),
.B(n_3669),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3864),
.B(n_3669),
.Y(n_3973)
);

AND2x2_ASAP7_75t_L g3974 ( 
.A(n_3867),
.B(n_3698),
.Y(n_3974)
);

HB1xp67_ASAP7_75t_L g3975 ( 
.A(n_3879),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_3886),
.Y(n_3976)
);

OR2x2_ASAP7_75t_L g3977 ( 
.A(n_3874),
.B(n_3543),
.Y(n_3977)
);

BUFx6f_ASAP7_75t_L g3978 ( 
.A(n_3736),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3812),
.B(n_3742),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3879),
.Y(n_3980)
);

INVx2_ASAP7_75t_L g3981 ( 
.A(n_3886),
.Y(n_3981)
);

OR2x2_ASAP7_75t_L g3982 ( 
.A(n_3824),
.B(n_3543),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3813),
.B(n_3709),
.Y(n_3983)
);

NOR2x1p5_ASAP7_75t_L g3984 ( 
.A(n_3736),
.B(n_3649),
.Y(n_3984)
);

AND2x2_ASAP7_75t_L g3985 ( 
.A(n_3814),
.B(n_3698),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3769),
.B(n_3642),
.Y(n_3986)
);

AND2x2_ASAP7_75t_L g3987 ( 
.A(n_3777),
.B(n_3642),
.Y(n_3987)
);

INVxp67_ASAP7_75t_L g3988 ( 
.A(n_3813),
.Y(n_3988)
);

INVx1_ASAP7_75t_L g3989 ( 
.A(n_3850),
.Y(n_3989)
);

AND2x4_ASAP7_75t_L g3990 ( 
.A(n_3761),
.B(n_3653),
.Y(n_3990)
);

INVx2_ASAP7_75t_L g3991 ( 
.A(n_3832),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3850),
.Y(n_3992)
);

INVx1_ASAP7_75t_SL g3993 ( 
.A(n_3738),
.Y(n_3993)
);

AND2x2_ASAP7_75t_L g3994 ( 
.A(n_3779),
.B(n_3642),
.Y(n_3994)
);

HB1xp67_ASAP7_75t_L g3995 ( 
.A(n_3809),
.Y(n_3995)
);

AND2x2_ASAP7_75t_L g3996 ( 
.A(n_3834),
.B(n_3599),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3851),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3894),
.B(n_3599),
.Y(n_3998)
);

BUFx2_ASAP7_75t_L g3999 ( 
.A(n_3738),
.Y(n_3999)
);

HB1xp67_ASAP7_75t_L g4000 ( 
.A(n_3851),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3891),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3891),
.Y(n_4002)
);

BUFx2_ASAP7_75t_L g4003 ( 
.A(n_3738),
.Y(n_4003)
);

BUFx2_ASAP7_75t_L g4004 ( 
.A(n_3894),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3806),
.B(n_3740),
.Y(n_4005)
);

INVx2_ASAP7_75t_L g4006 ( 
.A(n_3870),
.Y(n_4006)
);

BUFx2_ASAP7_75t_L g4007 ( 
.A(n_3894),
.Y(n_4007)
);

BUFx2_ASAP7_75t_L g4008 ( 
.A(n_3861),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3804),
.B(n_3612),
.Y(n_4009)
);

AOI22xp33_ASAP7_75t_SL g4010 ( 
.A1(n_3848),
.A2(n_3715),
.B1(n_3580),
.B2(n_3617),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_3817),
.B(n_3693),
.Y(n_4011)
);

INVx3_ASAP7_75t_L g4012 ( 
.A(n_3788),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3877),
.Y(n_4013)
);

OR2x2_ASAP7_75t_L g4014 ( 
.A(n_3775),
.B(n_3646),
.Y(n_4014)
);

INVx4_ASAP7_75t_L g4015 ( 
.A(n_3860),
.Y(n_4015)
);

AND2x2_ASAP7_75t_L g4016 ( 
.A(n_3899),
.B(n_3617),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3775),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3827),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3827),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3739),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3770),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3770),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3855),
.Y(n_4023)
);

NAND3xp33_ASAP7_75t_L g4024 ( 
.A(n_3817),
.B(n_3711),
.C(n_3729),
.Y(n_4024)
);

OR2x2_ASAP7_75t_L g4025 ( 
.A(n_3771),
.B(n_3749),
.Y(n_4025)
);

AND2x2_ASAP7_75t_L g4026 ( 
.A(n_3752),
.B(n_3638),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_3767),
.B(n_3638),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3798),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3798),
.Y(n_4029)
);

AND2x2_ASAP7_75t_L g4030 ( 
.A(n_3756),
.B(n_3638),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3811),
.Y(n_4031)
);

AND2x2_ASAP7_75t_L g4032 ( 
.A(n_3760),
.B(n_3653),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3811),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3896),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3746),
.B(n_3653),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3760),
.B(n_3778),
.Y(n_4036)
);

OR2x2_ASAP7_75t_L g4037 ( 
.A(n_3903),
.B(n_3646),
.Y(n_4037)
);

AND2x2_ASAP7_75t_L g4038 ( 
.A(n_3766),
.B(n_3566),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3800),
.B(n_3610),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3747),
.B(n_3592),
.Y(n_4040)
);

INVx3_ASAP7_75t_L g4041 ( 
.A(n_3782),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3900),
.Y(n_4042)
);

AND2x2_ASAP7_75t_L g4043 ( 
.A(n_3741),
.B(n_3619),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3838),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3838),
.Y(n_4045)
);

AND2x4_ASAP7_75t_L g4046 ( 
.A(n_3794),
.B(n_3862),
.Y(n_4046)
);

AND2x2_ASAP7_75t_L g4047 ( 
.A(n_3893),
.B(n_3619),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_3848),
.Y(n_4048)
);

AOI22xp33_ASAP7_75t_SL g4049 ( 
.A1(n_4005),
.A2(n_3750),
.B1(n_3751),
.B2(n_3863),
.Y(n_4049)
);

AOI22xp5_ASAP7_75t_L g4050 ( 
.A1(n_4048),
.A2(n_3863),
.B1(n_3841),
.B2(n_3898),
.Y(n_4050)
);

INVx2_ASAP7_75t_L g4051 ( 
.A(n_3915),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_4000),
.B(n_3868),
.Y(n_4052)
);

INVx2_ASAP7_75t_L g4053 ( 
.A(n_3970),
.Y(n_4053)
);

INVx2_ASAP7_75t_L g4054 ( 
.A(n_3970),
.Y(n_4054)
);

INVx2_ASAP7_75t_SL g4055 ( 
.A(n_3961),
.Y(n_4055)
);

AND2x4_ASAP7_75t_L g4056 ( 
.A(n_3914),
.B(n_3797),
.Y(n_4056)
);

AND2x2_ASAP7_75t_L g4057 ( 
.A(n_3986),
.B(n_3839),
.Y(n_4057)
);

AOI22xp33_ASAP7_75t_L g4058 ( 
.A1(n_4048),
.A2(n_3901),
.B1(n_3799),
.B2(n_3745),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_4023),
.B(n_3852),
.Y(n_4059)
);

BUFx2_ASAP7_75t_L g4060 ( 
.A(n_3999),
.Y(n_4060)
);

BUFx3_ASAP7_75t_L g4061 ( 
.A(n_3928),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3920),
.B(n_3801),
.Y(n_4062)
);

OR2x2_ASAP7_75t_L g4063 ( 
.A(n_3916),
.B(n_4021),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3920),
.B(n_3785),
.Y(n_4064)
);

OAI22xp5_ASAP7_75t_L g4065 ( 
.A1(n_4010),
.A2(n_3807),
.B1(n_3830),
.B2(n_3902),
.Y(n_4065)
);

AO21x2_ASAP7_75t_L g4066 ( 
.A1(n_3918),
.A2(n_3981),
.B(n_3976),
.Y(n_4066)
);

INVx2_ASAP7_75t_L g4067 ( 
.A(n_3970),
.Y(n_4067)
);

OAI21xp5_ASAP7_75t_SL g4068 ( 
.A1(n_4028),
.A2(n_3763),
.B(n_3880),
.Y(n_4068)
);

AOI22xp33_ASAP7_75t_L g4069 ( 
.A1(n_4025),
.A2(n_3745),
.B1(n_3783),
.B2(n_3750),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3975),
.B(n_3757),
.Y(n_4070)
);

BUFx2_ASAP7_75t_L g4071 ( 
.A(n_3999),
.Y(n_4071)
);

BUFx8_ASAP7_75t_L g4072 ( 
.A(n_3928),
.Y(n_4072)
);

HB1xp67_ASAP7_75t_L g4073 ( 
.A(n_3991),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3909),
.Y(n_4074)
);

AND2x4_ASAP7_75t_SL g4075 ( 
.A(n_4012),
.B(n_3762),
.Y(n_4075)
);

AOI21xp5_ASAP7_75t_L g4076 ( 
.A1(n_4011),
.A2(n_3807),
.B(n_3826),
.Y(n_4076)
);

INVx2_ASAP7_75t_L g4077 ( 
.A(n_3971),
.Y(n_4077)
);

OA21x2_ASAP7_75t_L g4078 ( 
.A1(n_4035),
.A2(n_3836),
.B(n_3837),
.Y(n_4078)
);

AOI22xp33_ASAP7_75t_L g4079 ( 
.A1(n_4025),
.A2(n_3793),
.B1(n_3818),
.B2(n_3882),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3910),
.Y(n_4080)
);

INVx4_ASAP7_75t_SL g4081 ( 
.A(n_3961),
.Y(n_4081)
);

OR2x2_ASAP7_75t_L g4082 ( 
.A(n_4022),
.B(n_3906),
.Y(n_4082)
);

AND2x6_ASAP7_75t_L g4083 ( 
.A(n_3993),
.B(n_3816),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_3986),
.B(n_3906),
.Y(n_4084)
);

BUFx3_ASAP7_75t_L g4085 ( 
.A(n_4003),
.Y(n_4085)
);

AOI22xp33_ASAP7_75t_L g4086 ( 
.A1(n_4029),
.A2(n_3768),
.B1(n_3889),
.B2(n_3865),
.Y(n_4086)
);

INVx2_ASAP7_75t_L g4087 ( 
.A(n_3971),
.Y(n_4087)
);

INVxp67_ASAP7_75t_L g4088 ( 
.A(n_3995),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3912),
.Y(n_4089)
);

O2A1O1Ixp33_ASAP7_75t_L g4090 ( 
.A1(n_4034),
.A2(n_3828),
.B(n_3844),
.C(n_3904),
.Y(n_4090)
);

INVx2_ASAP7_75t_L g4091 ( 
.A(n_3971),
.Y(n_4091)
);

AOI21xp33_ASAP7_75t_L g4092 ( 
.A1(n_4044),
.A2(n_3828),
.B(n_3884),
.Y(n_4092)
);

OAI221xp5_ASAP7_75t_L g4093 ( 
.A1(n_4045),
.A2(n_3892),
.B1(n_3869),
.B2(n_3890),
.C(n_3895),
.Y(n_4093)
);

BUFx2_ASAP7_75t_L g4094 ( 
.A(n_4003),
.Y(n_4094)
);

AOI221xp5_ASAP7_75t_L g4095 ( 
.A1(n_4031),
.A2(n_3759),
.B1(n_3885),
.B2(n_3786),
.C(n_3858),
.Y(n_4095)
);

INVx2_ASAP7_75t_L g4096 ( 
.A(n_3945),
.Y(n_4096)
);

BUFx6f_ASAP7_75t_L g4097 ( 
.A(n_3945),
.Y(n_4097)
);

INVxp67_ASAP7_75t_L g4098 ( 
.A(n_4033),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3921),
.Y(n_4099)
);

AOI21x1_ASAP7_75t_L g4100 ( 
.A1(n_4004),
.A2(n_4007),
.B(n_4036),
.Y(n_4100)
);

INVx2_ASAP7_75t_L g4101 ( 
.A(n_3945),
.Y(n_4101)
);

AND2x2_ASAP7_75t_L g4102 ( 
.A(n_3987),
.B(n_3957),
.Y(n_4102)
);

INVx2_ASAP7_75t_L g4103 ( 
.A(n_3945),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3933),
.Y(n_4104)
);

OR2x2_ASAP7_75t_L g4105 ( 
.A(n_3911),
.B(n_3786),
.Y(n_4105)
);

OAI21x1_ASAP7_75t_L g4106 ( 
.A1(n_3962),
.A2(n_3611),
.B(n_3647),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3976),
.B(n_3790),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_3936),
.Y(n_4108)
);

AO22x1_ASAP7_75t_L g4109 ( 
.A1(n_4046),
.A2(n_3764),
.B1(n_3805),
.B2(n_3810),
.Y(n_4109)
);

INVx2_ASAP7_75t_L g4110 ( 
.A(n_3978),
.Y(n_4110)
);

OAI22xp33_ASAP7_75t_L g4111 ( 
.A1(n_4024),
.A2(n_3560),
.B1(n_3559),
.B2(n_3680),
.Y(n_4111)
);

OAI21x1_ASAP7_75t_L g4112 ( 
.A1(n_3962),
.A2(n_3559),
.B(n_3632),
.Y(n_4112)
);

OAI221xp5_ASAP7_75t_L g4113 ( 
.A1(n_4020),
.A2(n_3819),
.B1(n_3847),
.B2(n_3856),
.C(n_3680),
.Y(n_4113)
);

AOI21xp5_ASAP7_75t_L g4114 ( 
.A1(n_4046),
.A2(n_3560),
.B(n_3632),
.Y(n_4114)
);

AND2x2_ASAP7_75t_L g4115 ( 
.A(n_3987),
.B(n_3661),
.Y(n_4115)
);

AO21x2_ASAP7_75t_L g4116 ( 
.A1(n_3981),
.A2(n_186),
.B(n_187),
.Y(n_4116)
);

OAI22xp5_ASAP7_75t_L g4117 ( 
.A1(n_4018),
.A2(n_3661),
.B1(n_189),
.B2(n_187),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3937),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_3957),
.B(n_188),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_3938),
.Y(n_4120)
);

AOI21xp5_ASAP7_75t_L g4121 ( 
.A1(n_4046),
.A2(n_188),
.B(n_189),
.Y(n_4121)
);

OR2x2_ASAP7_75t_L g4122 ( 
.A(n_3927),
.B(n_190),
.Y(n_4122)
);

NOR2xp33_ASAP7_75t_L g4123 ( 
.A(n_3988),
.B(n_190),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3941),
.Y(n_4124)
);

OAI21x1_ASAP7_75t_L g4125 ( 
.A1(n_3962),
.A2(n_191),
.B(n_193),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3942),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_3925),
.B(n_193),
.Y(n_4127)
);

OAI22xp5_ASAP7_75t_SL g4128 ( 
.A1(n_4019),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_4128)
);

OAI21xp33_ASAP7_75t_L g4129 ( 
.A1(n_4037),
.A2(n_194),
.B(n_195),
.Y(n_4129)
);

AOI221xp5_ASAP7_75t_L g4130 ( 
.A1(n_3989),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.C(n_200),
.Y(n_4130)
);

AOI22xp33_ASAP7_75t_L g4131 ( 
.A1(n_4036),
.A2(n_200),
.B1(n_197),
.B2(n_198),
.Y(n_4131)
);

OAI22xp5_ASAP7_75t_L g4132 ( 
.A1(n_4012),
.A2(n_4042),
.B1(n_4037),
.B2(n_3954),
.Y(n_4132)
);

INVxp33_ASAP7_75t_SL g4133 ( 
.A(n_3929),
.Y(n_4133)
);

AND4x1_ASAP7_75t_L g4134 ( 
.A(n_3994),
.B(n_203),
.C(n_201),
.D(n_202),
.Y(n_4134)
);

INVx1_ASAP7_75t_L g4135 ( 
.A(n_3944),
.Y(n_4135)
);

INVx2_ASAP7_75t_L g4136 ( 
.A(n_3978),
.Y(n_4136)
);

INVxp67_ASAP7_75t_L g4137 ( 
.A(n_3992),
.Y(n_4137)
);

AND2x4_ASAP7_75t_L g4138 ( 
.A(n_3914),
.B(n_201),
.Y(n_4138)
);

AOI21xp5_ASAP7_75t_L g4139 ( 
.A1(n_4040),
.A2(n_202),
.B(n_203),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3980),
.B(n_204),
.Y(n_4140)
);

O2A1O1Ixp33_ASAP7_75t_L g4141 ( 
.A1(n_4041),
.A2(n_207),
.B(n_205),
.C(n_206),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_3947),
.Y(n_4142)
);

OAI21x1_ASAP7_75t_L g4143 ( 
.A1(n_3930),
.A2(n_206),
.B(n_208),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_3978),
.Y(n_4144)
);

OR2x6_ASAP7_75t_L g4145 ( 
.A(n_3984),
.B(n_208),
.Y(n_4145)
);

OAI22xp5_ASAP7_75t_L g4146 ( 
.A1(n_4012),
.A2(n_212),
.B1(n_209),
.B2(n_210),
.Y(n_4146)
);

AOI22xp5_ASAP7_75t_L g4147 ( 
.A1(n_3979),
.A2(n_213),
.B1(n_210),
.B2(n_212),
.Y(n_4147)
);

AOI222xp33_ASAP7_75t_L g4148 ( 
.A1(n_3979),
.A2(n_216),
.B1(n_218),
.B2(n_213),
.C1(n_214),
.C2(n_217),
.Y(n_4148)
);

INVx2_ASAP7_75t_L g4149 ( 
.A(n_3978),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_3925),
.B(n_216),
.Y(n_4150)
);

OAI22xp5_ASAP7_75t_L g4151 ( 
.A1(n_3954),
.A2(n_222),
.B1(n_218),
.B2(n_220),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_3949),
.Y(n_4152)
);

HB1xp67_ASAP7_75t_L g4153 ( 
.A(n_3991),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3950),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_3968),
.Y(n_4155)
);

AOI22xp33_ASAP7_75t_L g4156 ( 
.A1(n_4027),
.A2(n_225),
.B1(n_220),
.B2(n_224),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3963),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_4004),
.Y(n_4158)
);

AOI22xp5_ASAP7_75t_L g4159 ( 
.A1(n_4027),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_4001),
.Y(n_4160)
);

BUFx2_ASAP7_75t_L g4161 ( 
.A(n_3907),
.Y(n_4161)
);

AOI22xp33_ASAP7_75t_SL g4162 ( 
.A1(n_4040),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_4007),
.Y(n_4163)
);

AOI22xp33_ASAP7_75t_L g4164 ( 
.A1(n_4038),
.A2(n_230),
.B1(n_227),
.B2(n_229),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_3997),
.B(n_229),
.Y(n_4165)
);

OAI21x1_ASAP7_75t_L g4166 ( 
.A1(n_3930),
.A2(n_232),
.B(n_233),
.Y(n_4166)
);

AO21x2_ASAP7_75t_L g4167 ( 
.A1(n_3964),
.A2(n_3965),
.B(n_3924),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_4002),
.Y(n_4168)
);

INVx2_ASAP7_75t_L g4169 ( 
.A(n_3930),
.Y(n_4169)
);

AND2x2_ASAP7_75t_L g4170 ( 
.A(n_3907),
.B(n_232),
.Y(n_4170)
);

BUFx12f_ASAP7_75t_L g4171 ( 
.A(n_4008),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3948),
.Y(n_4172)
);

BUFx2_ASAP7_75t_L g4173 ( 
.A(n_3994),
.Y(n_4173)
);

BUFx2_ASAP7_75t_L g4174 ( 
.A(n_3923),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_3948),
.Y(n_4175)
);

AOI22xp5_ASAP7_75t_L g4176 ( 
.A1(n_4032),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3952),
.Y(n_4177)
);

NOR2xp33_ASAP7_75t_L g4178 ( 
.A(n_4015),
.B(n_234),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_3952),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_3951),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_3969),
.Y(n_4181)
);

AOI21xp5_ASAP7_75t_L g4182 ( 
.A1(n_4006),
.A2(n_235),
.B(n_236),
.Y(n_4182)
);

BUFx6f_ASAP7_75t_L g4183 ( 
.A(n_4006),
.Y(n_4183)
);

AOI221xp5_ASAP7_75t_L g4184 ( 
.A1(n_4041),
.A2(n_240),
.B1(n_237),
.B2(n_238),
.C(n_241),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_3969),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_4074),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_4161),
.B(n_4017),
.Y(n_4187)
);

INVxp67_ASAP7_75t_SL g4188 ( 
.A(n_4062),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_4098),
.B(n_4062),
.Y(n_4189)
);

AND2x2_ASAP7_75t_L g4190 ( 
.A(n_4102),
.B(n_4173),
.Y(n_4190)
);

AOI33xp33_ASAP7_75t_L g4191 ( 
.A1(n_4049),
.A2(n_4032),
.A3(n_3964),
.B1(n_3965),
.B2(n_4030),
.B3(n_4026),
.Y(n_4191)
);

OAI321xp33_ASAP7_75t_L g4192 ( 
.A1(n_4065),
.A2(n_4026),
.A3(n_4030),
.B1(n_4013),
.B2(n_4014),
.C(n_4047),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4080),
.Y(n_4193)
);

AOI22xp33_ASAP7_75t_SL g4194 ( 
.A1(n_4065),
.A2(n_4041),
.B1(n_4047),
.B2(n_3934),
.Y(n_4194)
);

AND2x2_ASAP7_75t_L g4195 ( 
.A(n_4075),
.B(n_4039),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_4084),
.B(n_4039),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_4181),
.B(n_3958),
.Y(n_4197)
);

BUFx2_ASAP7_75t_L g4198 ( 
.A(n_4171),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4089),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4099),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_4104),
.Y(n_4201)
);

AND2x2_ASAP7_75t_L g4202 ( 
.A(n_4185),
.B(n_3958),
.Y(n_4202)
);

AND2x2_ASAP7_75t_L g4203 ( 
.A(n_4055),
.B(n_4038),
.Y(n_4203)
);

BUFx2_ASAP7_75t_L g4204 ( 
.A(n_4081),
.Y(n_4204)
);

AND2x2_ASAP7_75t_L g4205 ( 
.A(n_4057),
.B(n_3953),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4108),
.Y(n_4206)
);

INVx2_ASAP7_75t_SL g4207 ( 
.A(n_4072),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_4088),
.B(n_3959),
.Y(n_4208)
);

INVx2_ASAP7_75t_L g4209 ( 
.A(n_4081),
.Y(n_4209)
);

HB1xp67_ASAP7_75t_L g4210 ( 
.A(n_4167),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4118),
.Y(n_4211)
);

NOR2xp33_ASAP7_75t_SL g4212 ( 
.A(n_4129),
.B(n_4015),
.Y(n_4212)
);

AND2x2_ASAP7_75t_L g4213 ( 
.A(n_4056),
.B(n_3953),
.Y(n_4213)
);

INVx2_ASAP7_75t_L g4214 ( 
.A(n_4061),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_4056),
.B(n_3985),
.Y(n_4215)
);

AND2x2_ASAP7_75t_SL g4216 ( 
.A(n_4134),
.B(n_3990),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_4120),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_4124),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4126),
.Y(n_4219)
);

AND2x2_ASAP7_75t_L g4220 ( 
.A(n_4158),
.B(n_3985),
.Y(n_4220)
);

AND2x2_ASAP7_75t_L g4221 ( 
.A(n_4163),
.B(n_4085),
.Y(n_4221)
);

NAND3xp33_ASAP7_75t_L g4222 ( 
.A(n_4076),
.B(n_4014),
.C(n_3982),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_4135),
.Y(n_4223)
);

A2O1A1Ixp33_ASAP7_75t_L g4224 ( 
.A1(n_4129),
.A2(n_4068),
.B(n_4050),
.C(n_4090),
.Y(n_4224)
);

HB1xp67_ASAP7_75t_L g4225 ( 
.A(n_4167),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4142),
.Y(n_4226)
);

OR2x2_ASAP7_75t_L g4227 ( 
.A(n_4063),
.B(n_3982),
.Y(n_4227)
);

INVx3_ASAP7_75t_L g4228 ( 
.A(n_4072),
.Y(n_4228)
);

INVxp67_ASAP7_75t_L g4229 ( 
.A(n_4060),
.Y(n_4229)
);

OR2x2_ASAP7_75t_L g4230 ( 
.A(n_4064),
.B(n_3983),
.Y(n_4230)
);

INVx1_ASAP7_75t_SL g4231 ( 
.A(n_4071),
.Y(n_4231)
);

OR2x2_ASAP7_75t_L g4232 ( 
.A(n_4064),
.B(n_3932),
.Y(n_4232)
);

OR2x2_ASAP7_75t_L g4233 ( 
.A(n_4082),
.B(n_3923),
.Y(n_4233)
);

INVx3_ASAP7_75t_L g4234 ( 
.A(n_4097),
.Y(n_4234)
);

HB1xp67_ASAP7_75t_L g4235 ( 
.A(n_4094),
.Y(n_4235)
);

INVx2_ASAP7_75t_L g4236 ( 
.A(n_4097),
.Y(n_4236)
);

OA21x2_ASAP7_75t_L g4237 ( 
.A1(n_4107),
.A2(n_3924),
.B(n_3919),
.Y(n_4237)
);

BUFx2_ASAP7_75t_L g4238 ( 
.A(n_4145),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4152),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4154),
.Y(n_4240)
);

INVx2_ASAP7_75t_L g4241 ( 
.A(n_4097),
.Y(n_4241)
);

AOI22xp33_ASAP7_75t_L g4242 ( 
.A1(n_4058),
.A2(n_3955),
.B1(n_4015),
.B2(n_4043),
.Y(n_4242)
);

INVx1_ASAP7_75t_SL g4243 ( 
.A(n_4083),
.Y(n_4243)
);

AND2x2_ASAP7_75t_L g4244 ( 
.A(n_4170),
.B(n_3966),
.Y(n_4244)
);

AND2x2_ASAP7_75t_L g4245 ( 
.A(n_4096),
.B(n_3966),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4155),
.Y(n_4246)
);

AOI22xp5_ASAP7_75t_L g4247 ( 
.A1(n_4050),
.A2(n_4043),
.B1(n_3972),
.B2(n_3990),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_4160),
.Y(n_4248)
);

AND2x2_ASAP7_75t_L g4249 ( 
.A(n_4101),
.B(n_3972),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_4168),
.Y(n_4250)
);

AND2x2_ASAP7_75t_L g4251 ( 
.A(n_4103),
.B(n_3973),
.Y(n_4251)
);

OAI33xp33_ASAP7_75t_L g4252 ( 
.A1(n_4128),
.A2(n_3919),
.A3(n_3977),
.B1(n_3908),
.B2(n_3922),
.B3(n_3917),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4157),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_4059),
.B(n_3934),
.Y(n_4254)
);

BUFx2_ASAP7_75t_L g4255 ( 
.A(n_4145),
.Y(n_4255)
);

INVx3_ASAP7_75t_L g4256 ( 
.A(n_4100),
.Y(n_4256)
);

AOI21xp5_ASAP7_75t_L g4257 ( 
.A1(n_4068),
.A2(n_3955),
.B(n_3990),
.Y(n_4257)
);

INVx1_ASAP7_75t_SL g4258 ( 
.A(n_4083),
.Y(n_4258)
);

INVxp67_ASAP7_75t_L g4259 ( 
.A(n_4107),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_4172),
.Y(n_4260)
);

AND2x2_ASAP7_75t_L g4261 ( 
.A(n_4110),
.B(n_3973),
.Y(n_4261)
);

BUFx6f_ASAP7_75t_L g4262 ( 
.A(n_4138),
.Y(n_4262)
);

OR2x2_ASAP7_75t_L g4263 ( 
.A(n_4052),
.B(n_3956),
.Y(n_4263)
);

HB1xp67_ASAP7_75t_L g4264 ( 
.A(n_4174),
.Y(n_4264)
);

AND2x2_ASAP7_75t_L g4265 ( 
.A(n_4136),
.B(n_3974),
.Y(n_4265)
);

INVx5_ASAP7_75t_L g4266 ( 
.A(n_4145),
.Y(n_4266)
);

OAI22xp5_ASAP7_75t_L g4267 ( 
.A1(n_4069),
.A2(n_3908),
.B1(n_3913),
.B2(n_4009),
.Y(n_4267)
);

OA21x2_ASAP7_75t_L g4268 ( 
.A1(n_4070),
.A2(n_3926),
.B(n_3931),
.Y(n_4268)
);

INVx2_ASAP7_75t_L g4269 ( 
.A(n_4144),
.Y(n_4269)
);

HB1xp67_ASAP7_75t_L g4270 ( 
.A(n_4066),
.Y(n_4270)
);

AND2x2_ASAP7_75t_L g4271 ( 
.A(n_4149),
.B(n_3974),
.Y(n_4271)
);

OR2x2_ASAP7_75t_L g4272 ( 
.A(n_4180),
.B(n_4059),
.Y(n_4272)
);

AND2x2_ASAP7_75t_L g4273 ( 
.A(n_4127),
.B(n_3935),
.Y(n_4273)
);

HB1xp67_ASAP7_75t_L g4274 ( 
.A(n_4066),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4175),
.Y(n_4275)
);

AND2x4_ASAP7_75t_L g4276 ( 
.A(n_4051),
.B(n_3931),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4177),
.Y(n_4277)
);

NOR2xp33_ASAP7_75t_L g4278 ( 
.A(n_4133),
.B(n_4009),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4179),
.Y(n_4279)
);

AOI21x1_ASAP7_75t_L g4280 ( 
.A1(n_4119),
.A2(n_3926),
.B(n_3996),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4116),
.Y(n_4281)
);

NAND3xp33_ASAP7_75t_L g4282 ( 
.A(n_4079),
.B(n_3922),
.C(n_3917),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4116),
.Y(n_4283)
);

AND2x2_ASAP7_75t_L g4284 ( 
.A(n_4150),
.B(n_3935),
.Y(n_4284)
);

INVx1_ASAP7_75t_SL g4285 ( 
.A(n_4083),
.Y(n_4285)
);

OAI221xp5_ASAP7_75t_L g4286 ( 
.A1(n_4134),
.A2(n_3998),
.B1(n_3996),
.B2(n_3977),
.C(n_4016),
.Y(n_4286)
);

INVx3_ASAP7_75t_L g4287 ( 
.A(n_4138),
.Y(n_4287)
);

NOR2x1_ASAP7_75t_SL g4288 ( 
.A(n_4132),
.B(n_3913),
.Y(n_4288)
);

INVx4_ASAP7_75t_L g4289 ( 
.A(n_4083),
.Y(n_4289)
);

AND2x2_ASAP7_75t_L g4290 ( 
.A(n_4053),
.B(n_4016),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4137),
.Y(n_4291)
);

OR2x2_ASAP7_75t_L g4292 ( 
.A(n_4132),
.B(n_3955),
.Y(n_4292)
);

AND2x2_ASAP7_75t_L g4293 ( 
.A(n_4054),
.B(n_3943),
.Y(n_4293)
);

INVx3_ASAP7_75t_L g4294 ( 
.A(n_4183),
.Y(n_4294)
);

AOI22xp33_ASAP7_75t_L g4295 ( 
.A1(n_4095),
.A2(n_3998),
.B1(n_3960),
.B2(n_3940),
.Y(n_4295)
);

INVx2_ASAP7_75t_L g4296 ( 
.A(n_4183),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4073),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4153),
.Y(n_4298)
);

OAI211xp5_ASAP7_75t_SL g4299 ( 
.A1(n_4092),
.A2(n_3960),
.B(n_3967),
.C(n_3940),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4140),
.Y(n_4300)
);

AND2x4_ASAP7_75t_L g4301 ( 
.A(n_4067),
.B(n_3939),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4140),
.Y(n_4302)
);

INVx5_ASAP7_75t_L g4303 ( 
.A(n_4183),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_4105),
.B(n_3939),
.Y(n_4304)
);

OR2x2_ASAP7_75t_L g4305 ( 
.A(n_4122),
.B(n_3946),
.Y(n_4305)
);

AND2x2_ASAP7_75t_L g4306 ( 
.A(n_4077),
.B(n_4087),
.Y(n_4306)
);

INVx2_ASAP7_75t_L g4307 ( 
.A(n_4091),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_4216),
.B(n_4078),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4235),
.Y(n_4309)
);

INVx2_ASAP7_75t_L g4310 ( 
.A(n_4262),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4224),
.B(n_4078),
.Y(n_4311)
);

INVx2_ASAP7_75t_L g4312 ( 
.A(n_4262),
.Y(n_4312)
);

INVx1_ASAP7_75t_SL g4313 ( 
.A(n_4204),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_4235),
.Y(n_4314)
);

AND2x2_ASAP7_75t_L g4315 ( 
.A(n_4198),
.B(n_4178),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4264),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4264),
.Y(n_4317)
);

INVx3_ASAP7_75t_L g4318 ( 
.A(n_4262),
.Y(n_4318)
);

OR2x2_ASAP7_75t_L g4319 ( 
.A(n_4189),
.B(n_4165),
.Y(n_4319)
);

AND2x2_ASAP7_75t_L g4320 ( 
.A(n_4190),
.B(n_4169),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_4287),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4260),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4275),
.Y(n_4323)
);

OR2x2_ASAP7_75t_L g4324 ( 
.A(n_4189),
.B(n_4159),
.Y(n_4324)
);

AND2x4_ASAP7_75t_L g4325 ( 
.A(n_4266),
.B(n_4125),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4277),
.Y(n_4326)
);

BUFx2_ASAP7_75t_L g4327 ( 
.A(n_4287),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_SL g4328 ( 
.A(n_4216),
.B(n_4139),
.Y(n_4328)
);

AND2x2_ASAP7_75t_L g4329 ( 
.A(n_4238),
.B(n_4115),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_4259),
.B(n_4123),
.Y(n_4330)
);

INVx3_ASAP7_75t_L g4331 ( 
.A(n_4228),
.Y(n_4331)
);

INVxp67_ASAP7_75t_L g4332 ( 
.A(n_4212),
.Y(n_4332)
);

AND2x2_ASAP7_75t_L g4333 ( 
.A(n_4255),
.B(n_4278),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_4259),
.B(n_4159),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_4209),
.Y(n_4335)
);

INVx2_ASAP7_75t_L g4336 ( 
.A(n_4303),
.Y(n_4336)
);

BUFx2_ASAP7_75t_L g4337 ( 
.A(n_4266),
.Y(n_4337)
);

OR2x2_ASAP7_75t_L g4338 ( 
.A(n_4233),
.B(n_4176),
.Y(n_4338)
);

AND2x2_ASAP7_75t_L g4339 ( 
.A(n_4278),
.B(n_4092),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4279),
.Y(n_4340)
);

AND2x2_ASAP7_75t_L g4341 ( 
.A(n_4214),
.B(n_4143),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_4188),
.B(n_4086),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_4188),
.B(n_4176),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_4213),
.B(n_4166),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_4191),
.B(n_4147),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4186),
.Y(n_4346)
);

AND2x2_ASAP7_75t_L g4347 ( 
.A(n_4205),
.B(n_4162),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_4195),
.B(n_4121),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4193),
.Y(n_4349)
);

AND2x2_ASAP7_75t_L g4350 ( 
.A(n_4215),
.B(n_3946),
.Y(n_4350)
);

OR2x2_ASAP7_75t_L g4351 ( 
.A(n_4272),
.B(n_4164),
.Y(n_4351)
);

AND2x2_ASAP7_75t_L g4352 ( 
.A(n_4288),
.B(n_4182),
.Y(n_4352)
);

AND2x4_ASAP7_75t_L g4353 ( 
.A(n_4266),
.B(n_4147),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4199),
.Y(n_4354)
);

AND2x4_ASAP7_75t_L g4355 ( 
.A(n_4266),
.B(n_4231),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_L g4356 ( 
.A(n_4231),
.B(n_4184),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4200),
.Y(n_4357)
);

INVx2_ASAP7_75t_L g4358 ( 
.A(n_4303),
.Y(n_4358)
);

OR2x2_ASAP7_75t_L g4359 ( 
.A(n_4304),
.B(n_4117),
.Y(n_4359)
);

NOR2x1_ASAP7_75t_L g4360 ( 
.A(n_4289),
.B(n_4141),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4201),
.Y(n_4361)
);

OR2x2_ASAP7_75t_L g4362 ( 
.A(n_4304),
.B(n_4117),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_SL g4363 ( 
.A(n_4212),
.B(n_4151),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4206),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_4229),
.B(n_4148),
.Y(n_4365)
);

AND2x2_ASAP7_75t_L g4366 ( 
.A(n_4244),
.B(n_4151),
.Y(n_4366)
);

NOR2x1p5_ASAP7_75t_L g4367 ( 
.A(n_4228),
.B(n_4109),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4211),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_L g4369 ( 
.A(n_4229),
.B(n_4148),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4217),
.Y(n_4370)
);

HB1xp67_ASAP7_75t_L g4371 ( 
.A(n_4270),
.Y(n_4371)
);

INVxp67_ASAP7_75t_L g4372 ( 
.A(n_4286),
.Y(n_4372)
);

OR2x2_ASAP7_75t_L g4373 ( 
.A(n_4305),
.B(n_4156),
.Y(n_4373)
);

INVx4_ASAP7_75t_L g4374 ( 
.A(n_4207),
.Y(n_4374)
);

AND2x4_ASAP7_75t_L g4375 ( 
.A(n_4221),
.B(n_4249),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4218),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4219),
.Y(n_4377)
);

AOI22xp33_ASAP7_75t_L g4378 ( 
.A1(n_4194),
.A2(n_4093),
.B1(n_4130),
.B2(n_4128),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_4281),
.B(n_4146),
.Y(n_4379)
);

AND2x4_ASAP7_75t_L g4380 ( 
.A(n_4236),
.B(n_4106),
.Y(n_4380)
);

OR2x2_ASAP7_75t_L g4381 ( 
.A(n_4232),
.B(n_4114),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_4283),
.B(n_4146),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4223),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4303),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4226),
.Y(n_4385)
);

NAND2xp5_ASAP7_75t_L g4386 ( 
.A(n_4300),
.B(n_3967),
.Y(n_4386)
);

OR2x2_ASAP7_75t_L g4387 ( 
.A(n_4263),
.B(n_4111),
.Y(n_4387)
);

OR2x2_ASAP7_75t_L g4388 ( 
.A(n_4230),
.B(n_4113),
.Y(n_4388)
);

AND2x2_ASAP7_75t_L g4389 ( 
.A(n_4273),
.B(n_4112),
.Y(n_4389)
);

AND2x2_ASAP7_75t_L g4390 ( 
.A(n_4284),
.B(n_4131),
.Y(n_4390)
);

AND2x2_ASAP7_75t_L g4391 ( 
.A(n_4196),
.B(n_237),
.Y(n_4391)
);

AND2x2_ASAP7_75t_L g4392 ( 
.A(n_4187),
.B(n_238),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4239),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_L g4394 ( 
.A(n_4302),
.B(n_241),
.Y(n_4394)
);

INVx2_ASAP7_75t_L g4395 ( 
.A(n_4303),
.Y(n_4395)
);

OR2x2_ASAP7_75t_L g4396 ( 
.A(n_4208),
.B(n_242),
.Y(n_4396)
);

NAND2xp5_ASAP7_75t_SL g4397 ( 
.A(n_4194),
.B(n_243),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_4295),
.B(n_244),
.Y(n_4398)
);

NAND2xp5_ASAP7_75t_L g4399 ( 
.A(n_4295),
.B(n_244),
.Y(n_4399)
);

AND2x2_ASAP7_75t_SL g4400 ( 
.A(n_4289),
.B(n_245),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4240),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4246),
.Y(n_4402)
);

AND2x2_ASAP7_75t_L g4403 ( 
.A(n_4251),
.B(n_245),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_4248),
.B(n_246),
.Y(n_4404)
);

OR2x2_ASAP7_75t_L g4405 ( 
.A(n_4208),
.B(n_246),
.Y(n_4405)
);

INVx1_ASAP7_75t_SL g4406 ( 
.A(n_4243),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4250),
.Y(n_4407)
);

NAND2x1p5_ASAP7_75t_L g4408 ( 
.A(n_4294),
.B(n_248),
.Y(n_4408)
);

BUFx2_ASAP7_75t_L g4409 ( 
.A(n_4355),
.Y(n_4409)
);

NOR2x1_ASAP7_75t_L g4410 ( 
.A(n_4397),
.B(n_4286),
.Y(n_4410)
);

AND2x2_ASAP7_75t_L g4411 ( 
.A(n_4331),
.B(n_4290),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4371),
.Y(n_4412)
);

INVx2_ASAP7_75t_L g4413 ( 
.A(n_4374),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4309),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_4378),
.B(n_4253),
.Y(n_4415)
);

AND2x2_ASAP7_75t_SL g4416 ( 
.A(n_4311),
.B(n_4242),
.Y(n_4416)
);

NAND4xp75_ASAP7_75t_L g4417 ( 
.A(n_4311),
.B(n_4257),
.C(n_4237),
.D(n_4268),
.Y(n_4417)
);

AND2x2_ASAP7_75t_L g4418 ( 
.A(n_4331),
.B(n_4243),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_4372),
.B(n_4291),
.Y(n_4419)
);

NAND4xp75_ASAP7_75t_SL g4420 ( 
.A(n_4333),
.B(n_4237),
.C(n_4268),
.D(n_4280),
.Y(n_4420)
);

NOR2xp33_ASAP7_75t_L g4421 ( 
.A(n_4374),
.B(n_4400),
.Y(n_4421)
);

BUFx2_ASAP7_75t_SL g4422 ( 
.A(n_4355),
.Y(n_4422)
);

BUFx2_ASAP7_75t_L g4423 ( 
.A(n_4327),
.Y(n_4423)
);

INVx2_ASAP7_75t_SL g4424 ( 
.A(n_4318),
.Y(n_4424)
);

NAND4xp75_ASAP7_75t_L g4425 ( 
.A(n_4360),
.B(n_4308),
.C(n_4342),
.D(n_4328),
.Y(n_4425)
);

INVx1_ASAP7_75t_SL g4426 ( 
.A(n_4313),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4314),
.Y(n_4427)
);

INVx2_ASAP7_75t_L g4428 ( 
.A(n_4337),
.Y(n_4428)
);

HB1xp67_ASAP7_75t_L g4429 ( 
.A(n_4313),
.Y(n_4429)
);

OR2x2_ASAP7_75t_L g4430 ( 
.A(n_4338),
.B(n_4267),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_L g4431 ( 
.A(n_4398),
.B(n_4258),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4375),
.B(n_4258),
.Y(n_4432)
);

NOR2x1_ASAP7_75t_SL g4433 ( 
.A(n_4363),
.B(n_4222),
.Y(n_4433)
);

INVx3_ASAP7_75t_L g4434 ( 
.A(n_4318),
.Y(n_4434)
);

INVx1_ASAP7_75t_SL g4435 ( 
.A(n_4406),
.Y(n_4435)
);

XNOR2xp5_ASAP7_75t_L g4436 ( 
.A(n_4367),
.B(n_4267),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4375),
.B(n_4285),
.Y(n_4437)
);

INVx2_ASAP7_75t_L g4438 ( 
.A(n_4408),
.Y(n_4438)
);

NOR3xp33_ASAP7_75t_SL g4439 ( 
.A(n_4342),
.B(n_4192),
.C(n_4282),
.Y(n_4439)
);

NOR2xp33_ASAP7_75t_L g4440 ( 
.A(n_4315),
.B(n_4285),
.Y(n_4440)
);

INVx2_ASAP7_75t_L g4441 ( 
.A(n_4408),
.Y(n_4441)
);

AND2x2_ASAP7_75t_L g4442 ( 
.A(n_4366),
.B(n_4261),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_4310),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_4316),
.Y(n_4444)
);

INVx2_ASAP7_75t_L g4445 ( 
.A(n_4312),
.Y(n_4445)
);

NAND4xp75_ASAP7_75t_L g4446 ( 
.A(n_4343),
.B(n_4257),
.C(n_4345),
.D(n_4352),
.Y(n_4446)
);

INVx4_ASAP7_75t_L g4447 ( 
.A(n_4336),
.Y(n_4447)
);

AND2x2_ASAP7_75t_L g4448 ( 
.A(n_4329),
.B(n_4344),
.Y(n_4448)
);

NOR2xp33_ASAP7_75t_L g4449 ( 
.A(n_4396),
.B(n_4241),
.Y(n_4449)
);

INVx1_ASAP7_75t_L g4450 ( 
.A(n_4317),
.Y(n_4450)
);

NOR2xp33_ASAP7_75t_L g4451 ( 
.A(n_4405),
.B(n_4192),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4398),
.B(n_4269),
.Y(n_4452)
);

AND2x2_ASAP7_75t_L g4453 ( 
.A(n_4320),
.B(n_4265),
.Y(n_4453)
);

AND4x1_ASAP7_75t_L g4454 ( 
.A(n_4399),
.B(n_4242),
.C(n_4247),
.D(n_4252),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4322),
.Y(n_4455)
);

AND2x2_ASAP7_75t_L g4456 ( 
.A(n_4332),
.B(n_4271),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4323),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_4399),
.B(n_4254),
.Y(n_4458)
);

NOR2xp33_ASAP7_75t_L g4459 ( 
.A(n_4339),
.B(n_4234),
.Y(n_4459)
);

NAND4xp75_ASAP7_75t_L g4460 ( 
.A(n_4343),
.B(n_4298),
.C(n_4297),
.D(n_4254),
.Y(n_4460)
);

HB1xp67_ASAP7_75t_L g4461 ( 
.A(n_4353),
.Y(n_4461)
);

XNOR2xp5_ASAP7_75t_L g4462 ( 
.A(n_4347),
.B(n_4203),
.Y(n_4462)
);

NAND4xp75_ASAP7_75t_SL g4463 ( 
.A(n_4348),
.B(n_4306),
.C(n_4220),
.D(n_4245),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_4345),
.B(n_4406),
.Y(n_4464)
);

INVxp67_ASAP7_75t_SL g4465 ( 
.A(n_4353),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4365),
.B(n_4256),
.Y(n_4466)
);

XOR2x2_ASAP7_75t_L g4467 ( 
.A(n_4365),
.B(n_4292),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4326),
.Y(n_4468)
);

NOR2x1_ASAP7_75t_L g4469 ( 
.A(n_4358),
.B(n_4256),
.Y(n_4469)
);

NOR3xp33_ASAP7_75t_L g4470 ( 
.A(n_4369),
.B(n_4252),
.C(n_4234),
.Y(n_4470)
);

INVxp67_ASAP7_75t_L g4471 ( 
.A(n_4392),
.Y(n_4471)
);

XOR2x2_ASAP7_75t_L g4472 ( 
.A(n_4369),
.B(n_4197),
.Y(n_4472)
);

INVx3_ASAP7_75t_L g4473 ( 
.A(n_4321),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4340),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_4356),
.B(n_4296),
.Y(n_4475)
);

XOR2xp5_ASAP7_75t_L g4476 ( 
.A(n_4351),
.B(n_4202),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_L g4477 ( 
.A(n_4356),
.B(n_4307),
.Y(n_4477)
);

NAND4xp75_ASAP7_75t_L g4478 ( 
.A(n_4334),
.B(n_4293),
.C(n_4274),
.D(n_4270),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_4334),
.B(n_4324),
.Y(n_4479)
);

INVx2_ASAP7_75t_SL g4480 ( 
.A(n_4325),
.Y(n_4480)
);

AND2x2_ASAP7_75t_L g4481 ( 
.A(n_4335),
.B(n_4294),
.Y(n_4481)
);

INVx2_ASAP7_75t_L g4482 ( 
.A(n_4384),
.Y(n_4482)
);

INVx4_ASAP7_75t_L g4483 ( 
.A(n_4395),
.Y(n_4483)
);

XNOR2xp5_ASAP7_75t_L g4484 ( 
.A(n_4390),
.B(n_4227),
.Y(n_4484)
);

INVx2_ASAP7_75t_L g4485 ( 
.A(n_4325),
.Y(n_4485)
);

OAI22xp5_ASAP7_75t_L g4486 ( 
.A1(n_4359),
.A2(n_4274),
.B1(n_4225),
.B2(n_4210),
.Y(n_4486)
);

NAND3xp33_ASAP7_75t_SL g4487 ( 
.A(n_4362),
.B(n_4225),
.C(n_4210),
.Y(n_4487)
);

NAND4xp75_ASAP7_75t_SL g4488 ( 
.A(n_4341),
.B(n_4299),
.C(n_4276),
.D(n_4301),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4391),
.B(n_4276),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_4379),
.B(n_4301),
.Y(n_4490)
);

INVx2_ASAP7_75t_L g4491 ( 
.A(n_4350),
.Y(n_4491)
);

XNOR2x2_ASAP7_75t_L g4492 ( 
.A(n_4379),
.B(n_4382),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4346),
.Y(n_4493)
);

INVx2_ASAP7_75t_L g4494 ( 
.A(n_4403),
.Y(n_4494)
);

AND2x2_ASAP7_75t_L g4495 ( 
.A(n_4389),
.B(n_4299),
.Y(n_4495)
);

INVx2_ASAP7_75t_SL g4496 ( 
.A(n_4380),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4349),
.Y(n_4497)
);

AND2x2_ASAP7_75t_L g4498 ( 
.A(n_4373),
.B(n_248),
.Y(n_4498)
);

NAND4xp75_ASAP7_75t_SL g4499 ( 
.A(n_4330),
.B(n_251),
.C(n_249),
.D(n_250),
.Y(n_4499)
);

BUFx2_ASAP7_75t_L g4500 ( 
.A(n_4404),
.Y(n_4500)
);

AND2x4_ASAP7_75t_SL g4501 ( 
.A(n_4354),
.B(n_249),
.Y(n_4501)
);

XOR2xp5_ASAP7_75t_L g4502 ( 
.A(n_4388),
.B(n_250),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_L g4503 ( 
.A(n_4382),
.B(n_251),
.Y(n_4503)
);

AOI21xp5_ASAP7_75t_L g4504 ( 
.A1(n_4330),
.A2(n_252),
.B(n_253),
.Y(n_4504)
);

BUFx3_ASAP7_75t_L g4505 ( 
.A(n_4357),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_L g4506 ( 
.A(n_4394),
.B(n_253),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_L g4507 ( 
.A(n_4465),
.B(n_4394),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4492),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4429),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4461),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_4426),
.B(n_4319),
.Y(n_4511)
);

AND2x2_ASAP7_75t_L g4512 ( 
.A(n_4442),
.B(n_4361),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4426),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4435),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4435),
.Y(n_4515)
);

AND2x4_ASAP7_75t_L g4516 ( 
.A(n_4409),
.B(n_4480),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_4423),
.Y(n_4517)
);

INVx2_ASAP7_75t_L g4518 ( 
.A(n_4434),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4422),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4412),
.Y(n_4520)
);

INVxp67_ASAP7_75t_L g4521 ( 
.A(n_4421),
.Y(n_4521)
);

INVx2_ASAP7_75t_L g4522 ( 
.A(n_4434),
.Y(n_4522)
);

NAND2x1_ASAP7_75t_L g4523 ( 
.A(n_4410),
.B(n_4380),
.Y(n_4523)
);

NAND2xp5_ASAP7_75t_L g4524 ( 
.A(n_4416),
.B(n_4404),
.Y(n_4524)
);

HB1xp67_ASAP7_75t_SL g4525 ( 
.A(n_4502),
.Y(n_4525)
);

OR2x2_ASAP7_75t_L g4526 ( 
.A(n_4431),
.B(n_4387),
.Y(n_4526)
);

OR2x2_ASAP7_75t_L g4527 ( 
.A(n_4431),
.B(n_4381),
.Y(n_4527)
);

INVx1_ASAP7_75t_L g4528 ( 
.A(n_4414),
.Y(n_4528)
);

AND2x2_ASAP7_75t_L g4529 ( 
.A(n_4413),
.B(n_4364),
.Y(n_4529)
);

NOR2x1_ASAP7_75t_L g4530 ( 
.A(n_4425),
.B(n_4368),
.Y(n_4530)
);

INVxp67_ASAP7_75t_L g4531 ( 
.A(n_4433),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4448),
.B(n_4370),
.Y(n_4532)
);

AOI21xp5_ASAP7_75t_L g4533 ( 
.A1(n_4467),
.A2(n_4377),
.B(n_4376),
.Y(n_4533)
);

OAI21xp5_ASAP7_75t_SL g4534 ( 
.A1(n_4454),
.A2(n_4385),
.B(n_4383),
.Y(n_4534)
);

OR2x2_ASAP7_75t_L g4535 ( 
.A(n_4464),
.B(n_4475),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4427),
.Y(n_4536)
);

OAI21xp33_ASAP7_75t_L g4537 ( 
.A1(n_4439),
.A2(n_4401),
.B(n_4393),
.Y(n_4537)
);

NOR2xp33_ASAP7_75t_L g4538 ( 
.A(n_4438),
.B(n_4402),
.Y(n_4538)
);

OR2x2_ASAP7_75t_L g4539 ( 
.A(n_4464),
.B(n_4407),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4432),
.B(n_4386),
.Y(n_4540)
);

NOR2xp33_ASAP7_75t_L g4541 ( 
.A(n_4441),
.B(n_4440),
.Y(n_4541)
);

BUFx2_ASAP7_75t_L g4542 ( 
.A(n_4469),
.Y(n_4542)
);

OR2x6_ASAP7_75t_L g4543 ( 
.A(n_4504),
.B(n_4386),
.Y(n_4543)
);

BUFx2_ASAP7_75t_L g4544 ( 
.A(n_4447),
.Y(n_4544)
);

AND2x4_ASAP7_75t_L g4545 ( 
.A(n_4485),
.B(n_254),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4428),
.B(n_255),
.Y(n_4546)
);

AOI22xp5_ASAP7_75t_L g4547 ( 
.A1(n_4470),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4444),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4450),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4437),
.B(n_257),
.Y(n_4550)
);

AND2x2_ASAP7_75t_L g4551 ( 
.A(n_4411),
.B(n_258),
.Y(n_4551)
);

NAND3xp33_ASAP7_75t_SL g4552 ( 
.A(n_4504),
.B(n_4451),
.C(n_4430),
.Y(n_4552)
);

OR2x2_ASAP7_75t_L g4553 ( 
.A(n_4475),
.B(n_258),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_4473),
.B(n_259),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4482),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_4494),
.Y(n_4556)
);

AND2x4_ASAP7_75t_L g4557 ( 
.A(n_4418),
.B(n_260),
.Y(n_4557)
);

AND2x2_ASAP7_75t_L g4558 ( 
.A(n_4453),
.B(n_260),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4456),
.Y(n_4559)
);

AND2x2_ASAP7_75t_L g4560 ( 
.A(n_4489),
.B(n_261),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_SL g4561 ( 
.A(n_4436),
.B(n_261),
.Y(n_4561)
);

NOR2xp33_ASAP7_75t_L g4562 ( 
.A(n_4471),
.B(n_262),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4459),
.B(n_262),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4473),
.Y(n_4564)
);

NAND2xp5_ASAP7_75t_L g4565 ( 
.A(n_4424),
.B(n_4484),
.Y(n_4565)
);

AND2x2_ASAP7_75t_L g4566 ( 
.A(n_4481),
.B(n_263),
.Y(n_4566)
);

AND2x2_ASAP7_75t_L g4567 ( 
.A(n_4498),
.B(n_263),
.Y(n_4567)
);

AND2x2_ASAP7_75t_L g4568 ( 
.A(n_4491),
.B(n_264),
.Y(n_4568)
);

NOR2xp33_ASAP7_75t_L g4569 ( 
.A(n_4479),
.B(n_265),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4490),
.Y(n_4570)
);

AND2x4_ASAP7_75t_SL g4571 ( 
.A(n_4447),
.B(n_265),
.Y(n_4571)
);

OR2x2_ASAP7_75t_L g4572 ( 
.A(n_4477),
.B(n_267),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4490),
.Y(n_4573)
);

NOR2xp33_ASAP7_75t_L g4574 ( 
.A(n_4479),
.B(n_4452),
.Y(n_4574)
);

AND2x4_ASAP7_75t_L g4575 ( 
.A(n_4483),
.B(n_267),
.Y(n_4575)
);

NAND2x2_ASAP7_75t_L g4576 ( 
.A(n_4505),
.B(n_268),
.Y(n_4576)
);

NAND2x1_ASAP7_75t_L g4577 ( 
.A(n_4496),
.B(n_4483),
.Y(n_4577)
);

INVx2_ASAP7_75t_SL g4578 ( 
.A(n_4501),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4443),
.Y(n_4579)
);

OR2x2_ASAP7_75t_L g4580 ( 
.A(n_4477),
.B(n_268),
.Y(n_4580)
);

AND2x4_ASAP7_75t_L g4581 ( 
.A(n_4445),
.B(n_270),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_4462),
.B(n_270),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4455),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4457),
.Y(n_4584)
);

NOR2x1_ASAP7_75t_L g4585 ( 
.A(n_4417),
.B(n_272),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4468),
.Y(n_4586)
);

AND2x2_ASAP7_75t_L g4587 ( 
.A(n_4449),
.B(n_273),
.Y(n_4587)
);

AOI21xp33_ASAP7_75t_SL g4588 ( 
.A1(n_4466),
.A2(n_273),
.B(n_274),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4474),
.Y(n_4589)
);

AND2x2_ASAP7_75t_L g4590 ( 
.A(n_4500),
.B(n_274),
.Y(n_4590)
);

HB1xp67_ASAP7_75t_L g4591 ( 
.A(n_4420),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4493),
.Y(n_4592)
);

AOI21xp33_ASAP7_75t_SL g4593 ( 
.A1(n_4466),
.A2(n_275),
.B(n_277),
.Y(n_4593)
);

NOR2xp67_ASAP7_75t_L g4594 ( 
.A(n_4487),
.B(n_278),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_SL g4595 ( 
.A(n_4472),
.B(n_278),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_L g4596 ( 
.A(n_4476),
.B(n_280),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4497),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_4486),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4486),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_4419),
.B(n_280),
.Y(n_4600)
);

NAND2x1p5_ASAP7_75t_L g4601 ( 
.A(n_4577),
.B(n_4506),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4516),
.Y(n_4602)
);

AOI21xp5_ASAP7_75t_L g4603 ( 
.A1(n_4534),
.A2(n_4415),
.B(n_4503),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4510),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4510),
.Y(n_4605)
);

AO21x1_ASAP7_75t_L g4606 ( 
.A1(n_4508),
.A2(n_4503),
.B(n_4415),
.Y(n_4606)
);

OAI221xp5_ASAP7_75t_L g4607 ( 
.A1(n_4547),
.A2(n_4419),
.B1(n_4458),
.B2(n_4452),
.C(n_4495),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4509),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_L g4609 ( 
.A(n_4516),
.B(n_4460),
.Y(n_4609)
);

AOI22xp33_ASAP7_75t_L g4610 ( 
.A1(n_4508),
.A2(n_4458),
.B1(n_4488),
.B2(n_4420),
.Y(n_4610)
);

OAI21xp33_ASAP7_75t_L g4611 ( 
.A1(n_4585),
.A2(n_4506),
.B(n_4463),
.Y(n_4611)
);

OAI21xp33_ASAP7_75t_L g4612 ( 
.A1(n_4541),
.A2(n_4463),
.B(n_4446),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4509),
.Y(n_4613)
);

AOI22xp5_ASAP7_75t_L g4614 ( 
.A1(n_4552),
.A2(n_4478),
.B1(n_4488),
.B2(n_4499),
.Y(n_4614)
);

INVx2_ASAP7_75t_SL g4615 ( 
.A(n_4544),
.Y(n_4615)
);

OAI22xp5_ASAP7_75t_L g4616 ( 
.A1(n_4531),
.A2(n_4499),
.B1(n_283),
.B2(n_281),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_4519),
.B(n_282),
.Y(n_4617)
);

INVx2_ASAP7_75t_L g4618 ( 
.A(n_4571),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_L g4619 ( 
.A(n_4578),
.B(n_285),
.Y(n_4619)
);

OAI22x1_ASAP7_75t_L g4620 ( 
.A1(n_4542),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4513),
.Y(n_4621)
);

OAI22xp5_ASAP7_75t_L g4622 ( 
.A1(n_4523),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_4622)
);

OAI211xp5_ASAP7_75t_SL g4623 ( 
.A1(n_4524),
.A2(n_4537),
.B(n_4521),
.C(n_4530),
.Y(n_4623)
);

INVxp67_ASAP7_75t_L g4624 ( 
.A(n_4525),
.Y(n_4624)
);

AOI21xp5_ASAP7_75t_L g4625 ( 
.A1(n_4543),
.A2(n_288),
.B(n_290),
.Y(n_4625)
);

OAI22x1_ASAP7_75t_SL g4626 ( 
.A1(n_4514),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_4626)
);

OAI21xp33_ASAP7_75t_L g4627 ( 
.A1(n_4565),
.A2(n_291),
.B(n_292),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4515),
.Y(n_4628)
);

AOI31xp33_ASAP7_75t_L g4629 ( 
.A1(n_4595),
.A2(n_297),
.A3(n_293),
.B(n_294),
.Y(n_4629)
);

HB1xp67_ASAP7_75t_L g4630 ( 
.A(n_4575),
.Y(n_4630)
);

AOI32xp33_ASAP7_75t_L g4631 ( 
.A1(n_4574),
.A2(n_4598),
.A3(n_4599),
.B1(n_4569),
.B2(n_4561),
.Y(n_4631)
);

INVx2_ASAP7_75t_L g4632 ( 
.A(n_4575),
.Y(n_4632)
);

AOI21xp33_ASAP7_75t_L g4633 ( 
.A1(n_4543),
.A2(n_293),
.B(n_294),
.Y(n_4633)
);

BUFx3_ASAP7_75t_L g4634 ( 
.A(n_4517),
.Y(n_4634)
);

AOI22xp5_ASAP7_75t_L g4635 ( 
.A1(n_4594),
.A2(n_302),
.B1(n_299),
.B2(n_301),
.Y(n_4635)
);

INVx2_ASAP7_75t_L g4636 ( 
.A(n_4518),
.Y(n_4636)
);

AO21x1_ASAP7_75t_L g4637 ( 
.A1(n_4598),
.A2(n_299),
.B(n_301),
.Y(n_4637)
);

AND2x4_ASAP7_75t_L g4638 ( 
.A(n_4522),
.B(n_302),
.Y(n_4638)
);

AOI22xp33_ASAP7_75t_L g4639 ( 
.A1(n_4591),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4559),
.Y(n_4640)
);

AOI22xp33_ASAP7_75t_L g4641 ( 
.A1(n_4533),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_4641)
);

INVx4_ASAP7_75t_L g4642 ( 
.A(n_4581),
.Y(n_4642)
);

OAI31xp33_ASAP7_75t_L g4643 ( 
.A1(n_4535),
.A2(n_311),
.A3(n_309),
.B(n_310),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_4567),
.Y(n_4644)
);

OAI21xp5_ASAP7_75t_L g4645 ( 
.A1(n_4511),
.A2(n_4526),
.B(n_4599),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4558),
.Y(n_4646)
);

AO21x1_ASAP7_75t_L g4647 ( 
.A1(n_4588),
.A2(n_310),
.B(n_313),
.Y(n_4647)
);

AOI22xp5_ASAP7_75t_L g4648 ( 
.A1(n_4582),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_4648)
);

INVxp67_ASAP7_75t_L g4649 ( 
.A(n_4550),
.Y(n_4649)
);

NOR3xp33_ASAP7_75t_L g4650 ( 
.A(n_4507),
.B(n_314),
.C(n_316),
.Y(n_4650)
);

O2A1O1Ixp33_ASAP7_75t_L g4651 ( 
.A1(n_4593),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_4651)
);

AOI21xp5_ASAP7_75t_SL g4652 ( 
.A1(n_4557),
.A2(n_317),
.B(n_319),
.Y(n_4652)
);

INVx1_ASAP7_75t_SL g4653 ( 
.A(n_4590),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4554),
.Y(n_4654)
);

OAI21xp5_ASAP7_75t_SL g4655 ( 
.A1(n_4540),
.A2(n_319),
.B(n_320),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4512),
.Y(n_4656)
);

XOR2x2_ASAP7_75t_L g4657 ( 
.A(n_4596),
.B(n_4527),
.Y(n_4657)
);

OAI22xp33_ASAP7_75t_SL g4658 ( 
.A1(n_4576),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_4658)
);

NAND2x1p5_ASAP7_75t_L g4659 ( 
.A(n_4557),
.B(n_322),
.Y(n_4659)
);

BUFx3_ASAP7_75t_L g4660 ( 
.A(n_4566),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4551),
.Y(n_4661)
);

AOI21xp5_ASAP7_75t_L g4662 ( 
.A1(n_4546),
.A2(n_323),
.B(n_324),
.Y(n_4662)
);

INVxp67_ASAP7_75t_SL g4663 ( 
.A(n_4564),
.Y(n_4663)
);

OR2x2_ASAP7_75t_L g4664 ( 
.A(n_4539),
.B(n_4570),
.Y(n_4664)
);

NAND2x1p5_ASAP7_75t_L g4665 ( 
.A(n_4560),
.B(n_325),
.Y(n_4665)
);

OR2x2_ASAP7_75t_L g4666 ( 
.A(n_4573),
.B(n_326),
.Y(n_4666)
);

AOI31xp33_ASAP7_75t_L g4667 ( 
.A1(n_4556),
.A2(n_328),
.A3(n_326),
.B(n_327),
.Y(n_4667)
);

NAND3xp33_ASAP7_75t_L g4668 ( 
.A(n_4538),
.B(n_4520),
.C(n_4555),
.Y(n_4668)
);

OAI22xp5_ASAP7_75t_L g4669 ( 
.A1(n_4553),
.A2(n_331),
.B1(n_328),
.B2(n_330),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4545),
.Y(n_4670)
);

INVx2_ASAP7_75t_L g4671 ( 
.A(n_4545),
.Y(n_4671)
);

AOI221x1_ASAP7_75t_L g4672 ( 
.A1(n_4579),
.A2(n_332),
.B1(n_333),
.B2(n_335),
.C(n_336),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4568),
.Y(n_4673)
);

HB1xp67_ASAP7_75t_L g4674 ( 
.A(n_4581),
.Y(n_4674)
);

OAI22xp5_ASAP7_75t_L g4675 ( 
.A1(n_4572),
.A2(n_337),
.B1(n_333),
.B2(n_336),
.Y(n_4675)
);

XOR2x2_ASAP7_75t_L g4676 ( 
.A(n_4563),
.B(n_338),
.Y(n_4676)
);

AOI22xp5_ASAP7_75t_L g4677 ( 
.A1(n_4532),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.Y(n_4677)
);

OAI21xp5_ASAP7_75t_L g4678 ( 
.A1(n_4600),
.A2(n_339),
.B(n_341),
.Y(n_4678)
);

INVx2_ASAP7_75t_L g4679 ( 
.A(n_4529),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4587),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4580),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4528),
.Y(n_4682)
);

OAI22xp5_ASAP7_75t_L g4683 ( 
.A1(n_4562),
.A2(n_344),
.B1(n_341),
.B2(n_342),
.Y(n_4683)
);

OAI22xp5_ASAP7_75t_L g4684 ( 
.A1(n_4536),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.Y(n_4684)
);

OAI22xp33_ASAP7_75t_L g4685 ( 
.A1(n_4548),
.A2(n_348),
.B1(n_345),
.B2(n_347),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4630),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_4674),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_L g4688 ( 
.A(n_4602),
.B(n_4549),
.Y(n_4688)
);

NAND2xp33_ASAP7_75t_L g4689 ( 
.A(n_4631),
.B(n_4583),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_L g4690 ( 
.A(n_4615),
.B(n_4584),
.Y(n_4690)
);

OAI21xp5_ASAP7_75t_L g4691 ( 
.A1(n_4614),
.A2(n_4589),
.B(n_4586),
.Y(n_4691)
);

CKINVDCx16_ASAP7_75t_R g4692 ( 
.A(n_4660),
.Y(n_4692)
);

OR2x2_ASAP7_75t_L g4693 ( 
.A(n_4632),
.B(n_4592),
.Y(n_4693)
);

NAND3xp33_ASAP7_75t_L g4694 ( 
.A(n_4623),
.B(n_4597),
.C(n_349),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4670),
.Y(n_4695)
);

AOI222xp33_ASAP7_75t_L g4696 ( 
.A1(n_4610),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.C1(n_352),
.C2(n_353),
.Y(n_4696)
);

INVxp67_ASAP7_75t_L g4697 ( 
.A(n_4626),
.Y(n_4697)
);

OR2x2_ASAP7_75t_L g4698 ( 
.A(n_4671),
.B(n_4653),
.Y(n_4698)
);

HB1xp67_ASAP7_75t_L g4699 ( 
.A(n_4601),
.Y(n_4699)
);

OAI31xp33_ASAP7_75t_L g4700 ( 
.A1(n_4622),
.A2(n_355),
.A3(n_353),
.B(n_354),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4617),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4619),
.Y(n_4702)
);

INVx2_ASAP7_75t_L g4703 ( 
.A(n_4659),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4634),
.Y(n_4704)
);

NAND2xp5_ASAP7_75t_L g4705 ( 
.A(n_4624),
.B(n_354),
.Y(n_4705)
);

AND2x2_ASAP7_75t_L g4706 ( 
.A(n_4618),
.B(n_356),
.Y(n_4706)
);

OR2x2_ASAP7_75t_L g4707 ( 
.A(n_4642),
.B(n_356),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_4642),
.B(n_358),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4663),
.Y(n_4709)
);

NAND3xp33_ASAP7_75t_L g4710 ( 
.A(n_4631),
.B(n_358),
.C(n_359),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4656),
.Y(n_4711)
);

INVx2_ASAP7_75t_L g4712 ( 
.A(n_4665),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4638),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4638),
.Y(n_4714)
);

OAI22xp5_ASAP7_75t_L g4715 ( 
.A1(n_4641),
.A2(n_364),
.B1(n_361),
.B2(n_363),
.Y(n_4715)
);

OR2x2_ASAP7_75t_L g4716 ( 
.A(n_4661),
.B(n_361),
.Y(n_4716)
);

INVx1_ASAP7_75t_SL g4717 ( 
.A(n_4626),
.Y(n_4717)
);

INVx1_ASAP7_75t_SL g4718 ( 
.A(n_4609),
.Y(n_4718)
);

INVx2_ASAP7_75t_SL g4719 ( 
.A(n_4679),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4604),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_L g4721 ( 
.A(n_4616),
.B(n_363),
.Y(n_4721)
);

INVxp67_ASAP7_75t_L g4722 ( 
.A(n_4620),
.Y(n_4722)
);

AND2x2_ASAP7_75t_L g4723 ( 
.A(n_4646),
.B(n_365),
.Y(n_4723)
);

AOI22xp5_ASAP7_75t_L g4724 ( 
.A1(n_4606),
.A2(n_370),
.B1(n_366),
.B2(n_369),
.Y(n_4724)
);

AND2x2_ASAP7_75t_L g4725 ( 
.A(n_4644),
.B(n_369),
.Y(n_4725)
);

A2O1A1Ixp33_ASAP7_75t_L g4726 ( 
.A1(n_4633),
.A2(n_373),
.B(n_371),
.C(n_372),
.Y(n_4726)
);

AOI21xp5_ASAP7_75t_L g4727 ( 
.A1(n_4603),
.A2(n_371),
.B(n_372),
.Y(n_4727)
);

AND2x2_ASAP7_75t_L g4728 ( 
.A(n_4649),
.B(n_373),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_SL g4729 ( 
.A(n_4647),
.B(n_374),
.Y(n_4729)
);

OR2x2_ASAP7_75t_L g4730 ( 
.A(n_4636),
.B(n_374),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_4605),
.Y(n_4731)
);

OA21x2_ASAP7_75t_L g4732 ( 
.A1(n_4625),
.A2(n_376),
.B(n_377),
.Y(n_4732)
);

INVx1_ASAP7_75t_L g4733 ( 
.A(n_4608),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4680),
.B(n_376),
.Y(n_4734)
);

INVx1_ASAP7_75t_L g4735 ( 
.A(n_4613),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_4621),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4628),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4637),
.Y(n_4738)
);

CKINVDCx16_ASAP7_75t_R g4739 ( 
.A(n_4645),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4666),
.Y(n_4740)
);

INVx1_ASAP7_75t_SL g4741 ( 
.A(n_4676),
.Y(n_4741)
);

OAI21xp33_ASAP7_75t_L g4742 ( 
.A1(n_4612),
.A2(n_377),
.B(n_378),
.Y(n_4742)
);

OR2x2_ASAP7_75t_L g4743 ( 
.A(n_4664),
.B(n_379),
.Y(n_4743)
);

OR2x2_ASAP7_75t_L g4744 ( 
.A(n_4673),
.B(n_379),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4635),
.B(n_380),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_4635),
.B(n_381),
.Y(n_4746)
);

NAND2xp5_ASAP7_75t_L g4747 ( 
.A(n_4629),
.B(n_381),
.Y(n_4747)
);

AOI21xp33_ASAP7_75t_L g4748 ( 
.A1(n_4611),
.A2(n_382),
.B(n_383),
.Y(n_4748)
);

AND2x2_ASAP7_75t_L g4749 ( 
.A(n_4681),
.B(n_382),
.Y(n_4749)
);

OAI22xp5_ASAP7_75t_L g4750 ( 
.A1(n_4607),
.A2(n_383),
.B1(n_384),
.B2(n_386),
.Y(n_4750)
);

HB1xp67_ASAP7_75t_L g4751 ( 
.A(n_4640),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_L g4752 ( 
.A(n_4692),
.B(n_4655),
.Y(n_4752)
);

INVxp67_ASAP7_75t_SL g4753 ( 
.A(n_4699),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4686),
.Y(n_4754)
);

OAI22xp5_ASAP7_75t_L g4755 ( 
.A1(n_4739),
.A2(n_4639),
.B1(n_4668),
.B2(n_4648),
.Y(n_4755)
);

AOI21xp5_ASAP7_75t_L g4756 ( 
.A1(n_4689),
.A2(n_4657),
.B(n_4662),
.Y(n_4756)
);

OR2x2_ASAP7_75t_L g4757 ( 
.A(n_4717),
.B(n_4654),
.Y(n_4757)
);

INVxp33_ASAP7_75t_L g4758 ( 
.A(n_4729),
.Y(n_4758)
);

AOI322xp5_ASAP7_75t_L g4759 ( 
.A1(n_4697),
.A2(n_4738),
.A3(n_4724),
.B1(n_4722),
.B2(n_4718),
.C1(n_4741),
.C2(n_4742),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4687),
.Y(n_4760)
);

AND2x2_ASAP7_75t_L g4761 ( 
.A(n_4703),
.B(n_4678),
.Y(n_4761)
);

NOR2xp33_ASAP7_75t_L g4762 ( 
.A(n_4713),
.B(n_4627),
.Y(n_4762)
);

OAI21xp33_ASAP7_75t_L g4763 ( 
.A1(n_4724),
.A2(n_4650),
.B(n_4682),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4698),
.Y(n_4764)
);

AOI21xp33_ASAP7_75t_L g4765 ( 
.A1(n_4712),
.A2(n_4658),
.B(n_4651),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4707),
.Y(n_4766)
);

INVx2_ASAP7_75t_L g4767 ( 
.A(n_4714),
.Y(n_4767)
);

NAND2xp5_ASAP7_75t_L g4768 ( 
.A(n_4706),
.B(n_4643),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4708),
.Y(n_4769)
);

OR2x2_ASAP7_75t_L g4770 ( 
.A(n_4704),
.B(n_4693),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4751),
.Y(n_4771)
);

AND2x4_ASAP7_75t_L g4772 ( 
.A(n_4709),
.B(n_4672),
.Y(n_4772)
);

AND2x2_ASAP7_75t_L g4773 ( 
.A(n_4701),
.B(n_4652),
.Y(n_4773)
);

INVx2_ASAP7_75t_SL g4774 ( 
.A(n_4719),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4734),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4695),
.Y(n_4776)
);

INVx1_ASAP7_75t_SL g4777 ( 
.A(n_4743),
.Y(n_4777)
);

XNOR2xp5_ASAP7_75t_L g4778 ( 
.A(n_4694),
.B(n_4677),
.Y(n_4778)
);

AOI22xp33_ASAP7_75t_L g4779 ( 
.A1(n_4694),
.A2(n_4683),
.B1(n_4669),
.B2(n_4675),
.Y(n_4779)
);

NAND4xp25_ASAP7_75t_L g4780 ( 
.A(n_4691),
.B(n_4648),
.C(n_4684),
.D(n_4667),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4723),
.Y(n_4781)
);

NOR2x1_ASAP7_75t_L g4782 ( 
.A(n_4710),
.B(n_4685),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4725),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4728),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4705),
.Y(n_4785)
);

INVx2_ASAP7_75t_L g4786 ( 
.A(n_4716),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4688),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4749),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4700),
.B(n_384),
.Y(n_4789)
);

OAI31xp33_ASAP7_75t_L g4790 ( 
.A1(n_4710),
.A2(n_386),
.A3(n_387),
.B(n_389),
.Y(n_4790)
);

OAI22xp5_ASAP7_75t_SL g4791 ( 
.A1(n_4747),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.Y(n_4791)
);

INVx2_ASAP7_75t_L g4792 ( 
.A(n_4744),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4690),
.Y(n_4793)
);

OAI211xp5_ASAP7_75t_SL g4794 ( 
.A1(n_4742),
.A2(n_392),
.B(n_393),
.C(n_394),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4730),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4711),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4740),
.Y(n_4797)
);

NOR2xp33_ASAP7_75t_L g4798 ( 
.A(n_4721),
.B(n_394),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_L g4799 ( 
.A(n_4700),
.B(n_395),
.Y(n_4799)
);

INVx2_ASAP7_75t_L g4800 ( 
.A(n_4720),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4731),
.Y(n_4801)
);

INVx1_ASAP7_75t_L g4802 ( 
.A(n_4733),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_4735),
.Y(n_4803)
);

OAI311xp33_ASAP7_75t_L g4804 ( 
.A1(n_4696),
.A2(n_395),
.A3(n_396),
.B1(n_397),
.C1(n_398),
.Y(n_4804)
);

INVx2_ASAP7_75t_L g4805 ( 
.A(n_4732),
.Y(n_4805)
);

AOI211xp5_ASAP7_75t_L g4806 ( 
.A1(n_4750),
.A2(n_396),
.B(n_399),
.C(n_400),
.Y(n_4806)
);

AOI21xp33_ASAP7_75t_SL g4807 ( 
.A1(n_4732),
.A2(n_399),
.B(n_400),
.Y(n_4807)
);

AND2x4_ASAP7_75t_L g4808 ( 
.A(n_4736),
.B(n_401),
.Y(n_4808)
);

OR2x2_ASAP7_75t_L g4809 ( 
.A(n_4737),
.B(n_401),
.Y(n_4809)
);

HB1xp67_ASAP7_75t_L g4810 ( 
.A(n_4745),
.Y(n_4810)
);

OR2x2_ASAP7_75t_L g4811 ( 
.A(n_4702),
.B(n_404),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4746),
.Y(n_4812)
);

AND2x2_ASAP7_75t_L g4813 ( 
.A(n_4748),
.B(n_405),
.Y(n_4813)
);

OAI21xp5_ASAP7_75t_L g4814 ( 
.A1(n_4727),
.A2(n_405),
.B(n_407),
.Y(n_4814)
);

AOI221xp5_ASAP7_75t_L g4815 ( 
.A1(n_4755),
.A2(n_4715),
.B1(n_4726),
.B2(n_410),
.C(n_411),
.Y(n_4815)
);

INVx2_ASAP7_75t_L g4816 ( 
.A(n_4770),
.Y(n_4816)
);

O2A1O1Ixp33_ASAP7_75t_L g4817 ( 
.A1(n_4804),
.A2(n_408),
.B(n_409),
.C(n_411),
.Y(n_4817)
);

AOI211xp5_ASAP7_75t_L g4818 ( 
.A1(n_4807),
.A2(n_408),
.B(n_409),
.C(n_412),
.Y(n_4818)
);

NAND3xp33_ASAP7_75t_SL g4819 ( 
.A(n_4756),
.B(n_412),
.C(n_414),
.Y(n_4819)
);

INVx2_ASAP7_75t_L g4820 ( 
.A(n_4805),
.Y(n_4820)
);

CKINVDCx14_ASAP7_75t_R g4821 ( 
.A(n_4773),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_4759),
.B(n_415),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4753),
.Y(n_4823)
);

NOR2xp67_ASAP7_75t_L g4824 ( 
.A(n_4774),
.B(n_415),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4757),
.Y(n_4825)
);

OAI21xp33_ASAP7_75t_SL g4826 ( 
.A1(n_4759),
.A2(n_417),
.B(n_418),
.Y(n_4826)
);

AOI221xp5_ASAP7_75t_L g4827 ( 
.A1(n_4763),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.C(n_422),
.Y(n_4827)
);

AOI221xp5_ASAP7_75t_L g4828 ( 
.A1(n_4763),
.A2(n_420),
.B1(n_422),
.B2(n_423),
.C(n_424),
.Y(n_4828)
);

O2A1O1Ixp33_ASAP7_75t_L g4829 ( 
.A1(n_4790),
.A2(n_4772),
.B(n_4799),
.C(n_4789),
.Y(n_4829)
);

NAND3xp33_ASAP7_75t_L g4830 ( 
.A(n_4790),
.B(n_423),
.C(n_424),
.Y(n_4830)
);

NAND3xp33_ASAP7_75t_SL g4831 ( 
.A(n_4777),
.B(n_4758),
.C(n_4764),
.Y(n_4831)
);

AND2x2_ASAP7_75t_L g4832 ( 
.A(n_4767),
.B(n_426),
.Y(n_4832)
);

NOR3x1_ASAP7_75t_L g4833 ( 
.A(n_4780),
.B(n_426),
.C(n_427),
.Y(n_4833)
);

OR2x2_ASAP7_75t_L g4834 ( 
.A(n_4768),
.B(n_4772),
.Y(n_4834)
);

INVx1_ASAP7_75t_L g4835 ( 
.A(n_4791),
.Y(n_4835)
);

NOR2xp67_ASAP7_75t_L g4836 ( 
.A(n_4771),
.B(n_428),
.Y(n_4836)
);

NAND2xp33_ASAP7_75t_L g4837 ( 
.A(n_4782),
.B(n_431),
.Y(n_4837)
);

NAND2xp5_ASAP7_75t_L g4838 ( 
.A(n_4766),
.B(n_4762),
.Y(n_4838)
);

HB1xp67_ASAP7_75t_L g4839 ( 
.A(n_4752),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_SL g4840 ( 
.A(n_4806),
.B(n_431),
.Y(n_4840)
);

XNOR2x2_ASAP7_75t_L g4841 ( 
.A(n_4778),
.B(n_432),
.Y(n_4841)
);

NAND2xp5_ASAP7_75t_SL g4842 ( 
.A(n_4806),
.B(n_432),
.Y(n_4842)
);

NAND2xp5_ASAP7_75t_L g4843 ( 
.A(n_4775),
.B(n_433),
.Y(n_4843)
);

OAI21xp5_ASAP7_75t_SL g4844 ( 
.A1(n_4779),
.A2(n_435),
.B(n_436),
.Y(n_4844)
);

OR2x2_ASAP7_75t_L g4845 ( 
.A(n_4781),
.B(n_437),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4791),
.Y(n_4846)
);

NAND4xp25_ASAP7_75t_L g4847 ( 
.A(n_4765),
.B(n_437),
.C(n_438),
.D(n_440),
.Y(n_4847)
);

AND2x4_ASAP7_75t_L g4848 ( 
.A(n_4786),
.B(n_440),
.Y(n_4848)
);

AOI221xp5_ASAP7_75t_L g4849 ( 
.A1(n_4754),
.A2(n_441),
.B1(n_442),
.B2(n_443),
.C(n_444),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4783),
.B(n_4788),
.Y(n_4850)
);

AOI211x1_ASAP7_75t_L g4851 ( 
.A1(n_4814),
.A2(n_443),
.B(n_444),
.C(n_445),
.Y(n_4851)
);

AOI21xp5_ASAP7_75t_L g4852 ( 
.A1(n_4795),
.A2(n_445),
.B(n_446),
.Y(n_4852)
);

NOR2xp33_ASAP7_75t_L g4853 ( 
.A(n_4794),
.B(n_447),
.Y(n_4853)
);

NOR3xp33_ASAP7_75t_L g4854 ( 
.A(n_4812),
.B(n_447),
.C(n_448),
.Y(n_4854)
);

NOR2xp33_ASAP7_75t_L g4855 ( 
.A(n_4784),
.B(n_448),
.Y(n_4855)
);

AND2x2_ASAP7_75t_L g4856 ( 
.A(n_4761),
.B(n_451),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_L g4857 ( 
.A(n_4760),
.B(n_4792),
.Y(n_4857)
);

NOR2xp33_ASAP7_75t_L g4858 ( 
.A(n_4797),
.B(n_451),
.Y(n_4858)
);

NAND2xp5_ASAP7_75t_SL g4859 ( 
.A(n_4776),
.B(n_452),
.Y(n_4859)
);

INVx2_ASAP7_75t_L g4860 ( 
.A(n_4808),
.Y(n_4860)
);

NOR2xp67_ASAP7_75t_L g4861 ( 
.A(n_4809),
.B(n_4811),
.Y(n_4861)
);

AOI21xp33_ASAP7_75t_SL g4862 ( 
.A1(n_4796),
.A2(n_452),
.B(n_453),
.Y(n_4862)
);

INVx2_ASAP7_75t_L g4863 ( 
.A(n_4808),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4810),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4798),
.B(n_453),
.Y(n_4865)
);

AOI21xp5_ASAP7_75t_L g4866 ( 
.A1(n_4769),
.A2(n_454),
.B(n_455),
.Y(n_4866)
);

AOI21xp5_ASAP7_75t_L g4867 ( 
.A1(n_4831),
.A2(n_4829),
.B(n_4822),
.Y(n_4867)
);

AOI221xp5_ASAP7_75t_L g4868 ( 
.A1(n_4826),
.A2(n_4793),
.B1(n_4787),
.B2(n_4802),
.C(n_4801),
.Y(n_4868)
);

AND3x1_ASAP7_75t_L g4869 ( 
.A(n_4860),
.B(n_4800),
.C(n_4785),
.Y(n_4869)
);

INVx2_ASAP7_75t_L g4870 ( 
.A(n_4820),
.Y(n_4870)
);

NOR3xp33_ASAP7_75t_L g4871 ( 
.A(n_4819),
.B(n_4803),
.C(n_4813),
.Y(n_4871)
);

NOR3x1_ASAP7_75t_L g4872 ( 
.A(n_4844),
.B(n_454),
.C(n_456),
.Y(n_4872)
);

NAND2xp5_ASAP7_75t_SL g4873 ( 
.A(n_4824),
.B(n_4817),
.Y(n_4873)
);

AOI221xp5_ASAP7_75t_L g4874 ( 
.A1(n_4835),
.A2(n_456),
.B1(n_457),
.B2(n_458),
.C(n_459),
.Y(n_4874)
);

NOR3xp33_ASAP7_75t_L g4875 ( 
.A(n_4821),
.B(n_457),
.C(n_460),
.Y(n_4875)
);

AOI221xp5_ASAP7_75t_L g4876 ( 
.A1(n_4846),
.A2(n_462),
.B1(n_465),
.B2(n_466),
.C(n_467),
.Y(n_4876)
);

AOI221xp5_ASAP7_75t_L g4877 ( 
.A1(n_4823),
.A2(n_4830),
.B1(n_4837),
.B2(n_4815),
.C(n_4825),
.Y(n_4877)
);

AOI322xp5_ASAP7_75t_L g4878 ( 
.A1(n_4839),
.A2(n_465),
.A3(n_467),
.B1(n_469),
.B2(n_470),
.C1(n_471),
.C2(n_472),
.Y(n_4878)
);

AOI21xp5_ASAP7_75t_L g4879 ( 
.A1(n_4838),
.A2(n_469),
.B(n_470),
.Y(n_4879)
);

AOI22xp33_ASAP7_75t_L g4880 ( 
.A1(n_4816),
.A2(n_473),
.B1(n_474),
.B2(n_476),
.Y(n_4880)
);

AOI221xp5_ASAP7_75t_L g4881 ( 
.A1(n_4830),
.A2(n_476),
.B1(n_477),
.B2(n_478),
.C(n_479),
.Y(n_4881)
);

AOI221x1_ASAP7_75t_L g4882 ( 
.A1(n_4847),
.A2(n_477),
.B1(n_479),
.B2(n_480),
.C(n_481),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4836),
.Y(n_4883)
);

AOI22xp5_ASAP7_75t_L g4884 ( 
.A1(n_4853),
.A2(n_4864),
.B1(n_4834),
.B2(n_4856),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_L g4885 ( 
.A(n_4863),
.B(n_480),
.Y(n_4885)
);

NOR3x1_ASAP7_75t_L g4886 ( 
.A(n_4840),
.B(n_481),
.C(n_482),
.Y(n_4886)
);

AO22x2_ASAP7_75t_L g4887 ( 
.A1(n_4851),
.A2(n_482),
.B1(n_483),
.B2(n_485),
.Y(n_4887)
);

OAI22xp5_ASAP7_75t_SL g4888 ( 
.A1(n_4818),
.A2(n_483),
.B1(n_486),
.B2(n_487),
.Y(n_4888)
);

OAI22xp33_ASAP7_75t_L g4889 ( 
.A1(n_4857),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.Y(n_4889)
);

OAI221xp5_ASAP7_75t_SL g4890 ( 
.A1(n_4850),
.A2(n_489),
.B1(n_490),
.B2(n_491),
.C(n_492),
.Y(n_4890)
);

NAND3xp33_ASAP7_75t_SL g4891 ( 
.A(n_4818),
.B(n_489),
.C(n_491),
.Y(n_4891)
);

OAI21xp33_ASAP7_75t_SL g4892 ( 
.A1(n_4861),
.A2(n_492),
.B(n_493),
.Y(n_4892)
);

NAND3xp33_ASAP7_75t_SL g4893 ( 
.A(n_4827),
.B(n_493),
.C(n_494),
.Y(n_4893)
);

NOR2xp33_ASAP7_75t_L g4894 ( 
.A(n_4842),
.B(n_494),
.Y(n_4894)
);

AOI221x1_ASAP7_75t_L g4895 ( 
.A1(n_4854),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.C(n_499),
.Y(n_4895)
);

NOR2xp33_ASAP7_75t_L g4896 ( 
.A(n_4843),
.B(n_499),
.Y(n_4896)
);

AOI221xp5_ASAP7_75t_L g4897 ( 
.A1(n_4828),
.A2(n_501),
.B1(n_504),
.B2(n_505),
.C(n_506),
.Y(n_4897)
);

OA21x2_ASAP7_75t_L g4898 ( 
.A1(n_4858),
.A2(n_505),
.B(n_507),
.Y(n_4898)
);

AOI221xp5_ASAP7_75t_L g4899 ( 
.A1(n_4862),
.A2(n_507),
.B1(n_508),
.B2(n_509),
.C(n_510),
.Y(n_4899)
);

OAI211xp5_ASAP7_75t_L g4900 ( 
.A1(n_4849),
.A2(n_509),
.B(n_511),
.C(n_512),
.Y(n_4900)
);

OAI221xp5_ASAP7_75t_L g4901 ( 
.A1(n_4855),
.A2(n_513),
.B1(n_514),
.B2(n_515),
.C(n_516),
.Y(n_4901)
);

NOR3xp33_ASAP7_75t_L g4902 ( 
.A(n_4865),
.B(n_514),
.C(n_516),
.Y(n_4902)
);

AOI21xp5_ASAP7_75t_L g4903 ( 
.A1(n_4859),
.A2(n_517),
.B(n_518),
.Y(n_4903)
);

AOI221xp5_ASAP7_75t_L g4904 ( 
.A1(n_4832),
.A2(n_517),
.B1(n_519),
.B2(n_521),
.C(n_522),
.Y(n_4904)
);

NAND4xp25_ASAP7_75t_SL g4905 ( 
.A(n_4852),
.B(n_519),
.C(n_521),
.D(n_522),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4848),
.Y(n_4906)
);

OAI22xp5_ASAP7_75t_L g4907 ( 
.A1(n_4884),
.A2(n_4845),
.B1(n_4866),
.B2(n_4848),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4898),
.Y(n_4908)
);

AOI22xp5_ASAP7_75t_L g4909 ( 
.A1(n_4873),
.A2(n_4833),
.B1(n_4841),
.B2(n_526),
.Y(n_4909)
);

OAI22xp5_ASAP7_75t_L g4910 ( 
.A1(n_4869),
.A2(n_523),
.B1(n_524),
.B2(n_526),
.Y(n_4910)
);

OAI22xp5_ASAP7_75t_L g4911 ( 
.A1(n_4870),
.A2(n_528),
.B1(n_531),
.B2(n_532),
.Y(n_4911)
);

AOI22xp5_ASAP7_75t_L g4912 ( 
.A1(n_4871),
.A2(n_531),
.B1(n_533),
.B2(n_534),
.Y(n_4912)
);

AOI221xp5_ASAP7_75t_L g4913 ( 
.A1(n_4867),
.A2(n_533),
.B1(n_535),
.B2(n_536),
.C(n_537),
.Y(n_4913)
);

INVxp67_ASAP7_75t_SL g4914 ( 
.A(n_4883),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4898),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4888),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4887),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4887),
.Y(n_4918)
);

AOI221xp5_ASAP7_75t_L g4919 ( 
.A1(n_4877),
.A2(n_536),
.B1(n_537),
.B2(n_538),
.C(n_540),
.Y(n_4919)
);

INVx2_ASAP7_75t_L g4920 ( 
.A(n_4906),
.Y(n_4920)
);

HB1xp67_ASAP7_75t_L g4921 ( 
.A(n_4892),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_4885),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4872),
.Y(n_4923)
);

OAI31xp33_ASAP7_75t_L g4924 ( 
.A1(n_4900),
.A2(n_4889),
.A3(n_4905),
.B(n_4890),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4886),
.Y(n_4925)
);

OAI22xp5_ASAP7_75t_L g4926 ( 
.A1(n_4880),
.A2(n_538),
.B1(n_540),
.B2(n_541),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4894),
.Y(n_4927)
);

INVx1_ASAP7_75t_L g4928 ( 
.A(n_4891),
.Y(n_4928)
);

O2A1O1Ixp5_ASAP7_75t_SL g4929 ( 
.A1(n_4868),
.A2(n_4893),
.B(n_4875),
.C(n_4882),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4896),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4895),
.Y(n_4931)
);

AOI221xp5_ASAP7_75t_L g4932 ( 
.A1(n_4910),
.A2(n_4881),
.B1(n_4897),
.B2(n_4879),
.C(n_4903),
.Y(n_4932)
);

O2A1O1Ixp33_ASAP7_75t_L g4933 ( 
.A1(n_4921),
.A2(n_4902),
.B(n_4901),
.C(n_4876),
.Y(n_4933)
);

NAND4xp25_ASAP7_75t_L g4934 ( 
.A(n_4924),
.B(n_4899),
.C(n_4874),
.D(n_4904),
.Y(n_4934)
);

AND4x1_ASAP7_75t_L g4935 ( 
.A(n_4913),
.B(n_4878),
.C(n_543),
.D(n_544),
.Y(n_4935)
);

AOI211xp5_ASAP7_75t_L g4936 ( 
.A1(n_4907),
.A2(n_542),
.B(n_543),
.C(n_544),
.Y(n_4936)
);

AOI211xp5_ASAP7_75t_L g4937 ( 
.A1(n_4917),
.A2(n_542),
.B(n_545),
.C(n_546),
.Y(n_4937)
);

OAI21xp33_ASAP7_75t_L g4938 ( 
.A1(n_4923),
.A2(n_545),
.B(n_546),
.Y(n_4938)
);

AOI221xp5_ASAP7_75t_L g4939 ( 
.A1(n_4914),
.A2(n_548),
.B1(n_549),
.B2(n_550),
.C(n_551),
.Y(n_4939)
);

NOR2x1_ASAP7_75t_L g4940 ( 
.A(n_4908),
.B(n_4915),
.Y(n_4940)
);

AOI221xp5_ASAP7_75t_L g4941 ( 
.A1(n_4918),
.A2(n_548),
.B1(n_551),
.B2(n_552),
.C(n_553),
.Y(n_4941)
);

NOR4xp75_ASAP7_75t_L g4942 ( 
.A(n_4926),
.B(n_554),
.C(n_555),
.D(n_556),
.Y(n_4942)
);

AOI221xp5_ASAP7_75t_L g4943 ( 
.A1(n_4931),
.A2(n_554),
.B1(n_555),
.B2(n_557),
.C(n_558),
.Y(n_4943)
);

NAND3xp33_ASAP7_75t_SL g4944 ( 
.A(n_4909),
.B(n_557),
.C(n_559),
.Y(n_4944)
);

AOI222xp33_ASAP7_75t_L g4945 ( 
.A1(n_4928),
.A2(n_559),
.B1(n_560),
.B2(n_561),
.C1(n_562),
.C2(n_564),
.Y(n_4945)
);

AOI21xp5_ASAP7_75t_L g4946 ( 
.A1(n_4920),
.A2(n_560),
.B(n_565),
.Y(n_4946)
);

NAND2xp5_ASAP7_75t_L g4947 ( 
.A(n_4925),
.B(n_565),
.Y(n_4947)
);

AOI21xp5_ASAP7_75t_L g4948 ( 
.A1(n_4924),
.A2(n_566),
.B(n_567),
.Y(n_4948)
);

AOI321xp33_ASAP7_75t_SL g4949 ( 
.A1(n_4944),
.A2(n_4929),
.A3(n_4916),
.B1(n_4927),
.B2(n_4930),
.C(n_4922),
.Y(n_4949)
);

AOI22xp5_ASAP7_75t_L g4950 ( 
.A1(n_4934),
.A2(n_4919),
.B1(n_4912),
.B2(n_4911),
.Y(n_4950)
);

NOR2x1_ASAP7_75t_L g4951 ( 
.A(n_4940),
.B(n_566),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_SL g4952 ( 
.A(n_4937),
.B(n_1652),
.Y(n_4952)
);

OAI211xp5_ASAP7_75t_L g4953 ( 
.A1(n_4948),
.A2(n_586),
.B(n_589),
.C(n_592),
.Y(n_4953)
);

OAI321xp33_ASAP7_75t_L g4954 ( 
.A1(n_4932),
.A2(n_594),
.A3(n_595),
.B1(n_598),
.B2(n_599),
.C(n_600),
.Y(n_4954)
);

OAI211xp5_ASAP7_75t_SL g4955 ( 
.A1(n_4933),
.A2(n_603),
.B(n_604),
.C(n_606),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4947),
.Y(n_4956)
);

INVx5_ASAP7_75t_L g4957 ( 
.A(n_4938),
.Y(n_4957)
);

NAND3x1_ASAP7_75t_SL g4958 ( 
.A(n_4943),
.B(n_610),
.C(n_613),
.Y(n_4958)
);

AOI21xp33_ASAP7_75t_L g4959 ( 
.A1(n_4936),
.A2(n_615),
.B(n_617),
.Y(n_4959)
);

OAI211xp5_ASAP7_75t_SL g4960 ( 
.A1(n_4941),
.A2(n_618),
.B(n_620),
.C(n_622),
.Y(n_4960)
);

AOI22xp5_ASAP7_75t_L g4961 ( 
.A1(n_4950),
.A2(n_4945),
.B1(n_4939),
.B2(n_4946),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4951),
.Y(n_4962)
);

NOR2x1_ASAP7_75t_L g4963 ( 
.A(n_4953),
.B(n_4942),
.Y(n_4963)
);

AOI22xp5_ASAP7_75t_L g4964 ( 
.A1(n_4955),
.A2(n_4935),
.B1(n_1592),
.B2(n_1596),
.Y(n_4964)
);

OR2x2_ASAP7_75t_L g4965 ( 
.A(n_4956),
.B(n_625),
.Y(n_4965)
);

AOI21xp5_ASAP7_75t_L g4966 ( 
.A1(n_4959),
.A2(n_628),
.B(n_1592),
.Y(n_4966)
);

AOI211xp5_ASAP7_75t_L g4967 ( 
.A1(n_4960),
.A2(n_1596),
.B(n_1648),
.C(n_1621),
.Y(n_4967)
);

OR5x1_ASAP7_75t_L g4968 ( 
.A(n_4961),
.B(n_4949),
.C(n_4957),
.D(n_4963),
.E(n_4958),
.Y(n_4968)
);

AOI311xp33_ASAP7_75t_L g4969 ( 
.A1(n_4962),
.A2(n_4957),
.A3(n_4952),
.B(n_4954),
.C(n_1569),
.Y(n_4969)
);

NAND3xp33_ASAP7_75t_L g4970 ( 
.A(n_4964),
.B(n_4966),
.C(n_4965),
.Y(n_4970)
);

AND2x2_ASAP7_75t_L g4971 ( 
.A(n_4967),
.B(n_1329),
.Y(n_4971)
);

OAI321xp33_ASAP7_75t_L g4972 ( 
.A1(n_4961),
.A2(n_1596),
.A3(n_1648),
.B1(n_1621),
.B2(n_1569),
.C(n_1589),
.Y(n_4972)
);

NAND4xp75_ASAP7_75t_L g4973 ( 
.A(n_4962),
.B(n_1592),
.C(n_1648),
.D(n_1598),
.Y(n_4973)
);

INVx2_ASAP7_75t_L g4974 ( 
.A(n_4968),
.Y(n_4974)
);

OR3x2_ASAP7_75t_L g4975 ( 
.A(n_4969),
.B(n_1592),
.C(n_1648),
.Y(n_4975)
);

NOR2x1_ASAP7_75t_L g4976 ( 
.A(n_4973),
.B(n_4970),
.Y(n_4976)
);

INVx2_ASAP7_75t_L g4977 ( 
.A(n_4975),
.Y(n_4977)
);

INVx1_ASAP7_75t_L g4978 ( 
.A(n_4974),
.Y(n_4978)
);

OAI22xp5_ASAP7_75t_L g4979 ( 
.A1(n_4978),
.A2(n_4976),
.B1(n_4977),
.B2(n_4971),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4979),
.Y(n_4980)
);

NOR4xp25_ASAP7_75t_L g4981 ( 
.A(n_4980),
.B(n_4972),
.C(n_1592),
.D(n_1596),
.Y(n_4981)
);

AOI22xp33_ASAP7_75t_L g4982 ( 
.A1(n_4981),
.A2(n_1589),
.B1(n_1608),
.B2(n_1569),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_4982),
.Y(n_4983)
);

AOI22xp33_ASAP7_75t_L g4984 ( 
.A1(n_4983),
.A2(n_1589),
.B1(n_1608),
.B2(n_1569),
.Y(n_4984)
);

OA21x2_ASAP7_75t_L g4985 ( 
.A1(n_4984),
.A2(n_1596),
.B(n_1608),
.Y(n_4985)
);

BUFx3_ASAP7_75t_L g4986 ( 
.A(n_4985),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4986),
.B(n_1329),
.Y(n_4987)
);

AOI221xp5_ASAP7_75t_L g4988 ( 
.A1(n_4987),
.A2(n_1589),
.B1(n_1598),
.B2(n_1608),
.C(n_1329),
.Y(n_4988)
);

AOI211xp5_ASAP7_75t_L g4989 ( 
.A1(n_4988),
.A2(n_1589),
.B(n_1598),
.C(n_1682),
.Y(n_4989)
);


endmodule