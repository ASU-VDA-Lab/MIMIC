module fake_netlist_6_2439_n_1694 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1694);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1694;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g149 ( 
.A(n_10),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_60),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_25),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_47),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_34),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_66),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_72),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_43),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_108),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_20),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_32),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_27),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_77),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_135),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_10),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_32),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_16),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_8),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_0),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_37),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_26),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_2),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_91),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_85),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_24),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_69),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_74),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_4),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_133),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_129),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_84),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_40),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_68),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_7),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_79),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_1),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_40),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_47),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_146),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_30),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_33),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_35),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_65),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_51),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_101),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_62),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_42),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_114),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_78),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_33),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_111),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_128),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_106),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_38),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_38),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_142),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_124),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_63),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_97),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_81),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_16),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_102),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_98),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_25),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_18),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_9),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_21),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_76),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_96),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_56),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_100),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_35),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_12),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_140),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_132),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_4),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_82),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_127),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_88),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_3),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_141),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_53),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_73),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_46),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_58),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_123),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_70),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_67),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_42),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_44),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_24),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_27),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_23),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_13),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_87),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_75),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_21),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_90),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_0),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_93),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_7),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_59),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_22),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_83),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_57),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_36),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_94),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_39),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_136),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_20),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_9),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_145),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_46),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_23),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_137),
.Y(n_277)
);

BUFx2_ASAP7_75t_SL g278 ( 
.A(n_17),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_107),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_2),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_3),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_89),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_138),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_14),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_19),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_61),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_1),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_44),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_29),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_99),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_18),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_36),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_120),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_103),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_37),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_29),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_134),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_234),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_234),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_234),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_191),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_234),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_234),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_234),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_200),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_234),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_161),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_234),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_214),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_160),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_263),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_263),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_179),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_179),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_211),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_211),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_223),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_205),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_187),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_225),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_223),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_151),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_171),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_246),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_206),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_207),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_209),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_290),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_229),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_248),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_149),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_158),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_168),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_212),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_185),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_213),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_218),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_188),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_197),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_151),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_244),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_153),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_199),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_244),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_162),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_244),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_237),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_208),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_244),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_252),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_163),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_224),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_253),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_255),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_244),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_256),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_237),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_259),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_275),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_229),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_289),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_235),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_231),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_165),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_236),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_240),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_229),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_235),
.Y(n_372)
);

BUFx8_ASAP7_75t_L g373 ( 
.A(n_343),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_323),
.B(n_157),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_150),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_345),
.B(n_150),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_308),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_299),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_324),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_345),
.B(n_154),
.Y(n_380)
);

OAI21x1_ASAP7_75t_L g381 ( 
.A1(n_344),
.A2(n_190),
.B(n_176),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_324),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_324),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_320),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_325),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_339),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_300),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_300),
.Y(n_390)
);

XNOR2x2_ASAP7_75t_R g391 ( 
.A(n_363),
.B(n_5),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_301),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_301),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_310),
.B(n_159),
.Y(n_396)
);

AND2x6_ASAP7_75t_L g397 ( 
.A(n_344),
.B(n_171),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_303),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_302),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_303),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_304),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_311),
.A2(n_297),
.B1(n_296),
.B2(n_173),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_304),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_348),
.Y(n_404)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_348),
.Y(n_405)
);

INVx6_ASAP7_75t_L g406 ( 
.A(n_348),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_305),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_305),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_354),
.B(n_154),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_307),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_307),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_309),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_354),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_309),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_306),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_354),
.B(n_156),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_367),
.B(n_230),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_350),
.A2(n_198),
.B1(n_287),
.B2(n_181),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_319),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_326),
.B(n_232),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_331),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_333),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_321),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_334),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_368),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_327),
.B(n_286),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_350),
.B(n_237),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_368),
.B(n_176),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_334),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_347),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_335),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_335),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_337),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_368),
.B(n_156),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_349),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_314),
.B(n_167),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_371),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_328),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_343),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_430),
.B(n_314),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_378),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_374),
.B(n_360),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_378),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_388),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_416),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_404),
.Y(n_448)
);

NAND2x1p5_ASAP7_75t_L g449 ( 
.A(n_381),
.B(n_166),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_SL g451 ( 
.A(n_429),
.B(n_340),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_336),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_416),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_416),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_430),
.A2(n_418),
.B1(n_396),
.B2(n_389),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_432),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_432),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_432),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_427),
.B(n_338),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_404),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_437),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_437),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_382),
.Y(n_464)
);

INVx8_ASAP7_75t_L g465 ( 
.A(n_397),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_402),
.B(n_332),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_389),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_390),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_398),
.Y(n_469)
);

INVxp33_ASAP7_75t_SL g470 ( 
.A(n_399),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_427),
.B(n_355),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_405),
.B(n_369),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_390),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_L g476 ( 
.A(n_375),
.B(n_370),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

INVx8_ASAP7_75t_L g478 ( 
.A(n_397),
.Y(n_478)
);

BUFx10_ASAP7_75t_L g479 ( 
.A(n_421),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_393),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_374),
.B(n_360),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_396),
.B(n_167),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_403),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_388),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_403),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_393),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_418),
.B(n_421),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_428),
.B(n_169),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_403),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_405),
.B(n_404),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_428),
.B(n_315),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_400),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_410),
.Y(n_494)
);

NOR2x1p5_ASAP7_75t_L g495 ( 
.A(n_415),
.B(n_152),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_440),
.B(n_315),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_405),
.B(n_241),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_384),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_420),
.B(n_375),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_410),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_400),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_430),
.B(n_316),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_376),
.B(n_316),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_410),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_381),
.A2(n_352),
.B(n_349),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_441),
.B(n_317),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_401),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_376),
.B(n_169),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_401),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_407),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_407),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_413),
.Y(n_512)
);

BUFx6f_ASAP7_75t_SL g513 ( 
.A(n_413),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_408),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_381),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_408),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_411),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_413),
.B(n_243),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_397),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_411),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_412),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_412),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_414),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_406),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_380),
.B(n_170),
.Y(n_525)
);

NAND3xp33_ASAP7_75t_L g526 ( 
.A(n_414),
.B(n_194),
.C(n_190),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_422),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_397),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_438),
.B(n_317),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_379),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_380),
.B(n_170),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_379),
.Y(n_532)
);

BUFx6f_ASAP7_75t_SL g533 ( 
.A(n_391),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_441),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_422),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_406),
.B(n_245),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_406),
.B(n_247),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_424),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_424),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_387),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_406),
.B(n_250),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_409),
.B(n_220),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_406),
.B(n_258),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_379),
.Y(n_544)
);

AOI22x1_ASAP7_75t_L g545 ( 
.A1(n_426),
.A2(n_318),
.B1(n_330),
.B2(n_329),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_383),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_383),
.Y(n_547)
);

OA22x2_ASAP7_75t_L g548 ( 
.A1(n_438),
.A2(n_372),
.B1(n_366),
.B2(n_318),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_426),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_409),
.B(n_220),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_417),
.B(n_322),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_431),
.Y(n_552)
);

BUFx6f_ASAP7_75t_SL g553 ( 
.A(n_431),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_384),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_433),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_383),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_387),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_417),
.B(n_222),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_436),
.A2(n_278),
.B1(n_277),
.B2(n_204),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_433),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_436),
.B(n_260),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_434),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_385),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_385),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_423),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_384),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_394),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_385),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_395),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_395),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_423),
.B(n_322),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_439),
.B(n_329),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_434),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_435),
.B(n_330),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_395),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_439),
.B(n_366),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_394),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_L g578 ( 
.A(n_435),
.B(n_204),
.C(n_194),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_373),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_394),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_397),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_394),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_397),
.Y(n_583)
);

BUFx6f_ASAP7_75t_SL g584 ( 
.A(n_373),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_377),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_373),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_397),
.Y(n_587)
);

AND3x2_ASAP7_75t_L g588 ( 
.A(n_373),
.B(n_277),
.C(n_257),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_419),
.B(n_372),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_509),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_503),
.B(n_257),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_527),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_527),
.Y(n_593)
);

BUFx6f_ASAP7_75t_SL g594 ( 
.A(n_579),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_509),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_535),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_510),
.Y(n_597)
);

O2A1O1Ixp33_ASAP7_75t_L g598 ( 
.A1(n_488),
.A2(n_337),
.B(n_341),
.C(n_365),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_510),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_535),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_455),
.B(n_519),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_538),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_506),
.B(n_419),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_519),
.B(n_171),
.Y(n_604)
);

AND2x6_ASAP7_75t_L g605 ( 
.A(n_515),
.B(n_171),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_551),
.B(n_177),
.Y(n_606)
);

NAND3xp33_ASAP7_75t_L g607 ( 
.A(n_492),
.B(n_193),
.C(n_189),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_516),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_540),
.B(n_261),
.Y(n_609)
);

A2O1A1Ixp33_ASAP7_75t_L g610 ( 
.A1(n_529),
.A2(n_239),
.B(n_183),
.C(n_184),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_496),
.B(n_222),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_559),
.A2(n_267),
.B1(n_249),
.B2(n_233),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_565),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_565),
.Y(n_614)
);

OAI221xp5_ASAP7_75t_L g615 ( 
.A1(n_589),
.A2(n_402),
.B1(n_210),
.B2(n_291),
.C(n_186),
.Y(n_615)
);

OAI22x1_ASAP7_75t_R g616 ( 
.A1(n_585),
.A2(n_425),
.B1(n_386),
.B2(n_181),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_476),
.A2(n_262),
.B1(n_264),
.B2(n_295),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_529),
.B(n_182),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_442),
.B(n_341),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_519),
.B(n_171),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_516),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_443),
.B(n_192),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_506),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_444),
.B(n_269),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_481),
.B(n_269),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_538),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_519),
.B(n_244),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_540),
.B(n_557),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_517),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_443),
.B(n_196),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_539),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_557),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_517),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_522),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_489),
.B(n_271),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_522),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_534),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_445),
.B(n_215),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_571),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_539),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_581),
.B(n_244),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_534),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_549),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_450),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_448),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_450),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_470),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_581),
.B(n_219),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_485),
.B(n_342),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_499),
.A2(n_295),
.B1(n_294),
.B2(n_282),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_464),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_549),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_464),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_467),
.B(n_221),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_465),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_467),
.B(n_266),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_548),
.A2(n_274),
.B1(n_279),
.B2(n_283),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_581),
.B(n_298),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_R g659 ( 
.A(n_585),
.B(n_271),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_468),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_473),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_552),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_581),
.B(n_479),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_584),
.B(n_282),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_552),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_442),
.B(n_342),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_446),
.Y(n_667)
);

OAI221xp5_ASAP7_75t_L g668 ( 
.A1(n_482),
.A2(n_346),
.B1(n_365),
.B2(n_364),
.C(n_362),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_555),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_451),
.B(n_346),
.C(n_364),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_473),
.B(n_397),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_508),
.A2(n_353),
.B(n_362),
.C(n_361),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_477),
.B(n_397),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_479),
.B(n_294),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_502),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_477),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_555),
.Y(n_677)
);

OR2x2_ASAP7_75t_SL g678 ( 
.A(n_533),
.B(n_351),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_479),
.B(n_352),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_525),
.A2(n_361),
.B1(n_359),
.B2(n_351),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_502),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_560),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_560),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_480),
.B(n_358),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_572),
.B(n_195),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_480),
.B(n_358),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_L g687 ( 
.A(n_472),
.B(n_448),
.Y(n_687)
);

NAND2x1p5_ASAP7_75t_L g688 ( 
.A(n_528),
.B(n_353),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_562),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_479),
.B(n_201),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_548),
.A2(n_152),
.B1(n_155),
.B2(n_164),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_561),
.B(n_202),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_576),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_487),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_562),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_465),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_573),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_548),
.A2(n_155),
.B1(n_164),
.B2(n_172),
.Y(n_698)
);

AND2x6_ASAP7_75t_L g699 ( 
.A(n_515),
.B(n_356),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_484),
.Y(n_700)
);

INVx8_ASAP7_75t_L g701 ( 
.A(n_584),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_515),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_452),
.B(n_203),
.Y(n_703)
);

O2A1O1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_531),
.A2(n_359),
.B(n_357),
.C(n_356),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_487),
.B(n_357),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_460),
.A2(n_254),
.B1(n_216),
.B2(n_217),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_493),
.B(n_226),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_493),
.B(n_227),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_501),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_501),
.B(n_228),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_507),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_511),
.B(n_238),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_511),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_542),
.B(n_242),
.C(n_251),
.Y(n_714)
);

OAI22xp33_ASAP7_75t_L g715 ( 
.A1(n_459),
.A2(n_272),
.B1(n_175),
.B2(n_292),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_514),
.B(n_265),
.Y(n_716)
);

AND2x6_ASAP7_75t_SL g717 ( 
.A(n_533),
.B(n_313),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_514),
.Y(n_718)
);

O2A1O1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_550),
.A2(n_313),
.B(n_312),
.C(n_292),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_L g720 ( 
.A(n_471),
.B(n_273),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_574),
.B(n_261),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_573),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_574),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_466),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_558),
.B(n_174),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_520),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_495),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_520),
.B(n_178),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_521),
.B(n_523),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_521),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_523),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_512),
.B(n_312),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_518),
.B(n_288),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_553),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_587),
.B(n_288),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_447),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_453),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_580),
.Y(n_738)
);

NAND2x1_ASAP7_75t_L g739 ( 
.A(n_524),
.B(n_92),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_513),
.A2(n_284),
.B1(n_281),
.B2(n_280),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_453),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_580),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_454),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_491),
.B(n_284),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_524),
.B(n_484),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_484),
.B(n_281),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_582),
.Y(n_747)
);

AOI22x1_ASAP7_75t_L g748 ( 
.A1(n_449),
.A2(n_280),
.B1(n_276),
.B2(n_273),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_587),
.Y(n_749)
);

BUFx12f_ASAP7_75t_SL g750 ( 
.A(n_584),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_466),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_495),
.B(n_261),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_583),
.B(n_276),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_583),
.B(n_272),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_528),
.B(n_270),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_611),
.B(n_497),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_644),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_642),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_749),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_749),
.Y(n_760)
);

INVx4_ASAP7_75t_L g761 ( 
.A(n_701),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_SL g762 ( 
.A(n_611),
.B(n_578),
.C(n_180),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_639),
.B(n_484),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_601),
.A2(n_449),
.B1(n_513),
.B2(n_579),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_675),
.B(n_586),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_700),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_739),
.Y(n_767)
);

INVx5_ASAP7_75t_L g768 ( 
.A(n_699),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_646),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_700),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_646),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_685),
.B(n_498),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_693),
.B(n_553),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_651),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_632),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_651),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_637),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_685),
.B(n_498),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_653),
.Y(n_779)
);

AND2x6_ASAP7_75t_SL g780 ( 
.A(n_725),
.B(n_533),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_653),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_703),
.B(n_498),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_647),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_601),
.A2(n_606),
.B1(n_645),
.B2(n_591),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_623),
.B(n_449),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_667),
.Y(n_786)
);

BUFx12f_ASAP7_75t_L g787 ( 
.A(n_717),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_660),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_SL g789 ( 
.A(n_615),
.B(n_578),
.C(n_180),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_660),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_703),
.B(n_592),
.Y(n_791)
);

OR2x6_ASAP7_75t_L g792 ( 
.A(n_701),
.B(n_465),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_661),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_661),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_676),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_603),
.B(n_553),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_676),
.Y(n_797)
);

INVx6_ASAP7_75t_L g798 ( 
.A(n_619),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_702),
.A2(n_526),
.B1(n_505),
.B2(n_545),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_694),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_727),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_733),
.A2(n_513),
.B1(n_536),
.B2(n_537),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_729),
.A2(n_567),
.B1(n_554),
.B2(n_498),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_694),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_613),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_709),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_709),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_696),
.Y(n_808)
);

BUFx6f_ASAP7_75t_SL g809 ( 
.A(n_619),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_733),
.A2(n_541),
.B1(n_543),
.B2(n_554),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_711),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_711),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_614),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_604),
.A2(n_478),
.B(n_465),
.Y(n_814)
);

CKINVDCx11_ASAP7_75t_R g815 ( 
.A(n_616),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_593),
.B(n_554),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_713),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_635),
.A2(n_567),
.B1(n_554),
.B2(n_582),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_734),
.B(n_465),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_718),
.B(n_528),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_699),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_718),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_699),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_635),
.A2(n_567),
.B1(n_577),
.B2(n_469),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_596),
.B(n_600),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_730),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_730),
.B(n_731),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_681),
.B(n_567),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_731),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_609),
.B(n_588),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_699),
.Y(n_831)
);

OR2x4_ASAP7_75t_L g832 ( 
.A(n_725),
.B(n_624),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_602),
.B(n_474),
.Y(n_833)
);

AO21x1_ASAP7_75t_L g834 ( 
.A1(n_753),
.A2(n_563),
.B(n_544),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_723),
.B(n_566),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_626),
.B(n_474),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_590),
.Y(n_837)
);

NAND3xp33_ASAP7_75t_L g838 ( 
.A(n_624),
.B(n_545),
.C(n_268),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_595),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_659),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_631),
.B(n_640),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_595),
.B(n_566),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_649),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_643),
.B(n_475),
.Y(n_844)
);

INVx4_ASAP7_75t_L g845 ( 
.A(n_699),
.Y(n_845)
);

AND2x6_ASAP7_75t_L g846 ( 
.A(n_721),
.B(n_494),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_597),
.B(n_566),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_597),
.Y(n_848)
);

BUFx12f_ASAP7_75t_L g849 ( 
.A(n_678),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_599),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_666),
.Y(n_851)
);

INVx5_ASAP7_75t_L g852 ( 
.A(n_605),
.Y(n_852)
);

NOR3xp33_ASAP7_75t_SL g853 ( 
.A(n_715),
.B(n_178),
.C(n_268),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_652),
.B(n_662),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_666),
.Y(n_855)
);

OAI21xp33_ASAP7_75t_L g856 ( 
.A1(n_728),
.A2(n_270),
.B(n_526),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_659),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_665),
.B(n_475),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_674),
.B(n_483),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_608),
.Y(n_860)
);

NOR2x1p5_ASAP7_75t_L g861 ( 
.A(n_752),
.B(n_577),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_608),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_621),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_669),
.B(n_483),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_621),
.B(n_566),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_629),
.B(n_633),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_629),
.B(n_566),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_677),
.B(n_486),
.Y(n_868)
);

AND3x2_ASAP7_75t_SL g869 ( 
.A(n_702),
.B(n_6),
.C(n_8),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_633),
.B(n_634),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_750),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_682),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_679),
.A2(n_504),
.B1(n_500),
.B2(n_490),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_634),
.B(n_478),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_636),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_679),
.A2(n_504),
.B1(n_500),
.B2(n_490),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_636),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_683),
.B(n_486),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_689),
.B(n_494),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_724),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_695),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_697),
.B(n_454),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_722),
.B(n_544),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_726),
.B(n_456),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_663),
.Y(n_885)
);

OR2x2_ASAP7_75t_SL g886 ( 
.A(n_607),
.B(n_6),
.Y(n_886)
);

XOR2x2_ASAP7_75t_L g887 ( 
.A(n_625),
.B(n_11),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_738),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_618),
.A2(n_532),
.B1(n_530),
.B2(n_569),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_744),
.B(n_732),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_728),
.B(n_456),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_746),
.B(n_457),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_670),
.B(n_546),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_691),
.A2(n_457),
.B1(n_458),
.B2(n_461),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_625),
.B(n_478),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_594),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_707),
.Y(n_897)
);

NAND2x1p5_ASAP7_75t_L g898 ( 
.A(n_663),
.B(n_458),
.Y(n_898)
);

CKINVDCx11_ASAP7_75t_R g899 ( 
.A(n_706),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_594),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_736),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_708),
.B(n_710),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_742),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_737),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_747),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_712),
.B(n_462),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_741),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_741),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_743),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_671),
.B(n_478),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_690),
.B(n_462),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_716),
.B(n_463),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_674),
.B(n_564),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_714),
.B(n_705),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_622),
.B(n_463),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_751),
.B(n_563),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_735),
.Y(n_917)
);

NAND2x1p5_ASAP7_75t_L g918 ( 
.A(n_753),
.B(n_754),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_690),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_692),
.B(n_530),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_673),
.B(n_478),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_630),
.B(n_564),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_617),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_684),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_686),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_691),
.A2(n_532),
.B1(n_546),
.B2(n_569),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_692),
.B(n_568),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_881),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_881),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_895),
.A2(n_687),
.B(n_745),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_758),
.B(n_740),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_791),
.B(n_664),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_777),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_916),
.B(n_698),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_821),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_902),
.A2(n_719),
.B(n_754),
.C(n_720),
.Y(n_936)
);

INVx5_ASAP7_75t_L g937 ( 
.A(n_792),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_775),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_759),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_832),
.A2(n_657),
.B1(n_648),
.B2(n_658),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_777),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_813),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_890),
.B(n_897),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_832),
.B(n_650),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_789),
.A2(n_612),
.B(n_610),
.C(n_668),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_814),
.A2(n_658),
.B(n_648),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_757),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_769),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_851),
.B(n_698),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_L g950 ( 
.A1(n_887),
.A2(n_680),
.B(n_657),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_756),
.B(n_825),
.Y(n_951)
);

OR2x6_ASAP7_75t_L g952 ( 
.A(n_761),
.B(n_598),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_821),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_789),
.A2(n_638),
.B(n_654),
.C(n_656),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_814),
.A2(n_620),
.B(n_604),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_805),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_919),
.B(n_748),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_759),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_841),
.B(n_755),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_759),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_854),
.B(n_704),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_813),
.B(n_620),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_796),
.B(n_641),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_771),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_782),
.A2(n_688),
.B(n_627),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_772),
.A2(n_688),
.B(n_547),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_799),
.A2(n_672),
.B1(n_568),
.B2(n_547),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_917),
.A2(n_575),
.B(n_570),
.C(n_556),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_917),
.A2(n_575),
.B(n_570),
.C(n_556),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_778),
.A2(n_784),
.B(n_808),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_776),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_R g972 ( 
.A(n_783),
.B(n_605),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_763),
.B(n_605),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_786),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_843),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_760),
.B(n_575),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_779),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_924),
.B(n_570),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_773),
.B(n_556),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_762),
.A2(n_11),
.B(n_13),
.C(n_14),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_760),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_925),
.B(n_15),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_773),
.B(n_15),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_762),
.A2(n_17),
.B(n_19),
.C(n_22),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_880),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_923),
.B(n_26),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_SL g987 ( 
.A(n_840),
.B(n_28),
.C(n_31),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_760),
.B(n_86),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_781),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_801),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_891),
.B(n_34),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_872),
.B(n_39),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_856),
.A2(n_41),
.B(n_43),
.C(n_45),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_920),
.A2(n_927),
.B(n_859),
.C(n_838),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_764),
.A2(n_41),
.B(n_45),
.C(n_48),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_821),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_798),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_809),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_765),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_812),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_SL g1001 ( 
.A1(n_886),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_920),
.A2(n_49),
.B(n_50),
.C(n_52),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_906),
.A2(n_54),
.B(n_55),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_788),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_855),
.B(n_64),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_799),
.A2(n_71),
.B1(n_95),
.B2(n_104),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_830),
.B(n_105),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_914),
.B(n_109),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_918),
.A2(n_885),
.B1(n_785),
.B2(n_812),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_798),
.B(n_110),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_853),
.A2(n_113),
.B(n_115),
.C(n_116),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_798),
.B(n_119),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_912),
.A2(n_130),
.B(n_139),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_853),
.A2(n_888),
.B(n_903),
.C(n_905),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_790),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_765),
.B(n_861),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_846),
.B(n_828),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_927),
.A2(n_859),
.B(n_913),
.C(n_911),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_821),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_R g1020 ( 
.A(n_857),
.B(n_871),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_794),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_899),
.B(n_809),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_913),
.A2(n_828),
.B(n_802),
.C(n_829),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_774),
.B(n_793),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_800),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_L g1026 ( 
.A(n_815),
.B(n_896),
.C(n_761),
.Y(n_1026)
);

AND2x6_ASAP7_75t_L g1027 ( 
.A(n_885),
.B(n_823),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_SL g1028 ( 
.A1(n_810),
.A2(n_817),
.B(n_766),
.C(n_770),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_918),
.B(n_766),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_874),
.A2(n_892),
.B(n_921),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_R g1031 ( 
.A(n_900),
.B(n_780),
.Y(n_1031)
);

NAND3xp33_ASAP7_75t_L g1032 ( 
.A(n_893),
.B(n_822),
.C(n_807),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_L g1033 ( 
.A(n_896),
.B(n_835),
.C(n_845),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_846),
.B(n_817),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_846),
.B(n_804),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_885),
.A2(n_894),
.B1(n_811),
.B2(n_806),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_826),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_874),
.A2(n_910),
.B(n_921),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_823),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_910),
.A2(n_915),
.B(n_827),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_827),
.A2(n_922),
.B(n_852),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_835),
.A2(n_844),
.B(n_878),
.C(n_868),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_885),
.A2(n_894),
.B1(n_926),
.B2(n_795),
.Y(n_1043)
);

NOR2xp67_ASAP7_75t_SL g1044 ( 
.A(n_852),
.B(n_768),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_852),
.A2(n_898),
.B(n_803),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_833),
.A2(n_858),
.B(n_864),
.C(n_836),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_866),
.A2(n_870),
.B(n_926),
.Y(n_1047)
);

BUFx12f_ASAP7_75t_L g1048 ( 
.A(n_849),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_846),
.B(n_797),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_852),
.A2(n_898),
.B(n_816),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_893),
.B(n_883),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_842),
.A2(n_865),
.B(n_847),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_770),
.B(n_863),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_862),
.B(n_877),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_860),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_867),
.A2(n_866),
.B(n_870),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_SL g1057 ( 
.A1(n_848),
.A2(n_908),
.B(n_875),
.C(n_837),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_862),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_943),
.B(n_850),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_1056),
.A2(n_834),
.B(n_867),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_SL g1061 ( 
.A1(n_1014),
.A2(n_845),
.B(n_879),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_963),
.A2(n_818),
.B(n_824),
.C(n_882),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_951),
.B(n_883),
.Y(n_1063)
);

NAND2x1p5_ASAP7_75t_L g1064 ( 
.A(n_937),
.B(n_768),
.Y(n_1064)
);

OA21x2_ASAP7_75t_L g1065 ( 
.A1(n_994),
.A2(n_884),
.B(n_873),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_1038),
.A2(n_889),
.B(n_876),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1018),
.A2(n_907),
.B(n_909),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_970),
.A2(n_768),
.B(n_767),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1051),
.B(n_934),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1024),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1055),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_937),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_933),
.Y(n_1073)
);

AO21x2_ASAP7_75t_L g1074 ( 
.A1(n_1028),
.A2(n_820),
.B(n_839),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1040),
.A2(n_904),
.B(n_901),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_959),
.B(n_961),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_SL g1077 ( 
.A1(n_1006),
.A2(n_792),
.B(n_831),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_947),
.B(n_877),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_1030),
.A2(n_930),
.B(n_955),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_946),
.A2(n_767),
.B(n_792),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_948),
.Y(n_1081)
);

NOR2xp67_ASAP7_75t_SL g1082 ( 
.A(n_1048),
.B(n_787),
.Y(n_1082)
);

BUFx10_ASAP7_75t_L g1083 ( 
.A(n_1022),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_964),
.B(n_862),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_971),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_977),
.B(n_877),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1023),
.A2(n_819),
.B(n_869),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_937),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_965),
.A2(n_1046),
.B(n_1045),
.Y(n_1089)
);

AO32x2_ASAP7_75t_L g1090 ( 
.A1(n_1043),
.A2(n_869),
.A3(n_823),
.B1(n_831),
.B2(n_767),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_1016),
.B(n_819),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_R g1092 ( 
.A(n_985),
.B(n_831),
.Y(n_1092)
);

NOR2x1_ASAP7_75t_SL g1093 ( 
.A(n_952),
.B(n_819),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_989),
.B(n_767),
.Y(n_1094)
);

INVxp67_ASAP7_75t_SL g1095 ( 
.A(n_942),
.Y(n_1095)
);

AOI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_954),
.A2(n_991),
.B(n_995),
.Y(n_1096)
);

NOR2xp67_ASAP7_75t_L g1097 ( 
.A(n_990),
.B(n_975),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1042),
.A2(n_1043),
.B(n_1050),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1041),
.A2(n_966),
.B(n_936),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1047),
.A2(n_967),
.B(n_940),
.Y(n_1100)
);

AOI21x1_ASAP7_75t_L g1101 ( 
.A1(n_957),
.A2(n_1036),
.B(n_967),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1004),
.Y(n_1102)
);

BUFx4_ASAP7_75t_SL g1103 ( 
.A(n_956),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_938),
.Y(n_1104)
);

NOR2xp67_ASAP7_75t_L g1105 ( 
.A(n_941),
.B(n_997),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_931),
.B(n_974),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1047),
.A2(n_1036),
.B(n_945),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_949),
.B(n_962),
.Y(n_1108)
);

AOI221xp5_ASAP7_75t_SL g1109 ( 
.A1(n_993),
.A2(n_950),
.B1(n_980),
.B2(n_984),
.C(n_1002),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_999),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1009),
.A2(n_1017),
.B(n_973),
.Y(n_1111)
);

BUFx12f_ASAP7_75t_L g1112 ( 
.A(n_949),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_1006),
.A2(n_979),
.A3(n_1029),
.B(n_1035),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_928),
.Y(n_1114)
);

NAND2x1p5_ASAP7_75t_L g1115 ( 
.A(n_1044),
.B(n_958),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_944),
.B(n_986),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1054),
.A2(n_1032),
.B(n_932),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_998),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1032),
.A2(n_978),
.B(n_1057),
.Y(n_1119)
);

AO21x2_ASAP7_75t_L g1120 ( 
.A1(n_1034),
.A2(n_1049),
.B(n_976),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1015),
.B(n_1021),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1025),
.B(n_1037),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1007),
.B(n_929),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_968),
.A2(n_969),
.B(n_1053),
.Y(n_1124)
);

AND3x4_ASAP7_75t_L g1125 ( 
.A(n_1026),
.B(n_1005),
.C(n_1033),
.Y(n_1125)
);

AO31x2_ASAP7_75t_L g1126 ( 
.A1(n_983),
.A2(n_982),
.A3(n_1013),
.B(n_1003),
.Y(n_1126)
);

INVx4_ASAP7_75t_L g1127 ( 
.A(n_958),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_939),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1000),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1001),
.A2(n_1058),
.B1(n_1008),
.B2(n_1005),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1058),
.B(n_939),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1011),
.A2(n_988),
.B(n_1010),
.Y(n_1132)
);

OAI22x1_ASAP7_75t_L g1133 ( 
.A1(n_992),
.A2(n_1012),
.B1(n_981),
.B2(n_960),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_987),
.A2(n_981),
.B(n_960),
.C(n_953),
.Y(n_1134)
);

AOI21x1_ASAP7_75t_L g1135 ( 
.A1(n_952),
.A2(n_1027),
.B(n_953),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_935),
.B(n_1019),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_935),
.B(n_953),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_996),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_972),
.B(n_1020),
.Y(n_1139)
);

BUFx2_ASAP7_75t_R g1140 ( 
.A(n_1031),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1027),
.A2(n_996),
.B(n_1019),
.Y(n_1141)
);

O2A1O1Ixp5_ASAP7_75t_L g1142 ( 
.A1(n_1027),
.A2(n_488),
.B(n_932),
.C(n_957),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1019),
.A2(n_970),
.B(n_696),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1039),
.A2(n_951),
.B1(n_832),
.B2(n_943),
.Y(n_1144)
);

AND2x6_ASAP7_75t_L g1145 ( 
.A(n_935),
.B(n_953),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1056),
.A2(n_1038),
.B(n_1052),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_994),
.A2(n_1018),
.B(n_1040),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_951),
.B(n_943),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_951),
.A2(n_832),
.B1(n_943),
.B2(n_702),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_951),
.B(n_943),
.Y(n_1150)
);

AO31x2_ASAP7_75t_L g1151 ( 
.A1(n_994),
.A2(n_1018),
.A3(n_1023),
.B(n_834),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_956),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_986),
.A2(n_983),
.B1(n_466),
.B2(n_919),
.Y(n_1153)
);

BUFx10_ASAP7_75t_L g1154 ( 
.A(n_1022),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_943),
.B(n_628),
.Y(n_1155)
);

OAI21xp33_ASAP7_75t_L g1156 ( 
.A1(n_950),
.A2(n_685),
.B(n_611),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_935),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_937),
.Y(n_1158)
);

O2A1O1Ixp5_ASAP7_75t_L g1159 ( 
.A1(n_932),
.A2(n_488),
.B(n_957),
.C(n_970),
.Y(n_1159)
);

AOI221x1_ASAP7_75t_L g1160 ( 
.A1(n_970),
.A2(n_1006),
.B1(n_1002),
.B2(n_983),
.C(n_994),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1055),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_970),
.A2(n_696),
.B(n_655),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_970),
.A2(n_696),
.B(n_655),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1016),
.B(n_1051),
.Y(n_1164)
);

OA22x2_ASAP7_75t_L g1165 ( 
.A1(n_950),
.A2(n_1001),
.B1(n_402),
.B2(n_466),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1056),
.A2(n_1038),
.B(n_1052),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1055),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_994),
.A2(n_1018),
.A3(n_1023),
.B(n_834),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_951),
.B(n_943),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_994),
.A2(n_1018),
.A3(n_1023),
.B(n_834),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_951),
.B(n_943),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1056),
.A2(n_1038),
.B(n_1052),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1056),
.A2(n_1038),
.B(n_1052),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_956),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_994),
.A2(n_1023),
.B(n_1018),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_956),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_994),
.A2(n_1018),
.A3(n_1023),
.B(n_834),
.Y(n_1177)
);

NOR4xp25_ASAP7_75t_L g1178 ( 
.A(n_980),
.B(n_984),
.C(n_995),
.D(n_993),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_970),
.A2(n_696),
.B(n_655),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1024),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_956),
.Y(n_1181)
);

OR2x6_ASAP7_75t_L g1182 ( 
.A(n_956),
.B(n_761),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_943),
.B(n_308),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1056),
.A2(n_1038),
.B(n_1052),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_SL g1185 ( 
.A1(n_1018),
.A2(n_808),
.B(n_994),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1056),
.A2(n_1038),
.B(n_1052),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_970),
.A2(n_696),
.B(n_655),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1024),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_933),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_1020),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_943),
.B(n_308),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_950),
.A2(n_320),
.B1(n_321),
.B2(n_308),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_951),
.B(n_943),
.Y(n_1193)
);

BUFx10_ASAP7_75t_L g1194 ( 
.A(n_1022),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1148),
.B(n_1150),
.Y(n_1195)
);

AND2x6_ASAP7_75t_SL g1196 ( 
.A(n_1183),
.B(n_1191),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_1190),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1148),
.A2(n_1171),
.B1(n_1193),
.B2(n_1169),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1179),
.A2(n_1187),
.B(n_1166),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_1160),
.A2(n_1089),
.A3(n_1098),
.B(n_1099),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1146),
.A2(n_1173),
.B(n_1172),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1103),
.Y(n_1202)
);

OAI221xp5_ASAP7_75t_L g1203 ( 
.A1(n_1156),
.A2(n_1192),
.B1(n_1109),
.B2(n_1178),
.C(n_1165),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1076),
.B(n_1149),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1184),
.A2(n_1186),
.B(n_1079),
.Y(n_1205)
);

OA21x2_ASAP7_75t_L g1206 ( 
.A1(n_1100),
.A2(n_1147),
.B(n_1107),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1159),
.A2(n_1142),
.B(n_1117),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1075),
.A2(n_1066),
.B(n_1060),
.Y(n_1208)
);

AO21x2_ASAP7_75t_L g1209 ( 
.A1(n_1096),
.A2(n_1147),
.B(n_1100),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1104),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1081),
.Y(n_1211)
);

AND2x6_ASAP7_75t_L g1212 ( 
.A(n_1072),
.B(n_1088),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1116),
.B(n_1155),
.Y(n_1213)
);

CKINVDCx6p67_ASAP7_75t_R g1214 ( 
.A(n_1110),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_SL g1215 ( 
.A1(n_1096),
.A2(n_1087),
.B(n_1076),
.C(n_1132),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1152),
.Y(n_1216)
);

OR2x6_ASAP7_75t_L g1217 ( 
.A(n_1077),
.B(n_1185),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_1107),
.A2(n_1119),
.B(n_1101),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1067),
.A2(n_1087),
.B(n_1124),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1165),
.A2(n_1153),
.B1(n_1130),
.B2(n_1149),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1130),
.A2(n_1144),
.B(n_1132),
.C(n_1178),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1067),
.A2(n_1111),
.B(n_1109),
.Y(n_1222)
);

BUFx10_ASAP7_75t_L g1223 ( 
.A(n_1164),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1150),
.A2(n_1169),
.B1(n_1193),
.B2(n_1171),
.Y(n_1224)
);

AO21x2_ASAP7_75t_L g1225 ( 
.A1(n_1061),
.A2(n_1062),
.B(n_1135),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_SL g1226 ( 
.A1(n_1108),
.A2(n_1144),
.B1(n_1069),
.B2(n_1123),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1175),
.A2(n_1065),
.B(n_1141),
.Y(n_1227)
);

NOR2xp67_ASAP7_75t_L g1228 ( 
.A(n_1070),
.B(n_1180),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1133),
.A2(n_1093),
.A3(n_1094),
.B(n_1134),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1078),
.A2(n_1084),
.B(n_1086),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1121),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_SL g1232 ( 
.A1(n_1141),
.A2(n_1063),
.B(n_1086),
.Y(n_1232)
);

AO31x2_ASAP7_75t_L g1233 ( 
.A1(n_1078),
.A2(n_1084),
.A3(n_1122),
.B(n_1121),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1074),
.A2(n_1120),
.B(n_1122),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_SL g1235 ( 
.A1(n_1131),
.A2(n_1102),
.B(n_1161),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1140),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1091),
.B(n_1088),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1071),
.Y(n_1238)
);

INVxp67_ASAP7_75t_L g1239 ( 
.A(n_1106),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1125),
.A2(n_1112),
.B1(n_1188),
.B2(n_1085),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1157),
.Y(n_1241)
);

AOI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1065),
.A2(n_1167),
.B(n_1131),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1059),
.A2(n_1139),
.B(n_1095),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1157),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1129),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1073),
.A2(n_1105),
.B(n_1115),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1064),
.A2(n_1115),
.B(n_1158),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1151),
.A2(n_1170),
.B(n_1168),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1181),
.Y(n_1249)
);

AO222x2_ASAP7_75t_L g1250 ( 
.A1(n_1091),
.A2(n_1090),
.B1(n_1082),
.B2(n_1154),
.C1(n_1083),
.C2(n_1194),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1064),
.A2(n_1072),
.B(n_1158),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_R g1252 ( 
.A(n_1174),
.B(n_1176),
.Y(n_1252)
);

NAND2x1p5_ASAP7_75t_L g1253 ( 
.A(n_1127),
.B(n_1114),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1136),
.A2(n_1137),
.B(n_1138),
.Y(n_1254)
);

AO21x2_ASAP7_75t_L g1255 ( 
.A1(n_1074),
.A2(n_1120),
.B(n_1170),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1174),
.A2(n_1176),
.B1(n_1189),
.B2(n_1182),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1128),
.Y(n_1257)
);

CKINVDCx11_ASAP7_75t_R g1258 ( 
.A(n_1083),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1154),
.A2(n_1194),
.B1(n_1118),
.B2(n_1092),
.Y(n_1259)
);

OA21x2_ASAP7_75t_L g1260 ( 
.A1(n_1151),
.A2(n_1177),
.B(n_1170),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1151),
.A2(n_1177),
.B(n_1168),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1090),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1097),
.B(n_1127),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1168),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1090),
.A2(n_1182),
.B1(n_1145),
.B2(n_1126),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1177),
.A2(n_1113),
.B(n_1126),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_SL g1267 ( 
.A1(n_1126),
.A2(n_1113),
.B(n_1145),
.C(n_1182),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1145),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1113),
.A2(n_1080),
.B(n_1162),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1145),
.A2(n_1098),
.B(n_1160),
.Y(n_1270)
);

NAND2x1p5_ASAP7_75t_L g1271 ( 
.A(n_1072),
.B(n_937),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1080),
.A2(n_1163),
.B(n_1162),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1151),
.Y(n_1273)
);

NAND2x1p5_ASAP7_75t_L g1274 ( 
.A(n_1072),
.B(n_937),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1148),
.A2(n_1169),
.B1(n_1171),
.B2(n_1150),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1156),
.A2(n_1165),
.B1(n_887),
.B2(n_1001),
.Y(n_1276)
);

AOI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1068),
.A2(n_1080),
.B(n_1101),
.Y(n_1277)
);

OAI211xp5_ASAP7_75t_L g1278 ( 
.A1(n_1156),
.A2(n_488),
.B(n_615),
.C(n_950),
.Y(n_1278)
);

NAND2x1p5_ASAP7_75t_L g1279 ( 
.A(n_1072),
.B(n_937),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1165),
.A2(n_479),
.B1(n_1116),
.B2(n_373),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1103),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_SL g1282 ( 
.A1(n_1093),
.A2(n_1135),
.B(n_1087),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1157),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_SL g1284 ( 
.A1(n_1096),
.A2(n_1002),
.B(n_1006),
.C(n_1008),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1080),
.A2(n_1163),
.B(n_1162),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1089),
.A2(n_1080),
.B(n_1076),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1080),
.A2(n_1163),
.B(n_1162),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1156),
.A2(n_1100),
.B(n_950),
.C(n_1107),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1148),
.B(n_1150),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1091),
.B(n_1093),
.Y(n_1290)
);

OAI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1165),
.A2(n_832),
.B1(n_615),
.B2(n_1148),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1160),
.A2(n_1089),
.A3(n_1098),
.B(n_1099),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1080),
.A2(n_1143),
.B(n_1162),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1148),
.A2(n_1169),
.B1(n_1171),
.B2(n_1150),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1089),
.A2(n_1080),
.B(n_1076),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1157),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1091),
.B(n_1093),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1121),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1156),
.A2(n_488),
.B(n_481),
.C(n_444),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1121),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1104),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1116),
.B(n_1155),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1080),
.A2(n_1143),
.B(n_1162),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1116),
.B(n_1155),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1104),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1116),
.B(n_1155),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1080),
.A2(n_1163),
.B(n_1162),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1156),
.A2(n_1165),
.B1(n_887),
.B2(n_1001),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1116),
.B(n_1155),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1080),
.A2(n_1163),
.B(n_1162),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1072),
.B(n_937),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1091),
.B(n_1093),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1151),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_SL g1314 ( 
.A1(n_1096),
.A2(n_1002),
.B(n_1006),
.C(n_1008),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1081),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1069),
.B(n_1070),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1080),
.A2(n_1143),
.B(n_1162),
.Y(n_1317)
);

O2A1O1Ixp5_ASAP7_75t_L g1318 ( 
.A1(n_1096),
.A2(n_1100),
.B(n_1132),
.C(n_1147),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1091),
.B(n_1093),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_SL g1320 ( 
.A1(n_1093),
.A2(n_1135),
.B(n_1087),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1288),
.A2(n_1278),
.B(n_1203),
.C(n_1284),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1316),
.B(n_1239),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1195),
.B(n_1289),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1213),
.B(n_1302),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_SL g1325 ( 
.A1(n_1217),
.A2(n_1288),
.B(n_1224),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1198),
.B(n_1275),
.Y(n_1326)
);

INVxp67_ASAP7_75t_L g1327 ( 
.A(n_1238),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1238),
.Y(n_1328)
);

AOI21x1_ASAP7_75t_SL g1329 ( 
.A1(n_1273),
.A2(n_1313),
.B(n_1297),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1217),
.A2(n_1294),
.B(n_1299),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1276),
.A2(n_1308),
.B1(n_1220),
.B2(n_1240),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1231),
.B(n_1298),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1300),
.B(n_1304),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1284),
.A2(n_1314),
.B(n_1291),
.C(n_1221),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1252),
.Y(n_1335)
);

O2A1O1Ixp5_ASAP7_75t_L g1336 ( 
.A1(n_1318),
.A2(n_1207),
.B(n_1286),
.C(n_1295),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1306),
.B(n_1309),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1228),
.B(n_1243),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1233),
.B(n_1204),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1291),
.B(n_1220),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1256),
.Y(n_1341)
);

AOI21x1_ASAP7_75t_SL g1342 ( 
.A1(n_1273),
.A2(n_1313),
.B(n_1319),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_SL g1343 ( 
.A1(n_1217),
.A2(n_1263),
.B(n_1246),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1197),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1276),
.A2(n_1308),
.B1(n_1240),
.B2(n_1259),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1252),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1259),
.A2(n_1280),
.B1(n_1226),
.B2(n_1301),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1204),
.B(n_1211),
.Y(n_1348)
);

O2A1O1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1314),
.A2(n_1215),
.B(n_1232),
.C(n_1235),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1237),
.B(n_1254),
.Y(n_1350)
);

NOR2xp67_ASAP7_75t_L g1351 ( 
.A(n_1263),
.B(n_1281),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1315),
.B(n_1210),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_SL g1353 ( 
.A1(n_1206),
.A2(n_1270),
.B(n_1319),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1206),
.A2(n_1270),
.B(n_1319),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1290),
.B(n_1312),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1265),
.A2(n_1305),
.B1(n_1216),
.B2(n_1249),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1245),
.B(n_1257),
.Y(n_1357)
);

A2O1A1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1269),
.A2(n_1250),
.B(n_1312),
.C(n_1293),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1216),
.A2(n_1249),
.B1(n_1253),
.B2(n_1214),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1253),
.A2(n_1312),
.B1(n_1268),
.B2(n_1274),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1233),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1233),
.B(n_1230),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1271),
.A2(n_1311),
.B1(n_1279),
.B2(n_1202),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1202),
.A2(n_1236),
.B1(n_1197),
.B2(n_1250),
.Y(n_1364)
);

CKINVDCx6p67_ASAP7_75t_R g1365 ( 
.A(n_1258),
.Y(n_1365)
);

AOI21x1_ASAP7_75t_SL g1366 ( 
.A1(n_1209),
.A2(n_1267),
.B(n_1320),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1247),
.B(n_1251),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1233),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1223),
.B(n_1230),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1267),
.A2(n_1282),
.B(n_1264),
.C(n_1225),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1258),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1242),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1225),
.A2(n_1218),
.B(n_1219),
.C(n_1222),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1196),
.B(n_1223),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1229),
.B(n_1248),
.Y(n_1375)
);

AOI211xp5_ASAP7_75t_L g1376 ( 
.A1(n_1236),
.A2(n_1269),
.B(n_1317),
.C(n_1303),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1212),
.B(n_1296),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1229),
.B(n_1260),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1219),
.A2(n_1218),
.B1(n_1244),
.B2(n_1241),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1266),
.A2(n_1296),
.B(n_1244),
.Y(n_1380)
);

AOI21x1_ASAP7_75t_SL g1381 ( 
.A1(n_1277),
.A2(n_1200),
.B(n_1292),
.Y(n_1381)
);

O2A1O1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1234),
.A2(n_1255),
.B(n_1260),
.C(n_1261),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1283),
.B(n_1260),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1283),
.B(n_1261),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1248),
.B(n_1261),
.Y(n_1385)
);

AOI21x1_ASAP7_75t_SL g1386 ( 
.A1(n_1200),
.A2(n_1292),
.B(n_1227),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1248),
.A2(n_1266),
.B1(n_1262),
.B2(n_1200),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1266),
.B(n_1227),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1255),
.B(n_1208),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1201),
.B(n_1205),
.Y(n_1390)
);

AOI221x1_ASAP7_75t_SL g1391 ( 
.A1(n_1272),
.A2(n_1285),
.B1(n_1287),
.B2(n_1307),
.C(n_1310),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1285),
.A2(n_1199),
.B(n_584),
.Y(n_1392)
);

OA22x2_ASAP7_75t_L g1393 ( 
.A1(n_1199),
.A2(n_1001),
.B1(n_1125),
.B2(n_1153),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1213),
.B(n_1302),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1217),
.A2(n_584),
.B(n_963),
.Y(n_1395)
);

BUFx4f_ASAP7_75t_SL g1396 ( 
.A(n_1365),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1334),
.A2(n_1321),
.B(n_1325),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1367),
.Y(n_1398)
);

INVxp67_ASAP7_75t_L g1399 ( 
.A(n_1341),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1385),
.B(n_1388),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1383),
.B(n_1384),
.Y(n_1401)
);

NOR2x1_ASAP7_75t_L g1402 ( 
.A(n_1343),
.B(n_1330),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1367),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1369),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1362),
.Y(n_1405)
);

BUFx4f_ASAP7_75t_SL g1406 ( 
.A(n_1371),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1339),
.B(n_1375),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1326),
.B(n_1327),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1328),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1378),
.B(n_1361),
.Y(n_1410)
);

AOI221xp5_ASAP7_75t_L g1411 ( 
.A1(n_1331),
.A2(n_1334),
.B1(n_1321),
.B2(n_1345),
.C(n_1340),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1389),
.B(n_1353),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1390),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1368),
.B(n_1387),
.Y(n_1414)
);

OR2x6_ASAP7_75t_L g1415 ( 
.A(n_1392),
.B(n_1354),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1327),
.B(n_1323),
.Y(n_1416)
);

OR2x6_ASAP7_75t_L g1417 ( 
.A(n_1370),
.B(n_1358),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1338),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1347),
.B(n_1393),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1372),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1379),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1348),
.Y(n_1422)
);

AO21x2_ASAP7_75t_L g1423 ( 
.A1(n_1373),
.A2(n_1382),
.B(n_1370),
.Y(n_1423)
);

INVxp33_ASAP7_75t_L g1424 ( 
.A(n_1344),
.Y(n_1424)
);

AOI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1374),
.A2(n_1363),
.B(n_1393),
.Y(n_1425)
);

INVxp67_ASAP7_75t_L g1426 ( 
.A(n_1352),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1336),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1336),
.B(n_1373),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1355),
.B(n_1350),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1382),
.Y(n_1430)
);

OR2x6_ASAP7_75t_L g1431 ( 
.A(n_1395),
.B(n_1380),
.Y(n_1431)
);

NAND3xp33_ASAP7_75t_L g1432 ( 
.A(n_1349),
.B(n_1364),
.C(n_1376),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1332),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1349),
.Y(n_1434)
);

AO21x1_ASAP7_75t_SL g1435 ( 
.A1(n_1329),
.A2(n_1342),
.B(n_1366),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1400),
.B(n_1394),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1407),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1400),
.B(n_1357),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1398),
.B(n_1377),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1400),
.B(n_1386),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1407),
.B(n_1322),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1413),
.B(n_1356),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1413),
.B(n_1381),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1401),
.B(n_1324),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1422),
.B(n_1333),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1405),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1435),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1409),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1422),
.B(n_1391),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1401),
.B(n_1337),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1401),
.B(n_1412),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1409),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1409),
.Y(n_1453)
);

CKINVDCx16_ASAP7_75t_R g1454 ( 
.A(n_1417),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1423),
.A2(n_1366),
.B(n_1329),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1407),
.B(n_1335),
.Y(n_1456)
);

OAI31xp33_ASAP7_75t_L g1457 ( 
.A1(n_1449),
.A2(n_1432),
.A3(n_1419),
.B(n_1418),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1448),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1454),
.A2(n_1411),
.B1(n_1419),
.B2(n_1397),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1448),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1439),
.B(n_1403),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_SL g1462 ( 
.A1(n_1454),
.A2(n_1397),
.B1(n_1432),
.B2(n_1417),
.Y(n_1462)
);

OAI21xp33_ASAP7_75t_L g1463 ( 
.A1(n_1449),
.A2(n_1411),
.B(n_1417),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1456),
.B(n_1428),
.C(n_1417),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1454),
.A2(n_1402),
.B1(n_1417),
.B2(n_1418),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1451),
.B(n_1429),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1445),
.A2(n_1426),
.B1(n_1399),
.B2(n_1428),
.C(n_1408),
.Y(n_1467)
);

BUFx10_ASAP7_75t_L g1468 ( 
.A(n_1439),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1456),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1456),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1441),
.Y(n_1471)
);

OA222x2_ASAP7_75t_L g1472 ( 
.A1(n_1437),
.A2(n_1417),
.B1(n_1431),
.B2(n_1415),
.C1(n_1430),
.C2(n_1404),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1447),
.A2(n_1402),
.B(n_1346),
.C(n_1434),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1450),
.B(n_1426),
.Y(n_1474)
);

INVx5_ASAP7_75t_SL g1475 ( 
.A(n_1447),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_R g1476 ( 
.A(n_1447),
.B(n_1396),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1452),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1445),
.A2(n_1399),
.B1(n_1428),
.B2(n_1408),
.C(n_1421),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1441),
.B(n_1437),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1450),
.B(n_1433),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1452),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1441),
.A2(n_1434),
.B1(n_1424),
.B2(n_1430),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1455),
.A2(n_1427),
.B1(n_1396),
.B2(n_1421),
.Y(n_1483)
);

NAND2xp33_ASAP7_75t_R g1484 ( 
.A(n_1442),
.B(n_1431),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_SL g1485 ( 
.A1(n_1442),
.A2(n_1425),
.B(n_1359),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1452),
.Y(n_1486)
);

OAI322xp33_ASAP7_75t_L g1487 ( 
.A1(n_1453),
.A2(n_1416),
.A3(n_1433),
.B1(n_1410),
.B2(n_1405),
.C1(n_1414),
.C2(n_1420),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1439),
.B(n_1403),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1446),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_L g1490 ( 
.A(n_1443),
.B(n_1427),
.C(n_1420),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1447),
.A2(n_1425),
.B1(n_1431),
.B2(n_1351),
.Y(n_1491)
);

OR2x6_ASAP7_75t_L g1492 ( 
.A(n_1447),
.B(n_1431),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1447),
.A2(n_1431),
.B1(n_1416),
.B2(n_1406),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1458),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1492),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1492),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1492),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1468),
.Y(n_1498)
);

INVx4_ASAP7_75t_SL g1499 ( 
.A(n_1476),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1460),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1468),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1470),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_SL g1503 ( 
.A(n_1457),
.B(n_1447),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1470),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1489),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1467),
.B(n_1438),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1477),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1481),
.Y(n_1508)
);

INVxp67_ASAP7_75t_L g1509 ( 
.A(n_1490),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1462),
.A2(n_1455),
.B(n_1423),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1486),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1479),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1489),
.B(n_1446),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1471),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1480),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1474),
.B(n_1427),
.Y(n_1516)
);

NAND3xp33_ASAP7_75t_SL g1517 ( 
.A(n_1463),
.B(n_1459),
.C(n_1482),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1466),
.B(n_1440),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1487),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1469),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1478),
.B(n_1438),
.Y(n_1521)
);

NAND3xp33_ASAP7_75t_SL g1522 ( 
.A(n_1459),
.B(n_1442),
.C(n_1360),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1482),
.B(n_1438),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1461),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1488),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1494),
.Y(n_1526)
);

NAND3xp33_ASAP7_75t_L g1527 ( 
.A(n_1503),
.B(n_1483),
.C(n_1464),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1519),
.B(n_1509),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1495),
.B(n_1472),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1516),
.B(n_1512),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1503),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1494),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1500),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1516),
.B(n_1485),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1513),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1518),
.B(n_1475),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1500),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1513),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1519),
.B(n_1436),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1509),
.B(n_1521),
.Y(n_1540)
);

OAI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1517),
.A2(n_1473),
.B1(n_1465),
.B2(n_1491),
.C(n_1484),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1507),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1518),
.B(n_1475),
.Y(n_1543)
);

CKINVDCx16_ASAP7_75t_R g1544 ( 
.A(n_1517),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1505),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1513),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1518),
.B(n_1475),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1496),
.B(n_1497),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1496),
.B(n_1436),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1496),
.B(n_1436),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1496),
.B(n_1436),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1505),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1507),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1508),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1511),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1497),
.B(n_1440),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1506),
.B(n_1444),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1506),
.B(n_1444),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1520),
.B(n_1406),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1497),
.B(n_1524),
.Y(n_1560)
);

OR2x6_ASAP7_75t_L g1561 ( 
.A(n_1510),
.B(n_1415),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1520),
.B(n_1473),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1497),
.B(n_1524),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1544),
.A2(n_1522),
.B1(n_1510),
.B2(n_1499),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1545),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1544),
.B(n_1528),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1545),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1528),
.B(n_1523),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1536),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1562),
.Y(n_1570)
);

INVxp67_ASAP7_75t_SL g1571 ( 
.A(n_1562),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1552),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1555),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1552),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1539),
.B(n_1512),
.Y(n_1575)
);

NOR3xp33_ASAP7_75t_L g1576 ( 
.A(n_1540),
.B(n_1522),
.C(n_1493),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1526),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1539),
.B(n_1523),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1540),
.B(n_1514),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1536),
.B(n_1525),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1526),
.Y(n_1581)
);

INVxp67_ASAP7_75t_SL g1582 ( 
.A(n_1531),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1543),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1530),
.B(n_1515),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1530),
.B(n_1515),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1532),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1532),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1543),
.B(n_1525),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1548),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1533),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1533),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1548),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1537),
.Y(n_1593)
);

NOR2xp67_ASAP7_75t_L g1594 ( 
.A(n_1531),
.B(n_1498),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1537),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1547),
.B(n_1525),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1547),
.B(n_1525),
.Y(n_1597)
);

OAI21xp5_ASAP7_75t_SL g1598 ( 
.A1(n_1527),
.A2(n_1465),
.B(n_1493),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1594),
.B(n_1499),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1573),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1574),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1571),
.B(n_1549),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1583),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1582),
.B(n_1583),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1592),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1574),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_1583),
.Y(n_1607)
);

NAND2xp33_ASAP7_75t_L g1608 ( 
.A(n_1576),
.B(n_1564),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1570),
.B(n_1559),
.Y(n_1609)
);

NAND2x1_ASAP7_75t_L g1610 ( 
.A(n_1569),
.B(n_1529),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1589),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1566),
.B(n_1549),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1569),
.B(n_1560),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1565),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1567),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1572),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1580),
.B(n_1560),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1575),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1575),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1579),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1577),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1578),
.B(n_1534),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1573),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1604),
.B(n_1568),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1604),
.Y(n_1625)
);

O2A1O1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1608),
.A2(n_1598),
.B(n_1541),
.C(n_1527),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1609),
.A2(n_1541),
.B1(n_1605),
.B2(n_1617),
.Y(n_1627)
);

O2A1O1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1610),
.A2(n_1561),
.B(n_1529),
.C(n_1578),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1613),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1617),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1611),
.Y(n_1631)
);

AOI21xp33_ASAP7_75t_L g1632 ( 
.A1(n_1607),
.A2(n_1610),
.B(n_1618),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_SL g1633 ( 
.A1(n_1622),
.A2(n_1561),
.B1(n_1534),
.B2(n_1596),
.C(n_1597),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1611),
.Y(n_1634)
);

INVx1_ASAP7_75t_SL g1635 ( 
.A(n_1613),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1599),
.B(n_1580),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1601),
.Y(n_1637)
);

AOI321xp33_ASAP7_75t_L g1638 ( 
.A1(n_1612),
.A2(n_1602),
.A3(n_1622),
.B1(n_1603),
.B2(n_1615),
.C(n_1614),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1601),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1614),
.B(n_1588),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1606),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1603),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1629),
.B(n_1619),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1635),
.B(n_1620),
.Y(n_1644)
);

NOR2x1_ASAP7_75t_L g1645 ( 
.A(n_1631),
.B(n_1599),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1636),
.B(n_1599),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1625),
.B(n_1615),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1631),
.B(n_1616),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1634),
.B(n_1627),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1634),
.B(n_1616),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1630),
.B(n_1606),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1632),
.A2(n_1561),
.B1(n_1599),
.B2(n_1588),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1646),
.B(n_1640),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1651),
.Y(n_1654)
);

AOI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1649),
.A2(n_1626),
.B1(n_1640),
.B2(n_1633),
.C(n_1628),
.Y(n_1655)
);

OAI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1652),
.A2(n_1638),
.B1(n_1624),
.B2(n_1630),
.C(n_1561),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1645),
.A2(n_1636),
.B(n_1642),
.Y(n_1657)
);

NOR2x1_ASAP7_75t_L g1658 ( 
.A(n_1648),
.B(n_1650),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_SL g1659 ( 
.A1(n_1643),
.A2(n_1644),
.B(n_1647),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1649),
.A2(n_1642),
.B(n_1639),
.Y(n_1660)
);

AO21x1_ASAP7_75t_L g1661 ( 
.A1(n_1649),
.A2(n_1641),
.B(n_1637),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_SL g1662 ( 
.A1(n_1655),
.A2(n_1621),
.B(n_1597),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1661),
.A2(n_1656),
.B1(n_1653),
.B2(n_1659),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1658),
.A2(n_1621),
.B(n_1561),
.Y(n_1664)
);

NOR3xp33_ASAP7_75t_L g1665 ( 
.A(n_1654),
.B(n_1623),
.C(n_1600),
.Y(n_1665)
);

AOI221x1_ASAP7_75t_SL g1666 ( 
.A1(n_1660),
.A2(n_1623),
.B1(n_1600),
.B2(n_1581),
.C(n_1586),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1665),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1663),
.B(n_1657),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1662),
.B(n_1596),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1666),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1664),
.Y(n_1671)
);

NOR3xp33_ASAP7_75t_L g1672 ( 
.A(n_1663),
.B(n_1623),
.C(n_1600),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_R g1673 ( 
.A(n_1667),
.B(n_1671),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1668),
.A2(n_1561),
.B1(n_1563),
.B2(n_1499),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1672),
.A2(n_1590),
.B(n_1587),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1669),
.Y(n_1676)
);

NAND4xp25_ASAP7_75t_SL g1677 ( 
.A(n_1672),
.B(n_1595),
.C(n_1593),
.D(n_1591),
.Y(n_1677)
);

NOR3xp33_ASAP7_75t_L g1678 ( 
.A(n_1676),
.B(n_1670),
.C(n_1563),
.Y(n_1678)
);

NOR3xp33_ASAP7_75t_L g1679 ( 
.A(n_1677),
.B(n_1557),
.C(n_1558),
.Y(n_1679)
);

NOR2x1_ASAP7_75t_L g1680 ( 
.A(n_1675),
.B(n_1584),
.Y(n_1680)
);

NOR4xp75_ASAP7_75t_L g1681 ( 
.A(n_1678),
.B(n_1673),
.C(n_1674),
.D(n_1556),
.Y(n_1681)
);

OAI32xp33_ASAP7_75t_L g1682 ( 
.A1(n_1681),
.A2(n_1679),
.A3(n_1680),
.B1(n_1538),
.B2(n_1546),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1585),
.B1(n_1584),
.B2(n_1538),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1682),
.Y(n_1684)
);

OAI21x1_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1585),
.B(n_1535),
.Y(n_1685)
);

AO22x2_ASAP7_75t_L g1686 ( 
.A1(n_1683),
.A2(n_1538),
.B1(n_1535),
.B2(n_1546),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1686),
.A2(n_1535),
.B1(n_1546),
.B2(n_1555),
.Y(n_1687)
);

AOI22x1_ASAP7_75t_L g1688 ( 
.A1(n_1685),
.A2(n_1555),
.B1(n_1542),
.B2(n_1554),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1688),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1689),
.A2(n_1687),
.B1(n_1542),
.B2(n_1553),
.C(n_1554),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1690),
.A2(n_1556),
.B1(n_1553),
.B2(n_1499),
.Y(n_1691)
);

AOI322xp5_ASAP7_75t_L g1692 ( 
.A1(n_1691),
.A2(n_1501),
.A3(n_1502),
.B1(n_1504),
.B2(n_1551),
.C1(n_1550),
.C2(n_1498),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1692),
.A2(n_1499),
.B1(n_1551),
.B2(n_1550),
.Y(n_1693)
);

AOI211xp5_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1476),
.B(n_1558),
.C(n_1557),
.Y(n_1694)
);


endmodule