module fake_aes_12495_n_10 (n_1, n_2, n_0, n_10);
input n_1;
input n_2;
input n_0;
output n_10;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
BUFx6f_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
INVx1_ASAP7_75t_SL g6 ( .A(n_5), .Y(n_6) );
INVx1_ASAP7_75t_SL g7 ( .A(n_6), .Y(n_7) );
AO22x2_ASAP7_75t_L g8 ( .A1(n_7), .A2(n_1), .B1(n_2), .B2(n_5), .Y(n_8) );
INVxp67_ASAP7_75t_SL g9 ( .A(n_8), .Y(n_9) );
OAI222xp33_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_4), .B1(n_8), .B2(n_3), .C1(n_7), .C2(n_6), .Y(n_10) );
endmodule