module fake_jpeg_23351_n_228 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_27),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_38),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_25),
.B1(n_26),
.B2(n_14),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_24),
.B(n_22),
.C(n_17),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_19),
.B1(n_23),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_48),
.B1(n_37),
.B2(n_21),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_14),
.B1(n_26),
.B2(n_15),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_28),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_15),
.B1(n_24),
.B2(n_17),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_20),
.B1(n_34),
.B2(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_25),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_22),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_56),
.B(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_60),
.Y(n_80)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_66),
.B1(n_67),
.B2(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_54),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_37),
.B1(n_42),
.B2(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_37),
.B1(n_32),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_21),
.B1(n_50),
.B2(n_19),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_35),
.B1(n_32),
.B2(n_29),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_32),
.C(n_29),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_30),
.C(n_28),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_77),
.B(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_48),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_79),
.B(n_87),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_52),
.B1(n_39),
.B2(n_55),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_88),
.B1(n_70),
.B2(n_66),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_53),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_89),
.C(n_92),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_49),
.B(n_39),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_44),
.B1(n_19),
.B2(n_23),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_93),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_27),
.B(n_23),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_58),
.B(n_10),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_9),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_67),
.B(n_66),
.C(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_98),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_106),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_46),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_71),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_103),
.B(n_85),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_59),
.B1(n_69),
.B2(n_63),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_109),
.B1(n_87),
.B2(n_78),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_40),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_110),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_60),
.B1(n_30),
.B2(n_27),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_78),
.B1(n_75),
.B2(n_23),
.Y(n_128)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_30),
.C(n_46),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_86),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_96),
.B(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_81),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_117),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g119 ( 
.A(n_104),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_111),
.B1(n_108),
.B2(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_103),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_130),
.Y(n_143)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_116),
.Y(n_157)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_130),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_115),
.B(n_116),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_133),
.A2(n_112),
.B1(n_99),
.B2(n_109),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_123),
.B1(n_43),
.B2(n_62),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_142),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_124),
.B1(n_100),
.B2(n_127),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_146),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_126),
.A2(n_99),
.B1(n_103),
.B2(n_101),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_152),
.B1(n_125),
.B2(n_121),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_9),
.Y(n_148)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_9),
.Y(n_150)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_106),
.B1(n_46),
.B2(n_43),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_168),
.B1(n_136),
.B2(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_161),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_167),
.B(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_120),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_165),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_0),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_179),
.B1(n_161),
.B2(n_164),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_137),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_180),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_139),
.B(n_143),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_173),
.A2(n_177),
.B(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_175),
.B(n_153),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_167),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_135),
.B1(n_147),
.B2(n_152),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_150),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_148),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_182),
.C(n_155),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_138),
.C(n_62),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_185),
.B(n_188),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_170),
.B(n_180),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_192),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_0),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_191),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_153),
.C(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_194),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_166),
.C(n_164),
.Y(n_194)
);

OAI321xp33_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_188),
.A3(n_174),
.B1(n_163),
.B2(n_154),
.C(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_176),
.B1(n_170),
.B2(n_163),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_196),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_199),
.B(n_8),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_6),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_1),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_203),
.B(n_204),
.Y(n_211)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_202),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_208),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_6),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_196),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_206),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_199),
.C(n_198),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_215),
.A2(n_210),
.B(n_211),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_218),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_10),
.Y(n_218)
);

AOI211xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_222),
.B(n_11),
.C(n_12),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_216),
.B(n_213),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_223),
.A2(n_224),
.B(n_221),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_225),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_13),
.B(n_225),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);


endmodule