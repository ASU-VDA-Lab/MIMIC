module fake_jpeg_3595_n_174 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_56),
.Y(n_64)
);

CKINVDCx6p67_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_69),
.Y(n_80)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.Y(n_74)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_58),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_71),
.A2(n_58),
.B1(n_47),
.B2(n_49),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_44),
.B1(n_51),
.B2(n_53),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_44),
.B1(n_51),
.B2(n_53),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_55),
.C(n_54),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_76),
.C(n_80),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_62),
.B1(n_59),
.B2(n_48),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_69),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_59),
.B1(n_52),
.B2(n_57),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

CKINVDCx12_ASAP7_75t_R g91 ( 
.A(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_97),
.Y(n_114)
);

HAxp5_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_61),
.CON(n_93),
.SN(n_93)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_4),
.B(n_5),
.Y(n_108)
);

INVx2_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_95),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_100),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_61),
.C(n_18),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_21),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_61),
.B1(n_1),
.B2(n_2),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_102),
.B1(n_101),
.B2(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_0),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_116),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_82),
.B(n_5),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_108),
.B(n_8),
.Y(n_129)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_11),
.Y(n_135)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_4),
.B(n_7),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_108),
.B(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_7),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_23),
.C(n_43),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_133),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_125),
.C(n_129),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_12),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_27),
.C(n_41),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_134),
.B(n_135),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_11),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_136),
.B(n_138),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_12),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_25),
.C(n_39),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_28),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_143),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_118),
.B1(n_13),
.B2(n_14),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_146),
.B1(n_139),
.B2(n_128),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_133),
.C(n_123),
.Y(n_155)
);

AOI22x1_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_30),
.B1(n_16),
.B2(n_17),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_122),
.B(n_13),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_19),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_20),
.C(n_31),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_148),
.C(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_159),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_163),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_149),
.C(n_132),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_152),
.B1(n_132),
.B2(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_165),
.A2(n_160),
.B(n_152),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_160),
.B(n_146),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_170),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_166),
.A2(n_156),
.B(n_147),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_168),
.B(n_36),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_33),
.Y(n_174)
);


endmodule