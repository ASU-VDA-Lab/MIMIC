module fake_aes_7657_n_735 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_735);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_735;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g81 ( .A(n_36), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_5), .Y(n_82) );
INVx1_ASAP7_75t_SL g83 ( .A(n_73), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_66), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_65), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_17), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_25), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_41), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_0), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_43), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_75), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_77), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_47), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_71), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_24), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_11), .Y(n_96) );
BUFx10_ASAP7_75t_L g97 ( .A(n_29), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_20), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_14), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_76), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_54), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_80), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_38), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_6), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_40), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_23), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_42), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_16), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_30), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_58), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_74), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_44), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_1), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_7), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_34), .Y(n_115) );
NOR2xp67_ASAP7_75t_L g116 ( .A(n_22), .B(n_67), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_55), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_8), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_6), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_9), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_12), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_48), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_12), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_60), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_11), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_9), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_0), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_35), .Y(n_128) );
NOR2xp67_ASAP7_75t_L g129 ( .A(n_61), .B(n_68), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_56), .Y(n_130) );
BUFx12f_ASAP7_75t_L g131 ( .A(n_97), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_110), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_120), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_110), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_127), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_120), .B(n_1), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_101), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_95), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_95), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_122), .Y(n_141) );
CKINVDCx6p67_ASAP7_75t_R g142 ( .A(n_97), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_101), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_125), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_125), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_122), .B(n_2), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_81), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_85), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_87), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_108), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_91), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_92), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g155 ( .A1(n_127), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_97), .B(n_3), .Y(n_156) );
INVx5_ASAP7_75t_L g157 ( .A(n_116), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_94), .Y(n_158) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_130), .B(n_39), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_100), .Y(n_160) );
AND2x6_ASAP7_75t_L g161 ( .A(n_103), .B(n_37), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_106), .Y(n_162) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_109), .B(n_45), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_111), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_96), .B(n_4), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_124), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_104), .B(n_5), .Y(n_168) );
NOR2x1_ASAP7_75t_L g169 ( .A(n_113), .B(n_7), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_114), .B(n_8), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_119), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_121), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_83), .B(n_49), .Y(n_173) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_126), .B(n_50), .Y(n_174) );
BUFx12f_ASAP7_75t_L g175 ( .A(n_86), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_148), .B(n_86), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_135), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_137), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_137), .A2(n_118), .B1(n_99), .B2(n_84), .Y(n_179) );
BUFx10_ASAP7_75t_L g180 ( .A(n_147), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_135), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_137), .A2(n_90), .B1(n_84), .B2(n_105), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_147), .B(n_129), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_135), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_135), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_132), .Y(n_187) );
NAND2xp33_ASAP7_75t_L g188 ( .A(n_161), .B(n_102), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_136), .B(n_107), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_136), .B(n_98), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_139), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_147), .B(n_105), .Y(n_192) );
INVx4_ASAP7_75t_L g193 ( .A(n_161), .Y(n_193) );
INVx4_ASAP7_75t_L g194 ( .A(n_161), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_132), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_142), .B(n_10), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_159), .A2(n_115), .B1(n_112), .B2(n_90), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_172), .B(n_115), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_148), .B(n_117), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_172), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_134), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_139), .Y(n_203) );
INVx5_ASAP7_75t_L g204 ( .A(n_161), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_139), .Y(n_205) );
INVx4_ASAP7_75t_L g206 ( .A(n_161), .Y(n_206) );
BUFx10_ASAP7_75t_L g207 ( .A(n_159), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_142), .B(n_123), .Y(n_208) );
BUFx2_ASAP7_75t_L g209 ( .A(n_175), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_153), .B(n_93), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_172), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
BUFx4f_ASAP7_75t_L g213 ( .A(n_131), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_159), .B(n_112), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_163), .A2(n_123), .B1(n_89), .B2(n_82), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_175), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_171), .Y(n_218) );
BUFx12f_ASAP7_75t_L g219 ( .A(n_131), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_171), .Y(n_220) );
NOR2x1p5_ASAP7_75t_L g221 ( .A(n_146), .B(n_89), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_153), .B(n_82), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_174), .Y(n_223) );
INVx1_ASAP7_75t_SL g224 ( .A(n_174), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_139), .Y(n_225) );
AOI22xp33_ASAP7_75t_SL g226 ( .A1(n_174), .A2(n_10), .B1(n_13), .B2(n_14), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_149), .B(n_13), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_163), .B(n_52), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_149), .B(n_15), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_139), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_163), .B(n_51), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_140), .Y(n_232) );
OR2x2_ASAP7_75t_L g233 ( .A(n_150), .B(n_15), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_150), .A2(n_79), .B1(n_19), .B2(n_21), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_152), .B(n_18), .Y(n_235) );
INVx4_ASAP7_75t_L g236 ( .A(n_161), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_140), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_152), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_158), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_158), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_240) );
AND2x6_ASAP7_75t_L g241 ( .A(n_162), .B(n_46), .Y(n_241) );
OR2x6_ASAP7_75t_L g242 ( .A(n_156), .B(n_53), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_176), .B(n_162), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_201), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_239), .B(n_164), .Y(n_245) );
NAND2x1p5_ASAP7_75t_L g246 ( .A(n_213), .B(n_169), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_176), .B(n_200), .Y(n_247) );
OAI22x1_ASAP7_75t_L g248 ( .A1(n_221), .A2(n_155), .B1(n_169), .B2(n_166), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_200), .B(n_164), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_201), .B(n_166), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_218), .B(n_170), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_211), .Y(n_252) );
AND2x6_ASAP7_75t_SL g253 ( .A(n_208), .B(n_168), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_212), .B(n_146), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_219), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_194), .B(n_157), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_219), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_220), .B(n_161), .Y(n_258) );
INVxp67_ASAP7_75t_L g259 ( .A(n_222), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_213), .B(n_146), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_228), .A2(n_145), .B1(n_138), .B2(n_143), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_191), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_189), .B(n_133), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_224), .A2(n_145), .B1(n_143), .B2(n_138), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_187), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_191), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_190), .B(n_133), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_210), .B(n_144), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_193), .B(n_154), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_217), .B(n_144), .Y(n_270) );
NAND3xp33_ASAP7_75t_SL g271 ( .A(n_223), .B(n_151), .C(n_173), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_193), .B(n_154), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_184), .B(n_157), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_184), .B(n_157), .Y(n_274) );
O2A1O1Ixp5_ASAP7_75t_L g275 ( .A1(n_228), .A2(n_151), .B(n_173), .C(n_157), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_197), .B(n_157), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_178), .B(n_157), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_231), .A2(n_173), .B1(n_167), .B2(n_160), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_231), .A2(n_173), .B1(n_167), .B2(n_160), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_192), .B(n_173), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_180), .B(n_167), .Y(n_281) );
INVx2_ASAP7_75t_SL g282 ( .A(n_180), .Y(n_282) );
INVx4_ASAP7_75t_L g283 ( .A(n_180), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_195), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_192), .B(n_167), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_209), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_214), .B(n_167), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_196), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_192), .B(n_160), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_207), .A2(n_173), .B1(n_160), .B2(n_154), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_227), .B(n_160), .Y(n_291) );
NOR2x2_ASAP7_75t_L g292 ( .A(n_242), .B(n_173), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_194), .B(n_154), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_205), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_193), .B(n_154), .Y(n_295) );
OAI22xp5_ASAP7_75t_SL g296 ( .A1(n_215), .A2(n_141), .B1(n_140), .B2(n_62), .Y(n_296) );
NAND2x1p5_ASAP7_75t_L g297 ( .A(n_233), .B(n_141), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_229), .B(n_141), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_206), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_199), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_199), .Y(n_301) );
NAND2xp33_ASAP7_75t_L g302 ( .A(n_204), .B(n_141), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_202), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_214), .A2(n_141), .B1(n_140), .B2(n_63), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_206), .B(n_140), .Y(n_305) );
OAI221xp5_ASAP7_75t_L g306 ( .A1(n_179), .A2(n_57), .B1(n_59), .B2(n_64), .C(n_69), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_235), .B(n_78), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_199), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_179), .B(n_70), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_242), .B(n_72), .Y(n_310) );
INVxp33_ASAP7_75t_L g311 ( .A(n_216), .Y(n_311) );
OR2x6_ASAP7_75t_L g312 ( .A(n_242), .B(n_238), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_183), .B(n_215), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_286), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_270), .Y(n_315) );
XNOR2xp5_ASAP7_75t_L g316 ( .A(n_255), .B(n_198), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_300), .A2(n_198), .B1(n_183), .B2(n_226), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_283), .B(n_206), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_297), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_259), .B(n_207), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_259), .B(n_207), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_258), .A2(n_188), .B(n_236), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_285), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_245), .B(n_236), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_283), .B(n_236), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_297), .Y(n_326) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_300), .A2(n_188), .B(n_240), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_251), .B(n_241), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_SL g329 ( .A1(n_306), .A2(n_240), .B(n_234), .C(n_230), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_313), .B(n_241), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_299), .B(n_204), .Y(n_331) );
NOR2xp33_ASAP7_75t_SL g332 ( .A(n_257), .B(n_241), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_244), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_308), .Y(n_334) );
INVx4_ASAP7_75t_L g335 ( .A(n_310), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_299), .B(n_204), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_249), .B(n_241), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_310), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_289), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_243), .B(n_241), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_247), .B(n_204), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_312), .A2(n_234), .B1(n_181), .B2(n_177), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_299), .B(n_182), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_308), .B(n_205), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_301), .B(n_182), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_263), .B(n_177), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_280), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_299), .B(n_182), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_269), .A2(n_181), .B(n_186), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_265), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_312), .A2(n_186), .B1(n_182), .B2(n_185), .Y(n_351) );
OAI22xp5_ASAP7_75t_SL g352 ( .A1(n_312), .A2(n_230), .B1(n_232), .B2(n_237), .Y(n_352) );
A2O1A1Ixp33_ASAP7_75t_L g353 ( .A1(n_287), .A2(n_232), .B(n_237), .C(n_185), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_282), .B(n_185), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_269), .A2(n_185), .B(n_225), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_280), .B(n_203), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_262), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_267), .B(n_203), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_276), .B(n_203), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_266), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_309), .B(n_203), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_296), .A2(n_225), .B1(n_248), .B2(n_276), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_311), .B(n_225), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_284), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_250), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_288), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_253), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_260), .B(n_225), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_275), .A2(n_261), .B(n_287), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_317), .A2(n_254), .B1(n_252), .B2(n_246), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_315), .B(n_303), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_320), .B(n_254), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_320), .B(n_268), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_350), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_361), .A2(n_278), .B(n_279), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_328), .A2(n_307), .B(n_272), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_334), .A2(n_246), .B1(n_261), .B2(n_264), .Y(n_377) );
AO31x2_ASAP7_75t_L g378 ( .A1(n_342), .A2(n_298), .A3(n_291), .B(n_281), .Y(n_378) );
OAI21xp5_ASAP7_75t_L g379 ( .A1(n_340), .A2(n_304), .B(n_279), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_330), .A2(n_273), .B1(n_274), .B2(n_277), .Y(n_380) );
NAND3xp33_ASAP7_75t_SL g381 ( .A(n_314), .B(n_278), .C(n_290), .Y(n_381) );
AOI221x1_ASAP7_75t_L g382 ( .A1(n_327), .A2(n_271), .B1(n_281), .B2(n_292), .C(n_294), .Y(n_382) );
AOI21xp33_ASAP7_75t_L g383 ( .A1(n_321), .A2(n_256), .B(n_272), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_335), .B(n_290), .Y(n_384) );
NOR2xp33_ASAP7_75t_SL g385 ( .A(n_335), .B(n_295), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_361), .A2(n_295), .B(n_305), .Y(n_386) );
OAI21xp5_ASAP7_75t_L g387 ( .A1(n_337), .A2(n_293), .B(n_302), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_338), .B(n_365), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g389 ( .A1(n_324), .A2(n_329), .B(n_351), .C(n_323), .Y(n_389) );
BUFx4f_ASAP7_75t_SL g390 ( .A(n_367), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_322), .A2(n_341), .B(n_343), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_316), .A2(n_364), .B1(n_366), .B2(n_339), .C(n_338), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_363), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_358), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_347), .Y(n_395) );
BUFx12f_ASAP7_75t_L g396 ( .A(n_368), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_333), .B(n_319), .Y(n_397) );
OAI21x1_ASAP7_75t_L g398 ( .A1(n_369), .A2(n_355), .B(n_343), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_329), .A2(n_344), .B(n_356), .C(n_346), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g400 ( .A1(n_353), .A2(n_344), .B(n_331), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_357), .Y(n_401) );
AO32x2_ASAP7_75t_L g402 ( .A1(n_352), .A2(n_362), .A3(n_332), .B1(n_356), .B2(n_359), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_326), .A2(n_359), .B1(n_345), .B2(n_318), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_357), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_370), .A2(n_345), .B1(n_357), .B2(n_360), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_374), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_398), .A2(n_349), .B(n_348), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_392), .A2(n_325), .B1(n_354), .B2(n_357), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_371), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_371), .B(n_360), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_374), .B(n_331), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_373), .B(n_360), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_372), .B(n_360), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_388), .B(n_336), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_393), .B(n_395), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_395), .A2(n_399), .B1(n_380), .B2(n_389), .C(n_377), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_396), .A2(n_381), .B1(n_394), .B2(n_397), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g418 ( .A1(n_394), .A2(n_382), .B1(n_396), .B2(n_390), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_397), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_397), .Y(n_420) );
A2O1A1Ixp33_ASAP7_75t_L g421 ( .A1(n_400), .A2(n_379), .B(n_391), .C(n_376), .Y(n_421) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_401), .Y(n_422) );
NAND3xp33_ASAP7_75t_L g423 ( .A(n_382), .B(n_385), .C(n_384), .Y(n_423) );
OAI21x1_ASAP7_75t_L g424 ( .A1(n_398), .A2(n_375), .B(n_386), .Y(n_424) );
OAI21x1_ASAP7_75t_L g425 ( .A1(n_375), .A2(n_386), .B(n_404), .Y(n_425) );
OA21x2_ASAP7_75t_L g426 ( .A1(n_379), .A2(n_404), .B(n_387), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_385), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_401), .Y(n_428) );
AO31x2_ASAP7_75t_L g429 ( .A1(n_378), .A2(n_402), .A3(n_403), .B(n_383), .Y(n_429) );
AO31x2_ASAP7_75t_L g430 ( .A1(n_378), .A2(n_382), .A3(n_391), .B(n_342), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_378), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_378), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_402), .B(n_378), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_409), .Y(n_434) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_421), .A2(n_402), .B(n_423), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_406), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_425), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_431), .Y(n_438) );
AO21x2_ASAP7_75t_L g439 ( .A1(n_421), .A2(n_402), .B(n_432), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_424), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_410), .B(n_402), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_412), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_417), .A2(n_416), .B1(n_419), .B2(n_433), .Y(n_443) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_418), .A2(n_433), .B(n_427), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_422), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_417), .A2(n_414), .B1(n_411), .B2(n_418), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_420), .B(n_411), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_415), .Y(n_448) );
OAI221xp5_ASAP7_75t_SL g449 ( .A1(n_405), .A2(n_408), .B1(n_414), .B2(n_413), .C(n_428), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_426), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_422), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_426), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_422), .Y(n_453) );
BUFx3_ASAP7_75t_L g454 ( .A(n_422), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_426), .Y(n_455) );
BUFx4f_ASAP7_75t_L g456 ( .A(n_407), .Y(n_456) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_405), .A2(n_430), .B(n_429), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_407), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_407), .Y(n_459) );
OAI221xp5_ASAP7_75t_L g460 ( .A1(n_429), .A2(n_370), .B1(n_198), .B2(n_215), .C(n_392), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_429), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_429), .Y(n_462) );
OR2x6_ASAP7_75t_L g463 ( .A(n_430), .B(n_427), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_430), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_430), .Y(n_465) );
AND2x4_ASAP7_75t_SL g466 ( .A(n_410), .B(n_409), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_406), .Y(n_467) );
OR2x6_ASAP7_75t_L g468 ( .A(n_427), .B(n_352), .Y(n_468) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_421), .A2(n_424), .B(n_425), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_425), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_441), .B(n_439), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_438), .B(n_441), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_452), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_439), .B(n_464), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_438), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_439), .B(n_464), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_450), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_445), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_466), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_450), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_456), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_452), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_439), .B(n_461), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_452), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_461), .B(n_465), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_455), .B(n_463), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_455), .Y(n_487) );
INVx3_ASAP7_75t_L g488 ( .A(n_456), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_442), .B(n_467), .Y(n_489) );
INVxp67_ASAP7_75t_SL g490 ( .A(n_458), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_442), .B(n_467), .Y(n_491) );
INVxp67_ASAP7_75t_SL g492 ( .A(n_458), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_463), .B(n_457), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_443), .B(n_444), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_458), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_436), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_463), .B(n_457), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_463), .B(n_457), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_459), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_459), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_436), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_447), .B(n_443), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_448), .B(n_434), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_459), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_463), .B(n_457), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_440), .B(n_470), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_435), .B(n_462), .Y(n_507) );
INVx4_ASAP7_75t_L g508 ( .A(n_454), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_447), .B(n_446), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_437), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_435), .B(n_462), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_435), .B(n_444), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_435), .B(n_444), .Y(n_513) );
NOR2x1_ASAP7_75t_SL g514 ( .A(n_468), .B(n_454), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_460), .A2(n_468), .B1(n_444), .B2(n_466), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_451), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_445), .Y(n_517) );
INVx3_ASAP7_75t_L g518 ( .A(n_456), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_469), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_471), .B(n_456), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_472), .B(n_468), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_496), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_471), .B(n_469), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_471), .B(n_469), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_474), .B(n_469), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_472), .B(n_468), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_503), .B(n_466), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_496), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_501), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_474), .B(n_468), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_486), .B(n_454), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_501), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_489), .B(n_460), .Y(n_533) );
INVx4_ASAP7_75t_L g534 ( .A(n_479), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_475), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_475), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_481), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_474), .B(n_453), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_502), .A2(n_449), .B1(n_453), .B2(n_509), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_473), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_516), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_473), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_489), .Y(n_543) );
BUFx2_ASAP7_75t_L g544 ( .A(n_479), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_491), .B(n_449), .Y(n_545) );
OAI31xp33_ASAP7_75t_L g546 ( .A1(n_479), .A2(n_502), .A3(n_515), .B(n_494), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_491), .B(n_472), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_477), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_476), .B(n_483), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_473), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_482), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_509), .B(n_476), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_508), .B(n_514), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_476), .B(n_483), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_477), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_483), .B(n_486), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_480), .B(n_485), .Y(n_557) );
NAND2x1_ASAP7_75t_L g558 ( .A(n_481), .B(n_488), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_480), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_486), .B(n_485), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_485), .B(n_516), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_487), .B(n_493), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_487), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_481), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_514), .B(n_488), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_481), .B(n_488), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_487), .B(n_505), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_517), .Y(n_568) );
INVx4_ASAP7_75t_L g569 ( .A(n_508), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_517), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_482), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_493), .B(n_505), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_494), .B(n_482), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_494), .A2(n_518), .B1(n_488), .B2(n_508), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_484), .B(n_504), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_484), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_478), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_484), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_513), .B(n_515), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_478), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_575), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_561), .B(n_504), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_552), .B(n_513), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_541), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_522), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_560), .B(n_505), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_528), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_529), .Y(n_588) );
OR2x6_ASAP7_75t_L g589 ( .A(n_569), .B(n_518), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_549), .B(n_513), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_569), .B(n_518), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_560), .B(n_497), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_532), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_549), .B(n_507), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_556), .B(n_497), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_535), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_554), .B(n_490), .Y(n_597) );
NAND2x1_ASAP7_75t_L g598 ( .A(n_569), .B(n_508), .Y(n_598) );
INVxp67_ASAP7_75t_SL g599 ( .A(n_540), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_543), .B(n_507), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_547), .B(n_490), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_523), .B(n_507), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_557), .B(n_492), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_575), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_536), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_523), .B(n_512), .Y(n_606) );
INVx2_ASAP7_75t_SL g607 ( .A(n_534), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_556), .B(n_492), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_520), .B(n_498), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_524), .B(n_512), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_527), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_524), .B(n_511), .Y(n_612) );
AOI21xp33_ASAP7_75t_SL g613 ( .A1(n_553), .A2(n_518), .B(n_493), .Y(n_613) );
NOR2x1_ASAP7_75t_L g614 ( .A(n_534), .B(n_508), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_520), .B(n_497), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_540), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_542), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_548), .B(n_511), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_555), .Y(n_619) );
INVxp67_ASAP7_75t_L g620 ( .A(n_577), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_559), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_573), .B(n_498), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_568), .Y(n_623) );
NAND2x1_ASAP7_75t_L g624 ( .A(n_534), .B(n_498), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_539), .A2(n_495), .B1(n_499), .B2(n_500), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_573), .B(n_519), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_572), .B(n_495), .Y(n_627) );
AND2x2_ASAP7_75t_SL g628 ( .A(n_544), .B(n_495), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_572), .B(n_499), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_538), .B(n_499), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_538), .B(n_500), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_570), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_530), .B(n_500), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_565), .B(n_506), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_616), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_584), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_627), .B(n_567), .Y(n_637) );
AND2x4_ASAP7_75t_L g638 ( .A(n_624), .B(n_567), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_583), .B(n_545), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_585), .Y(n_640) );
BUFx2_ASAP7_75t_L g641 ( .A(n_589), .Y(n_641) );
INVx1_ASAP7_75t_SL g642 ( .A(n_611), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_629), .B(n_562), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_607), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_595), .B(n_562), .Y(n_645) );
OAI211xp5_ASAP7_75t_SL g646 ( .A1(n_620), .A2(n_546), .B(n_533), .C(n_579), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_617), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_586), .B(n_525), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_587), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_592), .B(n_531), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_601), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_589), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_620), .B(n_526), .Y(n_653) );
AOI21xp33_ASAP7_75t_L g654 ( .A1(n_625), .A2(n_580), .B(n_574), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_594), .B(n_526), .Y(n_655) );
NOR2xp67_ASAP7_75t_SL g656 ( .A(n_598), .B(n_544), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_588), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_593), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_583), .B(n_525), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_594), .B(n_521), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_596), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_605), .Y(n_662) );
INVx2_ASAP7_75t_SL g663 ( .A(n_589), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_590), .B(n_521), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_619), .Y(n_665) );
INVx2_ASAP7_75t_SL g666 ( .A(n_614), .Y(n_666) );
AND2x2_ASAP7_75t_SL g667 ( .A(n_628), .B(n_565), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_599), .Y(n_668) );
OAI21xp33_ASAP7_75t_L g669 ( .A1(n_590), .A2(n_530), .B(n_580), .Y(n_669) );
INVx1_ASAP7_75t_SL g670 ( .A(n_582), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_625), .A2(n_563), .B1(n_576), .B2(n_571), .C(n_578), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_621), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_623), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_640), .Y(n_674) );
BUFx3_ASAP7_75t_L g675 ( .A(n_666), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_648), .B(n_615), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_639), .B(n_606), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_646), .A2(n_606), .B1(n_610), .B2(n_612), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_668), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_666), .A2(n_628), .B(n_613), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g681 ( .A1(n_667), .A2(n_591), .B(n_565), .C(n_634), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_651), .B(n_610), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_670), .B(n_602), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_649), .Y(n_684) );
NOR2x1_ASAP7_75t_L g685 ( .A(n_641), .B(n_591), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_653), .A2(n_612), .B1(n_609), .B2(n_622), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_659), .B(n_602), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_668), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_657), .Y(n_689) );
INVx2_ASAP7_75t_SL g690 ( .A(n_642), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g691 ( .A1(n_667), .A2(n_634), .B(n_558), .C(n_608), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_658), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_652), .A2(n_622), .B1(n_597), .B2(n_558), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_653), .A2(n_531), .B1(n_566), .B2(n_632), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_661), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_662), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_665), .Y(n_697) );
NAND2xp33_ASAP7_75t_SL g698 ( .A(n_680), .B(n_656), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_691), .A2(n_663), .B1(n_669), .B2(n_644), .C(n_654), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_678), .A2(n_652), .B1(n_663), .B2(n_638), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_681), .A2(n_638), .B(n_671), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_693), .A2(n_638), .B1(n_664), .B2(n_636), .Y(n_702) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_681), .A2(n_664), .B(n_648), .C(n_650), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_674), .Y(n_704) );
OAI211xp5_ASAP7_75t_SL g705 ( .A1(n_690), .A2(n_685), .B(n_691), .C(n_694), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_687), .B(n_660), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_694), .A2(n_673), .B1(n_672), .B2(n_655), .C(n_600), .Y(n_707) );
INVxp67_ASAP7_75t_L g708 ( .A(n_675), .Y(n_708) );
OAI221xp5_ASAP7_75t_SL g709 ( .A1(n_686), .A2(n_600), .B1(n_603), .B2(n_645), .C(n_626), .Y(n_709) );
NAND3xp33_ASAP7_75t_SL g710 ( .A(n_683), .B(n_645), .C(n_643), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_677), .A2(n_633), .B1(n_630), .B2(n_631), .Y(n_711) );
AOI322xp5_ASAP7_75t_L g712 ( .A1(n_698), .A2(n_682), .A3(n_676), .B1(n_637), .B2(n_643), .C1(n_675), .C2(n_692), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_705), .A2(n_697), .B1(n_696), .B2(n_695), .C(n_689), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_699), .A2(n_684), .B1(n_688), .B2(n_679), .C(n_637), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_704), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_700), .A2(n_688), .B1(n_581), .B2(n_604), .Y(n_716) );
O2A1O1Ixp33_ASAP7_75t_L g717 ( .A1(n_708), .A2(n_618), .B(n_647), .C(n_635), .Y(n_717) );
BUFx2_ASAP7_75t_L g718 ( .A(n_703), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_709), .A2(n_626), .B1(n_618), .B2(n_647), .C(n_635), .Y(n_719) );
NAND5xp2_ASAP7_75t_L g720 ( .A(n_712), .B(n_701), .C(n_702), .D(n_707), .E(n_711), .Y(n_720) );
NAND4xp25_ASAP7_75t_L g721 ( .A(n_718), .B(n_710), .C(n_706), .D(n_566), .Y(n_721) );
OAI211xp5_ASAP7_75t_SL g722 ( .A1(n_714), .A2(n_537), .B(n_564), .C(n_599), .Y(n_722) );
NAND3xp33_ASAP7_75t_SL g723 ( .A(n_713), .B(n_519), .C(n_550), .Y(n_723) );
NOR3xp33_ASAP7_75t_L g724 ( .A(n_719), .B(n_537), .C(n_564), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_720), .B(n_716), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_724), .B(n_715), .Y(n_726) );
NOR3xp33_ASAP7_75t_L g727 ( .A(n_721), .B(n_717), .C(n_537), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_726), .Y(n_728) );
XNOR2x2_ASAP7_75t_SL g729 ( .A(n_725), .B(n_723), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_729), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_730), .Y(n_731) );
AOI222xp33_ASAP7_75t_L g732 ( .A1(n_731), .A2(n_728), .B1(n_722), .B2(n_727), .C1(n_566), .C2(n_564), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_732), .A2(n_531), .B(n_510), .Y(n_733) );
OR2x6_ASAP7_75t_L g734 ( .A(n_733), .B(n_551), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_734), .A2(n_551), .B1(n_550), .B2(n_542), .Y(n_735) );
endmodule