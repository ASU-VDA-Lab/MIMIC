module fake_jpeg_14170_n_405 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_405);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_405;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_52),
.B(n_61),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_30),
.B1(n_38),
.B2(n_36),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_62),
.Y(n_91)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_69),
.B(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_23),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_26),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_25),
.B(n_0),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_27),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_74),
.B(n_107),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_76),
.A2(n_36),
.B1(n_38),
.B2(n_33),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_31),
.B1(n_25),
.B2(n_38),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_81),
.A2(n_30),
.B1(n_28),
.B2(n_21),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_35),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_108),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_40),
.A2(n_26),
.B1(n_29),
.B2(n_23),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_102),
.B(n_109),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_40),
.A2(n_26),
.B1(n_29),
.B2(n_23),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_25),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_39),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_45),
.A2(n_26),
.B1(n_23),
.B2(n_31),
.Y(n_109)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

BUFx2_ASAP7_75t_SL g176 ( 
.A(n_113),
.Y(n_176)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_114),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_77),
.Y(n_116)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_118),
.A2(n_131),
.B1(n_147),
.B2(n_30),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_100),
.B(n_106),
.C(n_91),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_139),
.B(n_143),
.Y(n_153)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_141),
.B1(n_35),
.B2(n_36),
.Y(n_155)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_76),
.A2(n_34),
.B1(n_32),
.B2(n_19),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_46),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_136),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_44),
.B(n_57),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_63),
.B(n_59),
.Y(n_163)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_47),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_98),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_31),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_48),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_51),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_148),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_41),
.B1(n_43),
.B2(n_53),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_48),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_145),
.Y(n_167)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_87),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_80),
.A2(n_34),
.B1(n_32),
.B2(n_19),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_104),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_87),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_102),
.A2(n_34),
.B(n_32),
.C(n_35),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_28),
.B(n_33),
.Y(n_165)
);

AO22x1_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_90),
.B1(n_85),
.B2(n_42),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_151),
.B(n_179),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_163),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_54),
.C(n_65),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_174),
.C(n_180),
.Y(n_196)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_99),
.A3(n_23),
.B1(n_50),
.B2(n_104),
.Y(n_161)
);

OR2x2_ASAP7_75t_SL g194 ( 
.A(n_161),
.B(n_150),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_96),
.B1(n_105),
.B2(n_83),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_162),
.A2(n_144),
.B1(n_130),
.B2(n_122),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_165),
.A2(n_166),
.B(n_135),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_119),
.A2(n_28),
.B(n_33),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_136),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_169),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_172),
.A2(n_142),
.B1(n_99),
.B2(n_146),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_115),
.B(n_101),
.C(n_92),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_120),
.A2(n_18),
.B(n_21),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_18),
.B(n_21),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_92),
.C(n_56),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_86),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_148),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_183),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_137),
.B1(n_125),
.B2(n_114),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_197),
.B1(n_201),
.B2(n_160),
.Y(n_229)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_193),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_149),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_199),
.C(n_205),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_183),
.Y(n_191)
);

NAND2xp33_ASAP7_75t_SL g248 ( 
.A(n_191),
.B(n_203),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_218),
.B(n_151),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_134),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_184),
.B(n_159),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_132),
.B1(n_105),
.B2(n_96),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_121),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_200),
.B(n_210),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_209),
.B1(n_191),
.B2(n_185),
.Y(n_230)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_174),
.C(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_145),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_217),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_155),
.A2(n_144),
.B1(n_49),
.B2(n_66),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_181),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_116),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_213),
.Y(n_247)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_160),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g213 ( 
.A(n_153),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_158),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_167),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_SL g216 ( 
.A(n_151),
.B(n_18),
.C(n_129),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_128),
.C(n_123),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

A2O1A1O1Ixp25_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_184),
.B(n_159),
.C(n_152),
.D(n_162),
.Y(n_220)
);

OA21x2_ASAP7_75t_SL g253 ( 
.A1(n_220),
.A2(n_240),
.B(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_221),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_187),
.B1(n_195),
.B2(n_201),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_225),
.A2(n_246),
.B1(n_249),
.B2(n_185),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_207),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_231),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_228),
.A2(n_203),
.B(n_188),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_229),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_274)
);

OA22x2_ASAP7_75t_L g266 ( 
.A1(n_230),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_197),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_167),
.B1(n_177),
.B2(n_152),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_234),
.A2(n_242),
.B1(n_244),
.B2(n_251),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_238),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_176),
.B(n_167),
.C(n_177),
.D(n_129),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_204),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_1),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_192),
.A2(n_154),
.B1(n_156),
.B2(n_86),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_192),
.A2(n_154),
.B1(n_156),
.B2(n_124),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_126),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_250),
.C(n_24),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_195),
.A2(n_113),
.B1(n_117),
.B2(n_75),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_75),
.B1(n_170),
.B2(n_73),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_196),
.B(n_164),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_209),
.A2(n_67),
.B1(n_68),
.B2(n_170),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_252),
.A2(n_263),
.B1(n_271),
.B2(n_274),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_253),
.A2(n_254),
.B(n_257),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_248),
.A2(n_217),
.B(n_194),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_221),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_255),
.B(n_259),
.Y(n_303)
);

OAI22x1_ASAP7_75t_L g257 ( 
.A1(n_219),
.A2(n_206),
.B1(n_214),
.B2(n_199),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_208),
.Y(n_258)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

NAND3xp33_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_215),
.C(n_196),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_260),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_243),
.A2(n_129),
.B(n_164),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_262),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_224),
.B(n_202),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_225),
.A2(n_164),
.B1(n_23),
.B2(n_42),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_164),
.Y(n_265)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_266),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_24),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_272),
.C(n_279),
.Y(n_293)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_236),
.A2(n_24),
.B1(n_3),
.B2(n_4),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_221),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_273),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_233),
.B(n_1),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_235),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_223),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_281),
.B1(n_239),
.B2(n_237),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_228),
.A2(n_5),
.B(n_6),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_278),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_222),
.B(n_250),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_224),
.B(n_5),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_223),
.B(n_6),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_301),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_222),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_290),
.C(n_294),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_245),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_260),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_239),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_238),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_234),
.C(n_249),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_254),
.B(n_246),
.C(n_237),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_230),
.C(n_232),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_302),
.C(n_306),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_265),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_240),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_256),
.A2(n_275),
.B1(n_262),
.B2(n_268),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_304),
.A2(n_263),
.B1(n_242),
.B2(n_231),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_232),
.C(n_227),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_298),
.A2(n_268),
.B1(n_253),
.B2(n_267),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_310),
.A2(n_304),
.B1(n_300),
.B2(n_284),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_280),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_311),
.B(n_317),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_264),
.B(n_261),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_312),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_283),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_328),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_281),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_285),
.Y(n_318)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_255),
.C(n_273),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_325),
.C(n_326),
.Y(n_335)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_301),
.Y(n_320)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_307),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_321),
.B(n_322),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_289),
.A2(n_264),
.B(n_252),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_323),
.A2(n_291),
.B1(n_284),
.B2(n_297),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g324 ( 
.A1(n_282),
.A2(n_274),
.B(n_241),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_293),
.B(n_227),
.C(n_244),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_256),
.C(n_243),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_277),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_327),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_283),
.A2(n_278),
.B(n_251),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_303),
.B(n_266),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_329),
.A2(n_271),
.B1(n_266),
.B2(n_220),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_295),
.C(n_290),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_292),
.C(n_286),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_338),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_332),
.A2(n_319),
.B1(n_313),
.B2(n_314),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_309),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_347),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_334),
.A2(n_336),
.B1(n_347),
.B2(n_344),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_309),
.A2(n_310),
.B1(n_328),
.B2(n_312),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_336),
.A2(n_323),
.B1(n_266),
.B2(n_8),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_302),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_343),
.B(n_348),
.Y(n_349)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_341),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_316),
.C(n_326),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_351),
.B(n_352),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_335),
.B(n_313),
.C(n_325),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_346),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_353),
.A2(n_354),
.B1(n_340),
.B2(n_338),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_337),
.B(n_314),
.Y(n_356)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_356),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_330),
.Y(n_357)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_357),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_308),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_359),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_315),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_360),
.A2(n_362),
.B(n_340),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_332),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_SL g362 ( 
.A(n_343),
.B(n_6),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_14),
.B1(n_7),
.B2(n_8),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_341),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_368),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_366),
.B(n_367),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_331),
.C(n_333),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_8),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_372),
.B(n_6),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_339),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_374),
.B(n_363),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_350),
.A2(n_349),
.B(n_351),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_375),
.A2(n_10),
.B(n_11),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_355),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_376),
.A2(n_385),
.B(n_366),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_371),
.A2(n_358),
.B(n_361),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_377),
.A2(n_372),
.B(n_370),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_379),
.B(n_383),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_381),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_9),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_9),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_11),
.Y(n_393)
);

BUFx24_ASAP7_75t_SL g386 ( 
.A(n_382),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_386),
.B(n_387),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_378),
.B(n_368),
.C(n_374),
.Y(n_388)
);

MAJx2_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_380),
.C(n_13),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_12),
.C(n_14),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_378),
.A2(n_11),
.B(n_12),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_392),
.A2(n_12),
.B(n_13),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_393),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_394),
.B(n_390),
.C(n_391),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_395),
.B(n_398),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_400),
.A2(n_401),
.B(n_397),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_396),
.Y(n_401)
);

BUFx24_ASAP7_75t_SL g403 ( 
.A(n_402),
.Y(n_403)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_403),
.Y(n_404)
);

AOI21x1_ASAP7_75t_L g405 ( 
.A1(n_404),
.A2(n_399),
.B(n_12),
.Y(n_405)
);


endmodule