module fake_aes_3051_n_629 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_629);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_629;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g70 ( .A(n_39), .Y(n_70) );
NOR2xp33_ASAP7_75t_L g71 ( .A(n_22), .B(n_32), .Y(n_71) );
CKINVDCx5p33_ASAP7_75t_R g72 ( .A(n_58), .Y(n_72) );
INVxp33_ASAP7_75t_SL g73 ( .A(n_35), .Y(n_73) );
INVxp67_ASAP7_75t_SL g74 ( .A(n_30), .Y(n_74) );
BUFx2_ASAP7_75t_L g75 ( .A(n_54), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_31), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_42), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_64), .Y(n_78) );
INVxp33_ASAP7_75t_L g79 ( .A(n_48), .Y(n_79) );
INVxp67_ASAP7_75t_L g80 ( .A(n_49), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_69), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_52), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_63), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_27), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_34), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_12), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_62), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_3), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_65), .Y(n_89) );
BUFx2_ASAP7_75t_L g90 ( .A(n_55), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_18), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_14), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_33), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_36), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_51), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_40), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_67), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_13), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_20), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_3), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_7), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_12), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_57), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_8), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_47), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_59), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_45), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_18), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_14), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_60), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_4), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_61), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_13), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_53), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_66), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_50), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_11), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_106), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_75), .B(n_0), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_70), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_83), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_70), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g124 ( .A(n_75), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_76), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_77), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_90), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_77), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g129 ( .A(n_90), .B(n_0), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_78), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_88), .B(n_1), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_86), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_108), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_78), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_81), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_79), .B(n_1), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_85), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_85), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_88), .B(n_2), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_92), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_101), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_98), .Y(n_145) );
BUFx10_ASAP7_75t_L g146 ( .A(n_72), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_87), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_87), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_111), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_98), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_102), .B(n_2), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_89), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
BUFx2_ASAP7_75t_L g155 ( .A(n_102), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_109), .B(n_4), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_93), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_95), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_109), .B(n_5), .Y(n_159) );
CKINVDCx16_ASAP7_75t_R g160 ( .A(n_96), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_157), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_157), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_157), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_127), .B(n_80), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_155), .B(n_117), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_124), .B(n_73), .Y(n_166) );
INVx8_ASAP7_75t_L g167 ( .A(n_131), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_155), .B(n_117), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_160), .B(n_105), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_157), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_146), .Y(n_171) );
AND2x6_ASAP7_75t_L g172 ( .A(n_131), .B(n_97), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_157), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_124), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_157), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_146), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_120), .A2(n_107), .B(n_96), .C(n_103), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_119), .B(n_91), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_122), .Y(n_181) );
OR2x2_ASAP7_75t_L g182 ( .A(n_160), .B(n_100), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_122), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_138), .B(n_99), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_122), .Y(n_185) );
INVxp67_ASAP7_75t_SL g186 ( .A(n_119), .Y(n_186) );
NOR2x1_ASAP7_75t_L g187 ( .A(n_120), .B(n_115), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_122), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_138), .B(n_94), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_132), .B(n_114), .Y(n_192) );
CKINVDCx8_ASAP7_75t_R g193 ( .A(n_118), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_130), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_131), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_136), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_130), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_119), .B(n_113), .Y(n_198) );
AO22x2_ASAP7_75t_L g199 ( .A1(n_131), .A2(n_103), .B1(n_112), .B2(n_107), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_131), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_136), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_133), .B(n_97), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_145), .B(n_104), .Y(n_203) );
NOR2xp33_ASAP7_75t_SL g204 ( .A(n_149), .B(n_110), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_130), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_130), .Y(n_206) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_121), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_145), .B(n_112), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_138), .B(n_82), .Y(n_209) );
INVxp67_ASAP7_75t_L g210 ( .A(n_159), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_142), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_123), .B(n_93), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_151), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_135), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_135), .B(n_116), .Y(n_215) );
INVx2_ASAP7_75t_SL g216 ( .A(n_135), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_135), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_123), .B(n_74), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_140), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_140), .Y(n_220) );
AO22x2_ASAP7_75t_L g221 ( .A1(n_129), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_140), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_217), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_174), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_186), .B(n_159), .Y(n_225) );
NAND3xp33_ASAP7_75t_SL g226 ( .A(n_174), .B(n_144), .C(n_129), .Y(n_226) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_213), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_208), .B(n_148), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_211), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_217), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_195), .B(n_140), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_217), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_181), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_171), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_196), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_195), .B(n_150), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_181), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_195), .B(n_150), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_211), .Y(n_239) );
INVx2_ASAP7_75t_SL g240 ( .A(n_198), .Y(n_240) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_213), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_198), .B(n_159), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_167), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_183), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_183), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_185), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_184), .B(n_158), .Y(n_247) );
OAI22xp5_ASAP7_75t_SL g248 ( .A1(n_193), .A2(n_141), .B1(n_156), .B2(n_152), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_210), .A2(n_141), .B(n_156), .C(n_152), .Y(n_249) );
INVx4_ASAP7_75t_L g250 ( .A(n_167), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_207), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_195), .B(n_150), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_185), .Y(n_253) );
INVx5_ASAP7_75t_L g254 ( .A(n_172), .Y(n_254) );
OR2x2_ASAP7_75t_L g255 ( .A(n_182), .B(n_158), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_167), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_208), .B(n_154), .Y(n_257) );
OR2x6_ASAP7_75t_L g258 ( .A(n_167), .B(n_154), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_196), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_203), .B(n_137), .Y(n_260) );
INVx2_ASAP7_75t_SL g261 ( .A(n_198), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_188), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_198), .B(n_137), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_200), .A2(n_125), .B(n_134), .C(n_148), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_190), .B(n_139), .Y(n_265) );
BUFx4f_ASAP7_75t_L g266 ( .A(n_172), .Y(n_266) );
NOR2xp33_ASAP7_75t_R g267 ( .A(n_193), .B(n_153), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_199), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_196), .Y(n_269) );
NOR3xp33_ASAP7_75t_SL g270 ( .A(n_166), .B(n_125), .C(n_126), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_199), .A2(n_147), .B1(n_126), .B2(n_139), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_188), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_182), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_179), .B(n_147), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_171), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_194), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_167), .A2(n_134), .B(n_128), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_194), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_197), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_197), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_205), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_209), .B(n_128), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_196), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_209), .B(n_153), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_215), .B(n_153), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_196), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_205), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_215), .B(n_153), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_243), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_224), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_250), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_258), .A2(n_199), .B1(n_200), .B2(n_215), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_231), .A2(n_177), .B(n_199), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_268), .A2(n_242), .B1(n_240), .B2(n_261), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_263), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_287), .Y(n_296) );
INVx2_ASAP7_75t_SL g297 ( .A(n_258), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_233), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_258), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_242), .B(n_203), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_225), .B(n_179), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_287), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_250), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_248), .A2(n_172), .B1(n_164), .B2(n_204), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_224), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_237), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_251), .Y(n_307) );
OAI22xp5_ASAP7_75t_SL g308 ( .A1(n_229), .A2(n_169), .B1(n_221), .B2(n_215), .Y(n_308) );
BUFx12f_ASAP7_75t_L g309 ( .A(n_229), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_243), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_250), .B(n_165), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g312 ( .A1(n_264), .A2(n_178), .B(n_168), .C(n_165), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_242), .B(n_168), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_225), .A2(n_172), .B1(n_221), .B2(n_218), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_244), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_282), .A2(n_172), .B1(n_202), .B2(n_180), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_225), .B(n_172), .Y(n_317) );
INVx3_ASAP7_75t_SL g318 ( .A(n_239), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_243), .Y(n_319) );
INVx6_ASAP7_75t_L g320 ( .A(n_243), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_254), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_256), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_227), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_263), .B(n_187), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_263), .B(n_187), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_256), .Y(n_326) );
INVx5_ASAP7_75t_L g327 ( .A(n_254), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_266), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_282), .B(n_172), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_274), .B(n_228), .Y(n_330) );
INVx4_ASAP7_75t_SL g331 ( .A(n_234), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_245), .Y(n_332) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_264), .A2(n_212), .B(n_162), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_274), .B(n_180), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_274), .B(n_189), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_246), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_266), .A2(n_191), .B1(n_189), .B2(n_221), .Y(n_337) );
OAI21xp33_ASAP7_75t_L g338 ( .A1(n_247), .A2(n_191), .B(n_177), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_L g339 ( .A1(n_273), .A2(n_222), .B(n_206), .C(n_220), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_311), .A2(n_226), .B1(n_241), .B2(n_255), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_305), .B(n_257), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_298), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_307), .B(n_260), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_311), .A2(n_265), .B1(n_247), .B2(n_284), .Y(n_344) );
AOI222xp33_ASAP7_75t_SL g345 ( .A1(n_308), .A2(n_150), .B1(n_143), .B2(n_136), .C1(n_221), .C2(n_201), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_311), .B(n_265), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_296), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_298), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_313), .A2(n_231), .B1(n_252), .B2(n_238), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_330), .B(n_249), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_306), .B(n_270), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_299), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_329), .A2(n_277), .B(n_236), .Y(n_353) );
AOI21xp33_ASAP7_75t_L g354 ( .A1(n_337), .A2(n_271), .B(n_234), .Y(n_354) );
NAND3x1_ASAP7_75t_L g355 ( .A(n_304), .B(n_71), .C(n_267), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_306), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_292), .A2(n_288), .B1(n_285), .B2(n_272), .Y(n_357) );
CKINVDCx14_ASAP7_75t_R g358 ( .A(n_290), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_293), .A2(n_235), .B(n_259), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_296), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_319), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_313), .A2(n_238), .B1(n_236), .B2(n_252), .Y(n_362) );
OAI22xp33_ASAP7_75t_L g363 ( .A1(n_307), .A2(n_290), .B1(n_318), .B2(n_323), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_301), .B(n_223), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_315), .Y(n_365) );
BUFx2_ASAP7_75t_SL g366 ( .A(n_327), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_300), .A2(n_267), .B1(n_192), .B2(n_222), .C(n_220), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_299), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_297), .B(n_254), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_302), .Y(n_370) );
OA21x2_ASAP7_75t_L g371 ( .A1(n_314), .A2(n_176), .B(n_175), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_342), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_346), .B(n_300), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_357), .A2(n_297), .B1(n_334), .B2(n_294), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_361), .Y(n_375) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_357), .B(n_334), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_361), .Y(n_377) );
OAI211xp5_ASAP7_75t_L g378 ( .A1(n_340), .A2(n_312), .B(n_339), .C(n_316), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_346), .B(n_335), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_343), .A2(n_309), .B1(n_334), .B2(n_335), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_351), .A2(n_309), .B1(n_318), .B2(n_324), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_341), .A2(n_295), .B1(n_317), .B2(n_338), .C(n_325), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_342), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_348), .B(n_315), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_351), .A2(n_325), .B1(n_324), .B2(n_332), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_345), .A2(n_344), .B1(n_350), .B2(n_363), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_350), .A2(n_336), .B1(n_332), .B2(n_302), .Y(n_387) );
AO221x2_ASAP7_75t_L g388 ( .A1(n_345), .A2(n_336), .B1(n_8), .B2(n_9), .C(n_10), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_355), .A2(n_275), .B1(n_291), .B2(n_303), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_348), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_352), .A2(n_291), .B1(n_303), .B2(n_322), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_358), .A2(n_326), .B1(n_322), .B2(n_333), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_356), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_367), .A2(n_326), .B1(n_333), .B2(n_291), .Y(n_394) );
AOI222xp33_ASAP7_75t_L g395 ( .A1(n_356), .A2(n_279), .B1(n_281), .B2(n_253), .C1(n_262), .C2(n_276), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_352), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_347), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_368), .A2(n_326), .B1(n_333), .B2(n_303), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_365), .B(n_310), .Y(n_399) );
NAND4xp25_ASAP7_75t_SL g400 ( .A(n_381), .B(n_365), .C(n_354), .D(n_355), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_376), .A2(n_354), .B1(n_370), .B2(n_347), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_385), .A2(n_349), .B1(n_362), .B2(n_368), .C(n_364), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_397), .Y(n_403) );
NAND3xp33_ASAP7_75t_L g404 ( .A(n_388), .B(n_371), .C(n_370), .Y(n_404) );
OAI222xp33_ASAP7_75t_L g405 ( .A1(n_386), .A2(n_347), .B1(n_360), .B2(n_370), .C1(n_364), .C2(n_361), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_376), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_372), .B(n_360), .Y(n_407) );
AO21x2_ASAP7_75t_L g408 ( .A1(n_387), .A2(n_359), .B(n_353), .Y(n_408) );
AND2x6_ASAP7_75t_SL g409 ( .A(n_373), .B(n_369), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_376), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_372), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g412 ( .A1(n_378), .A2(n_359), .B(n_371), .Y(n_412) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_397), .Y(n_413) );
OAI21x1_ASAP7_75t_SL g414 ( .A1(n_383), .A2(n_371), .B(n_360), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_384), .B(n_361), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_384), .B(n_371), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_396), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_388), .A2(n_366), .B1(n_289), .B2(n_369), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_383), .Y(n_419) );
NAND3xp33_ASAP7_75t_SL g420 ( .A(n_392), .B(n_143), .C(n_201), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_397), .B(n_390), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_390), .B(n_393), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_386), .B(n_310), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_393), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_379), .A2(n_143), .B1(n_216), .B2(n_219), .C(n_206), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_375), .Y(n_426) );
AO21x2_ASAP7_75t_L g427 ( .A1(n_391), .A2(n_162), .B(n_175), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_379), .B(n_366), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_395), .B(n_278), .Y(n_429) );
OAI211xp5_ASAP7_75t_SL g430 ( .A1(n_380), .A2(n_176), .B(n_214), .C(n_219), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_388), .B(n_369), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_388), .B(n_289), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_399), .B(n_374), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_398), .B(n_394), .C(n_395), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_411), .B(n_377), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_419), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_419), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_403), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_416), .B(n_375), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_416), .B(n_375), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_424), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_403), .B(n_375), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_421), .B(n_377), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_424), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_421), .B(n_377), .Y(n_446) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_404), .B(n_377), .Y(n_447) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_413), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_415), .B(n_6), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_422), .B(n_389), .Y(n_450) );
INVx2_ASAP7_75t_SL g451 ( .A(n_426), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_422), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_415), .B(n_9), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_414), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_406), .B(n_10), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_406), .B(n_11), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_409), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_414), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_408), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_410), .B(n_15), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_408), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_407), .B(n_382), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_426), .B(n_331), .Y(n_463) );
OAI31xp33_ASAP7_75t_L g464 ( .A1(n_400), .A2(n_275), .A3(n_369), .B(n_216), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_408), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_407), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_433), .B(n_214), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_410), .B(n_15), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_431), .B(n_16), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_433), .B(n_16), .Y(n_470) );
INVx3_ASAP7_75t_L g471 ( .A(n_426), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_409), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_404), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_431), .B(n_331), .Y(n_474) );
AOI211xp5_ASAP7_75t_L g475 ( .A1(n_405), .A2(n_319), .B(n_232), .C(n_230), .Y(n_475) );
CKINVDCx8_ASAP7_75t_R g476 ( .A(n_418), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g477 ( .A(n_434), .B(n_319), .C(n_163), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_428), .B(n_17), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_401), .B(n_331), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_401), .B(n_331), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_412), .A2(n_319), .B(n_254), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_434), .B(n_17), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_427), .Y(n_483) );
NOR3xp33_ASAP7_75t_L g484 ( .A(n_482), .B(n_417), .C(n_402), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_454), .Y(n_485) );
INVx2_ASAP7_75t_SL g486 ( .A(n_436), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_472), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_437), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g489 ( .A1(n_482), .A2(n_429), .B1(n_423), .B2(n_412), .C(n_430), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_440), .B(n_428), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_448), .B(n_432), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_452), .B(n_432), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_472), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_440), .B(n_427), .Y(n_494) );
NAND2x1p5_ASAP7_75t_SL g495 ( .A(n_447), .B(n_427), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_441), .B(n_19), .Y(n_496) );
NOR4xp25_ASAP7_75t_SL g497 ( .A(n_457), .B(n_425), .C(n_420), .D(n_19), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_437), .Y(n_498) );
NAND2xp33_ASAP7_75t_R g499 ( .A(n_457), .B(n_21), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_438), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_439), .Y(n_501) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_469), .A2(n_320), .B1(n_319), .B2(n_321), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_444), .B(n_173), .Y(n_503) );
OAI31xp33_ASAP7_75t_L g504 ( .A1(n_470), .A2(n_321), .A3(n_280), .B(n_232), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_442), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_446), .B(n_173), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_446), .B(n_170), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_442), .B(n_170), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_448), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_475), .A2(n_327), .B(n_328), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_445), .B(n_443), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_478), .Y(n_512) );
NAND2xp33_ASAP7_75t_SL g513 ( .A(n_460), .B(n_328), .Y(n_513) );
NAND2xp33_ASAP7_75t_L g514 ( .A(n_460), .B(n_328), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_435), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_443), .B(n_163), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_478), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_451), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_443), .B(n_161), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_469), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_458), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_449), .B(n_161), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_451), .B(n_23), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g524 ( .A(n_460), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_449), .B(n_230), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_458), .B(n_24), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_439), .B(n_25), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_453), .B(n_223), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_439), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_453), .B(n_320), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_476), .Y(n_531) );
BUFx2_ASAP7_75t_SL g532 ( .A(n_487), .Y(n_532) );
OAI221xp5_ASAP7_75t_SL g533 ( .A1(n_504), .A2(n_464), .B1(n_468), .B2(n_456), .C(n_455), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_488), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_524), .A2(n_476), .B1(n_475), .B2(n_455), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_488), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_498), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_520), .A2(n_476), .B1(n_456), .B2(n_468), .Y(n_538) );
OAI21xp33_ASAP7_75t_L g539 ( .A1(n_520), .A2(n_447), .B(n_473), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_484), .A2(n_462), .B1(n_466), .B2(n_474), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_531), .A2(n_462), .B1(n_474), .B2(n_467), .Y(n_541) );
OAI222xp33_ASAP7_75t_L g542 ( .A1(n_512), .A2(n_483), .B1(n_479), .B2(n_480), .C1(n_454), .C2(n_473), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_500), .Y(n_543) );
XNOR2x1_ASAP7_75t_L g544 ( .A(n_493), .B(n_467), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_531), .A2(n_450), .B1(n_480), .B2(n_479), .Y(n_545) );
AOI21xp33_ASAP7_75t_L g546 ( .A1(n_499), .A2(n_464), .B(n_483), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_509), .Y(n_547) );
INVxp33_ASAP7_75t_L g548 ( .A(n_496), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_517), .B(n_511), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_509), .B(n_471), .Y(n_550) );
NOR4xp25_ASAP7_75t_SL g551 ( .A(n_513), .B(n_477), .C(n_465), .D(n_459), .Y(n_551) );
AOI321xp33_ASAP7_75t_SL g552 ( .A1(n_497), .A2(n_473), .A3(n_465), .B1(n_461), .B2(n_459), .C(n_38), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_500), .Y(n_553) );
O2A1O1Ixp33_ASAP7_75t_L g554 ( .A1(n_514), .A2(n_459), .B(n_465), .C(n_461), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_514), .A2(n_481), .B(n_454), .Y(n_555) );
OAI21xp33_ASAP7_75t_SL g556 ( .A1(n_491), .A2(n_471), .B(n_481), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_486), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_489), .A2(n_463), .B1(n_461), .B2(n_471), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_505), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_513), .A2(n_327), .B(n_283), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_526), .B(n_327), .Y(n_561) );
NOR2xp67_ASAP7_75t_SL g562 ( .A(n_523), .B(n_327), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_515), .B(n_26), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_486), .Y(n_564) );
AOI322xp5_ASAP7_75t_L g565 ( .A1(n_496), .A2(n_28), .A3(n_29), .B1(n_37), .B2(n_41), .C1(n_43), .C2(n_44), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_L g566 ( .A1(n_526), .A2(n_286), .B(n_269), .C(n_259), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_510), .A2(n_283), .B(n_328), .Y(n_567) );
XNOR2x1_ASAP7_75t_L g568 ( .A(n_490), .B(n_46), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g569 ( .A1(n_491), .A2(n_320), .B1(n_328), .B2(n_283), .Y(n_569) );
XNOR2xp5_ASAP7_75t_L g570 ( .A(n_544), .B(n_502), .Y(n_570) );
NOR4xp25_ASAP7_75t_SL g571 ( .A(n_561), .B(n_521), .C(n_515), .D(n_495), .Y(n_571) );
INVxp67_ASAP7_75t_L g572 ( .A(n_532), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_566), .A2(n_518), .B(n_523), .Y(n_573) );
NAND2xp33_ASAP7_75t_SL g574 ( .A(n_548), .B(n_494), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g575 ( .A1(n_533), .A2(n_492), .B1(n_528), .B2(n_525), .C(n_530), .Y(n_575) );
XOR2xp5_ASAP7_75t_L g576 ( .A(n_568), .B(n_494), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_549), .B(n_522), .Y(n_577) );
O2A1O1Ixp33_ASAP7_75t_SL g578 ( .A1(n_546), .A2(n_527), .B(n_485), .C(n_529), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_566), .A2(n_527), .B(n_501), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_559), .Y(n_580) );
XOR2x2_ASAP7_75t_L g581 ( .A(n_538), .B(n_507), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_557), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_540), .B(n_506), .Y(n_583) );
CKINVDCx20_ASAP7_75t_L g584 ( .A(n_562), .Y(n_584) );
AND2x2_ASAP7_75t_SL g585 ( .A(n_558), .B(n_495), .Y(n_585) );
XOR2x2_ASAP7_75t_L g586 ( .A(n_533), .B(n_503), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_550), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_534), .B(n_508), .Y(n_588) );
XOR2x2_ASAP7_75t_L g589 ( .A(n_535), .B(n_519), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_536), .B(n_508), .Y(n_590) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_547), .B(n_564), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_537), .B(n_516), .Y(n_592) );
INVxp67_ASAP7_75t_SL g593 ( .A(n_554), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_591), .B(n_539), .Y(n_594) );
INVxp67_ASAP7_75t_L g595 ( .A(n_572), .Y(n_595) );
XOR2x2_ASAP7_75t_L g596 ( .A(n_570), .B(n_541), .Y(n_596) );
OAI21xp33_ASAP7_75t_SL g597 ( .A1(n_585), .A2(n_560), .B(n_555), .Y(n_597) );
OAI21xp33_ASAP7_75t_L g598 ( .A1(n_593), .A2(n_556), .B(n_545), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_578), .A2(n_542), .B(n_567), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_575), .A2(n_542), .B1(n_553), .B2(n_543), .C(n_554), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_582), .Y(n_601) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_584), .B(n_563), .Y(n_602) );
NAND4xp25_ASAP7_75t_L g603 ( .A(n_583), .B(n_565), .C(n_552), .D(n_569), .Y(n_603) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_587), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_580), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_574), .B(n_551), .C(n_516), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_592), .Y(n_607) );
BUFx2_ASAP7_75t_L g608 ( .A(n_604), .Y(n_608) );
AO22x2_ASAP7_75t_L g609 ( .A1(n_595), .A2(n_576), .B1(n_573), .B2(n_579), .Y(n_609) );
AOI222xp33_ASAP7_75t_L g610 ( .A1(n_596), .A2(n_586), .B1(n_581), .B2(n_589), .C1(n_577), .C2(n_592), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_594), .A2(n_571), .B1(n_588), .B2(n_590), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_600), .B(n_607), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_598), .A2(n_320), .B1(n_235), .B2(n_283), .C(n_56), .Y(n_613) );
XOR2x2_ASAP7_75t_L g614 ( .A(n_602), .B(n_68), .Y(n_614) );
XOR2xp5_ASAP7_75t_L g615 ( .A(n_603), .B(n_606), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_L g616 ( .A1(n_605), .A2(n_597), .B(n_598), .C(n_595), .Y(n_616) );
NAND4xp75_ASAP7_75t_L g617 ( .A(n_602), .B(n_597), .C(n_594), .D(n_600), .Y(n_617) );
AOI22x1_ASAP7_75t_L g618 ( .A1(n_599), .A2(n_570), .B1(n_532), .B2(n_601), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_614), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_610), .B(n_612), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_608), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_621), .Y(n_622) );
OA22x2_ASAP7_75t_L g623 ( .A1(n_620), .A2(n_615), .B1(n_611), .B2(n_617), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_619), .A2(n_618), .B1(n_609), .B2(n_613), .Y(n_624) );
BUFx2_ASAP7_75t_L g625 ( .A(n_622), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_623), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_625), .Y(n_627) );
OAI31xp33_ASAP7_75t_L g628 ( .A1(n_627), .A2(n_626), .A3(n_625), .B(n_616), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_628), .A2(n_624), .B(n_619), .Y(n_629) );
endmodule