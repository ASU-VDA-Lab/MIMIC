module fake_netlist_6_925_n_1540 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1540);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1540;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_167;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_302;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1240;

INVxp67_ASAP7_75t_L g146 ( 
.A(n_46),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_73),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_56),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_1),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_31),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_96),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_16),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_20),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_61),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_45),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_9),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_0),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_19),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_112),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_44),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_4),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_100),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_7),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_39),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_106),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_127),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_24),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_37),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_50),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_80),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_97),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_36),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_5),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_134),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_63),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_64),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_74),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_24),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_107),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_82),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_37),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_142),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_109),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_11),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_143),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_99),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_10),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_84),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_98),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_123),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_55),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_49),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_59),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_136),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_138),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_14),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_94),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_101),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_124),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_110),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_32),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_93),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_35),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_28),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_77),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_25),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_69),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_60),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_40),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_32),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_76),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_1),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_39),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_44),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_48),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_108),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_70),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_75),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_129),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_25),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_28),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_65),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_122),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_95),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_29),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_104),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_111),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_137),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_35),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_36),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_131),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_86),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_19),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_135),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_51),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_27),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_141),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_17),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_38),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_12),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_114),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_38),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_12),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_49),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_41),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_20),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_14),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_13),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_4),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_6),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_121),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_113),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_88),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_21),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_33),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_40),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_52),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_27),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_30),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_11),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_43),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_81),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_92),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_62),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_120),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_132),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_78),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_116),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_144),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_43),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_58),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_91),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_89),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_87),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_237),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_237),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_237),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_174),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_237),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_159),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_175),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_237),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_181),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_184),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_208),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_189),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_208),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_190),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_208),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_185),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_208),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_192),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_193),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_208),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_173),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_164),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_266),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_146),
.B(n_0),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_210),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_164),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_198),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_200),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_205),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_172),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_172),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_194),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_206),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_194),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_187),
.B(n_2),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_251),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_251),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_260),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_209),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_214),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_195),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_216),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_219),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_223),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_232),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_216),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_234),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_176),
.B(n_2),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_151),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_148),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_152),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_236),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_186),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_221),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_242),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_148),
.B(n_165),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_238),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_240),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_156),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_162),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_177),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_201),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_182),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_221),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_291),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g356 ( 
.A(n_294),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_289),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_324),
.A2(n_161),
.B1(n_226),
.B2(n_259),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_300),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_289),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_298),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_165),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_346),
.B(n_204),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_299),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_301),
.B(n_204),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_296),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_306),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_302),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_296),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_303),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_306),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_307),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_304),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_308),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_304),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_309),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_316),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_293),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_317),
.B(n_229),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_287),
.Y(n_382)
);

OAI21x1_ASAP7_75t_L g383 ( 
.A1(n_287),
.A2(n_231),
.B(n_154),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_305),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_288),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_309),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_318),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_322),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_288),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_328),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_290),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_290),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_R g393 ( 
.A(n_330),
.B(n_263),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_314),
.B(n_271),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_292),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_345),
.A2(n_168),
.B1(n_166),
.B2(n_218),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_333),
.B(n_229),
.Y(n_397)
);

NAND2xp33_ASAP7_75t_R g398 ( 
.A(n_334),
.B(n_149),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_292),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_295),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_295),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_337),
.B(n_176),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_342),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_297),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_297),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_339),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_347),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_348),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_339),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_341),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_340),
.B(n_338),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_350),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_350),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_332),
.B(n_211),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_343),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_332),
.B(n_211),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_312),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_331),
.Y(n_418)
);

AND3x2_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_349),
.C(n_155),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_386),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_380),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_331),
.Y(n_422)
);

OAI22xp33_ASAP7_75t_L g423 ( 
.A1(n_359),
.A2(n_335),
.B1(n_255),
.B2(n_178),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_386),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g425 ( 
.A(n_396),
.Y(n_425)
);

AND2x2_ASAP7_75t_SL g426 ( 
.A(n_394),
.B(n_180),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_364),
.B(n_150),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_367),
.B(n_314),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_369),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_381),
.B(n_180),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_397),
.B(n_180),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_364),
.B(n_312),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_369),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_393),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_355),
.B(n_180),
.Y(n_436)
);

BUFx4f_ASAP7_75t_L g437 ( 
.A(n_414),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_395),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_365),
.B(n_310),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_395),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_362),
.B(n_180),
.Y(n_441)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_377),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_400),
.Y(n_443)
);

BUFx8_ASAP7_75t_SL g444 ( 
.A(n_384),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_401),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_414),
.A2(n_207),
.B1(n_245),
.B2(n_215),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_365),
.B(n_344),
.Y(n_447)
);

AND2x6_ASAP7_75t_L g448 ( 
.A(n_401),
.B(n_217),
.Y(n_448)
);

INVx5_ASAP7_75t_L g449 ( 
.A(n_377),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_344),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_366),
.B(n_217),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_382),
.B(n_199),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_372),
.B(n_217),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_336),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_382),
.B(n_220),
.Y(n_456)
);

OR2x6_ASAP7_75t_L g457 ( 
.A(n_416),
.B(n_313),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_361),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_385),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_359),
.B(n_354),
.Y(n_462)
);

BUFx4f_ASAP7_75t_L g463 ( 
.A(n_416),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_416),
.B(n_336),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_368),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_383),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_369),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_391),
.Y(n_469)
);

OR2x6_ASAP7_75t_L g470 ( 
.A(n_416),
.B(n_188),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_383),
.A2(n_213),
.B1(n_248),
.B2(n_270),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_374),
.B(n_351),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_376),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_379),
.B(n_217),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_391),
.Y(n_475)
);

OR2x6_ASAP7_75t_L g476 ( 
.A(n_406),
.B(n_197),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_415),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_392),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_387),
.B(n_352),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_369),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_388),
.B(n_351),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_390),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_403),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_407),
.B(n_353),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_408),
.B(n_235),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_399),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_356),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_358),
.B(n_353),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_SL g490 ( 
.A(n_406),
.B(n_276),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_399),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_396),
.B(n_311),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_358),
.B(n_275),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_369),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_356),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_404),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_409),
.A2(n_267),
.B1(n_272),
.B2(n_202),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_356),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_368),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_404),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_369),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_360),
.B(n_149),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_368),
.Y(n_503)
);

AND2x4_ASAP7_75t_SL g504 ( 
.A(n_409),
.B(n_271),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_410),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_360),
.B(n_153),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_405),
.B(n_235),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_405),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_413),
.B(n_235),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_412),
.B(n_311),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_412),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_371),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_363),
.B(n_153),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_371),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_413),
.A2(n_235),
.B1(n_239),
.B2(n_285),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_357),
.B(n_363),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_378),
.B(n_235),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_357),
.B(n_243),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_378),
.A2(n_239),
.B1(n_286),
.B2(n_249),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_357),
.B(n_244),
.Y(n_520)
);

OR2x6_ASAP7_75t_L g521 ( 
.A(n_370),
.B(n_147),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_377),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_370),
.B(n_157),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_375),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_371),
.A2(n_239),
.B1(n_230),
.B2(n_228),
.Y(n_525)
);

AND2x2_ASAP7_75t_SL g526 ( 
.A(n_373),
.B(n_239),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_389),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_402),
.B(n_246),
.Y(n_528)
);

AO21x2_ASAP7_75t_L g529 ( 
.A1(n_411),
.A2(n_196),
.B(n_203),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_411),
.B(n_315),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_411),
.A2(n_252),
.B1(n_183),
.B2(n_222),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_402),
.B(n_253),
.Y(n_532)
);

INVx4_ASAP7_75t_SL g533 ( 
.A(n_369),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_364),
.Y(n_534)
);

INVx5_ASAP7_75t_L g535 ( 
.A(n_377),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_361),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_364),
.B(n_239),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_422),
.B(n_157),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_422),
.B(n_160),
.Y(n_539)
);

INVx8_ASAP7_75t_L g540 ( 
.A(n_457),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_444),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_505),
.B(n_271),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_453),
.A2(n_163),
.B(n_264),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_438),
.B(n_169),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_511),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_417),
.B(n_160),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_440),
.B(n_179),
.Y(n_547)
);

A2O1A1Ixp33_ASAP7_75t_L g548 ( 
.A1(n_437),
.A2(n_212),
.B(n_247),
.C(n_265),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_510),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_461),
.B(n_472),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_437),
.B(n_281),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_435),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_443),
.B(n_167),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_439),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_456),
.A2(n_329),
.B(n_327),
.Y(n_555)
);

BUFx6f_ASAP7_75t_SL g556 ( 
.A(n_473),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_445),
.B(n_171),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_475),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_433),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_504),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_527),
.B(n_269),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_472),
.B(n_269),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_L g563 ( 
.A(n_418),
.B(n_274),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_534),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_475),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_481),
.B(n_277),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_420),
.B(n_277),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_420),
.B(n_278),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_424),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_487),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_424),
.B(n_278),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_504),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_481),
.B(n_279),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_487),
.Y(n_574)
);

A2O1A1Ixp33_ASAP7_75t_L g575 ( 
.A1(n_463),
.A2(n_279),
.B(n_280),
.C(n_283),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_484),
.B(n_280),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_484),
.B(n_283),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_491),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_426),
.A2(n_156),
.B1(n_158),
.B2(n_166),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_426),
.B(n_284),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_427),
.B(n_191),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_491),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_524),
.B(n_224),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_530),
.B(n_225),
.Y(n_584)
);

NOR3xp33_ASAP7_75t_L g585 ( 
.A(n_423),
.B(n_227),
.C(n_233),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_473),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_482),
.Y(n_587)
);

A2O1A1Ixp33_ASAP7_75t_L g588 ( 
.A1(n_455),
.A2(n_326),
.B(n_325),
.C(n_323),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_427),
.B(n_250),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_447),
.B(n_326),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_447),
.B(n_241),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_529),
.B(n_254),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_492),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_529),
.B(n_256),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_516),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_429),
.B(n_158),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_528),
.B(n_325),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_470),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_428),
.B(n_261),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_496),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_532),
.B(n_321),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_493),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_496),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_450),
.B(n_168),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_500),
.B(n_321),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_500),
.B(n_320),
.Y(n_606)
);

NOR2xp67_ASAP7_75t_L g607 ( 
.A(n_479),
.B(n_66),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_482),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_467),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_490),
.Y(n_610)
);

BUFx5_ASAP7_75t_L g611 ( 
.A(n_467),
.Y(n_611)
);

CKINVDCx8_ASAP7_75t_R g612 ( 
.A(n_476),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_489),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_450),
.B(n_436),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_526),
.B(n_319),
.Y(n_615)
);

OR2x2_ASAP7_75t_SL g616 ( 
.A(n_462),
.B(n_319),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_526),
.B(n_455),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g618 ( 
.A(n_488),
.B(n_282),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_489),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_476),
.B(n_3),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_464),
.B(n_282),
.Y(n_621)
);

BUFx5_ASAP7_75t_L g622 ( 
.A(n_451),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_464),
.B(n_273),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_518),
.A2(n_273),
.B(n_268),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_502),
.B(n_268),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_502),
.B(n_506),
.Y(n_626)
);

NOR3x1_ASAP7_75t_L g627 ( 
.A(n_531),
.B(n_262),
.C(n_261),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_506),
.B(n_262),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_434),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_515),
.A2(n_259),
.B1(n_258),
.B2(n_257),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_434),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_457),
.A2(n_258),
.B1(n_257),
.B2(n_218),
.Y(n_632)
);

INVx8_ASAP7_75t_L g633 ( 
.A(n_457),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_470),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_436),
.B(n_170),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_458),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_458),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_513),
.B(n_140),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_L g639 ( 
.A(n_537),
.B(n_139),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_513),
.B(n_128),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_441),
.A2(n_117),
.B1(n_105),
.B2(n_103),
.Y(n_641)
);

BUFx5_ASAP7_75t_L g642 ( 
.A(n_459),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_466),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_441),
.B(n_3),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_523),
.B(n_85),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_499),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_452),
.B(n_6),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_520),
.A2(n_79),
.B(n_72),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_431),
.B(n_71),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_431),
.B(n_68),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_432),
.B(n_67),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_432),
.B(n_57),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_515),
.A2(n_471),
.B1(n_446),
.B2(n_519),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_471),
.A2(n_8),
.B1(n_9),
.B2(n_13),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_452),
.B(n_454),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_460),
.B(n_54),
.Y(n_656)
);

INVx8_ASAP7_75t_L g657 ( 
.A(n_470),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_454),
.B(n_15),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_L g659 ( 
.A1(n_425),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_503),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_512),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_512),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_514),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_465),
.B(n_53),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_R g665 ( 
.A(n_498),
.B(n_18),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_419),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_495),
.B(n_21),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_474),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_469),
.B(n_47),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_537),
.B(n_22),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_476),
.B(n_23),
.Y(n_671)
);

AO221x1_ASAP7_75t_L g672 ( 
.A1(n_423),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.C(n_31),
.Y(n_672)
);

AND2x2_ASAP7_75t_SL g673 ( 
.A(n_519),
.B(n_446),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_478),
.B(n_33),
.Y(n_674)
);

NOR3xp33_ASAP7_75t_L g675 ( 
.A(n_486),
.B(n_34),
.C(n_41),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_485),
.B(n_508),
.Y(n_676)
);

AND2x6_ASAP7_75t_SL g677 ( 
.A(n_521),
.B(n_34),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_559),
.Y(n_678)
);

NAND2x1_ASAP7_75t_L g679 ( 
.A(n_629),
.B(n_480),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_626),
.B(n_483),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_556),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_550),
.B(n_477),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_653),
.A2(n_497),
.B1(n_525),
.B2(n_521),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_550),
.B(n_421),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_643),
.A2(n_494),
.B(n_480),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_595),
.B(n_536),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_602),
.B(n_521),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_673),
.A2(n_653),
.B(n_615),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_558),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_602),
.B(n_522),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_613),
.B(n_536),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_564),
.B(n_501),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_614),
.A2(n_655),
.B(n_619),
.Y(n_693)
);

INVx5_ASAP7_75t_L g694 ( 
.A(n_629),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_539),
.A2(n_509),
.B(n_525),
.C(n_517),
.Y(n_695)
);

AOI21x1_ASAP7_75t_L g696 ( 
.A1(n_676),
.A2(n_468),
.B(n_507),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_573),
.B(n_430),
.Y(n_697)
);

AND2x6_ASAP7_75t_SL g698 ( 
.A(n_620),
.B(n_42),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_600),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_590),
.B(n_533),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_631),
.A2(n_535),
.B(n_449),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_597),
.B(n_601),
.Y(n_702)
);

OAI321xp33_ASAP7_75t_L g703 ( 
.A1(n_659),
.A2(n_42),
.A3(n_45),
.B1(n_46),
.B2(n_448),
.C(n_533),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_565),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_631),
.A2(n_442),
.B(n_449),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_596),
.B(n_442),
.Y(n_706)
);

AO21x1_ASAP7_75t_L g707 ( 
.A1(n_638),
.A2(n_448),
.B(n_442),
.Y(n_707)
);

AOI21x1_ASAP7_75t_L g708 ( 
.A1(n_676),
.A2(n_442),
.B(n_449),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_604),
.A2(n_449),
.B(n_535),
.C(n_448),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_640),
.A2(n_448),
.B1(n_535),
.B2(n_645),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_593),
.B(n_562),
.Y(n_711)
);

NOR2xp67_ASAP7_75t_L g712 ( 
.A(n_560),
.B(n_572),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_598),
.B(n_634),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_540),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_551),
.A2(n_589),
.B(n_581),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_551),
.A2(n_603),
.B(n_574),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_570),
.A2(n_578),
.B(n_582),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_592),
.A2(n_594),
.B(n_625),
.C(n_628),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_643),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_563),
.B(n_549),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_540),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_540),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_644),
.A2(n_658),
.B(n_647),
.C(n_580),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_542),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_546),
.B(n_604),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_546),
.B(n_585),
.C(n_579),
.Y(n_726)
);

CKINVDCx10_ASAP7_75t_R g727 ( 
.A(n_556),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_567),
.A2(n_568),
.B(n_571),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_649),
.A2(n_652),
.B(n_651),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_650),
.A2(n_605),
.B(n_606),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_624),
.A2(n_538),
.B(n_623),
.C(n_621),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_545),
.B(n_666),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_646),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_610),
.B(n_671),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_646),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_624),
.A2(n_599),
.B(n_675),
.C(n_584),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_618),
.B(n_654),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_663),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_591),
.A2(n_577),
.B1(n_566),
.B2(n_554),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_639),
.A2(n_656),
.B(n_664),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_667),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_584),
.A2(n_675),
.B(n_654),
.C(n_575),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_637),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_660),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_579),
.A2(n_668),
.B1(n_630),
.B2(n_616),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_611),
.B(n_642),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_544),
.B(n_547),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_630),
.A2(n_659),
.B1(n_641),
.B2(n_632),
.Y(n_748)
);

AO21x1_ASAP7_75t_L g749 ( 
.A1(n_648),
.A2(n_670),
.B(n_669),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_611),
.B(n_622),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_662),
.A2(n_636),
.B(n_661),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_588),
.A2(n_543),
.B(n_674),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_553),
.A2(n_561),
.B(n_557),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_611),
.B(n_622),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_583),
.B(n_585),
.C(n_635),
.Y(n_755)
);

OAI22xp33_ASAP7_75t_L g756 ( 
.A1(n_612),
.A2(n_633),
.B1(n_620),
.B2(n_657),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_611),
.B(n_642),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_611),
.B(n_642),
.Y(n_758)
);

OAI21xp5_ASAP7_75t_L g759 ( 
.A1(n_543),
.A2(n_548),
.B(n_555),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_R g760 ( 
.A(n_541),
.B(n_586),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_552),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_672),
.A2(n_622),
.B1(n_642),
.B2(n_671),
.Y(n_762)
);

BUFx8_ASAP7_75t_SL g763 ( 
.A(n_587),
.Y(n_763)
);

AND2x4_ASAP7_75t_SL g764 ( 
.A(n_620),
.B(n_608),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_622),
.B(n_642),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_622),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_633),
.A2(n_657),
.B(n_642),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_627),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_607),
.B(n_633),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_657),
.B(n_677),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_665),
.Y(n_771)
);

BUFx4f_ASAP7_75t_L g772 ( 
.A(n_665),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_550),
.B(n_602),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_564),
.B(n_598),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_626),
.A2(n_539),
.B(n_655),
.C(n_596),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_595),
.B(n_626),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_626),
.B(n_602),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_556),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_558),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_L g780 ( 
.A(n_573),
.B(n_576),
.C(n_539),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_558),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_602),
.B(n_542),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_542),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_614),
.B(n_461),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_626),
.B(n_602),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_550),
.B(n_602),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_626),
.B(n_602),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_626),
.B(n_602),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_600),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_626),
.B(n_602),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_558),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_617),
.A2(n_673),
.B(n_609),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_558),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_617),
.A2(n_673),
.B(n_609),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_564),
.B(n_598),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_626),
.A2(n_539),
.B(n_655),
.C(n_596),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_569),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_626),
.B(n_602),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_614),
.B(n_461),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_626),
.A2(n_539),
.B(n_655),
.C(n_596),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_550),
.B(n_602),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_550),
.B(n_602),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_542),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_614),
.B(n_461),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_614),
.B(n_461),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_600),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_602),
.B(n_542),
.Y(n_818)
);

OAI21xp33_ASAP7_75t_L g819 ( 
.A1(n_596),
.A2(n_576),
.B(n_573),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_626),
.A2(n_539),
.B(n_655),
.C(n_596),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_552),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_558),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_626),
.B(n_602),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_600),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_552),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_550),
.B(n_602),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_653),
.A2(n_673),
.B1(n_654),
.B2(n_626),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_569),
.A2(n_463),
.B(n_437),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_626),
.B(n_602),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_629),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_819),
.A2(n_780),
.B1(n_725),
.B2(n_726),
.Y(n_835)
);

AOI21xp33_ASAP7_75t_L g836 ( 
.A1(n_742),
.A2(n_748),
.B(n_831),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_693),
.B(n_776),
.Y(n_837)
);

NOR2xp67_ASAP7_75t_L g838 ( 
.A(n_724),
.B(n_812),
.Y(n_838)
);

AOI21xp33_ASAP7_75t_L g839 ( 
.A1(n_748),
.A2(n_831),
.B(n_745),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_693),
.B(n_776),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_775),
.A2(n_802),
.B(n_806),
.C(n_820),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_685),
.A2(n_696),
.B(n_708),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_783),
.B(n_818),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_754),
.A2(n_758),
.B(n_757),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_716),
.A2(n_786),
.B(n_782),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_678),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_773),
.A2(n_808),
.B1(n_809),
.B2(n_830),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_743),
.Y(n_848)
);

OAI21x1_ASAP7_75t_L g849 ( 
.A1(n_795),
.A2(n_799),
.B(n_798),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_744),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_788),
.B(n_777),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_729),
.A2(n_728),
.B(n_715),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_755),
.A2(n_745),
.B1(n_737),
.B2(n_680),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_834),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_800),
.A2(n_810),
.B(n_807),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_811),
.A2(n_817),
.B(n_816),
.Y(n_856)
);

OAI21x1_ASAP7_75t_L g857 ( 
.A1(n_822),
.A2(n_827),
.B(n_823),
.Y(n_857)
);

AO21x1_ASAP7_75t_L g858 ( 
.A1(n_718),
.A2(n_688),
.B(n_794),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_829),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_682),
.B(n_684),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_730),
.A2(n_740),
.B(n_747),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_699),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_791),
.Y(n_863)
);

OAI21x1_ASAP7_75t_L g864 ( 
.A1(n_828),
.A2(n_832),
.B(n_751),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_834),
.Y(n_865)
);

AO31x2_ASAP7_75t_L g866 ( 
.A1(n_749),
.A2(n_707),
.A3(n_731),
.B(n_695),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_834),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_787),
.B(n_789),
.Y(n_868)
);

AO21x1_ASAP7_75t_L g869 ( 
.A1(n_688),
.A2(n_794),
.B(n_797),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_815),
.Y(n_870)
);

OAI21x1_ASAP7_75t_L g871 ( 
.A1(n_717),
.A2(n_701),
.B(n_705),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_790),
.B(n_792),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_679),
.A2(n_686),
.B(n_752),
.Y(n_873)
);

OAI21x1_ASAP7_75t_L g874 ( 
.A1(n_686),
.A2(n_752),
.B(n_766),
.Y(n_874)
);

NAND3xp33_ASAP7_75t_SL g875 ( 
.A(n_739),
.B(n_736),
.C(n_833),
.Y(n_875)
);

AOI21xp33_ASAP7_75t_L g876 ( 
.A1(n_683),
.A2(n_723),
.B(n_785),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_732),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_697),
.A2(n_700),
.B(n_702),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_761),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_735),
.Y(n_880)
);

NAND3xp33_ASAP7_75t_SL g881 ( 
.A(n_804),
.B(n_825),
.C(n_821),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_738),
.Y(n_882)
);

OA22x2_ASAP7_75t_L g883 ( 
.A1(n_741),
.A2(n_784),
.B1(n_768),
.B2(n_734),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_733),
.Y(n_884)
);

OAI22x1_ASAP7_75t_L g885 ( 
.A1(n_687),
.A2(n_734),
.B1(n_711),
.B2(n_770),
.Y(n_885)
);

NAND2xp33_ASAP7_75t_SL g886 ( 
.A(n_714),
.B(n_722),
.Y(n_886)
);

NAND2x1p5_ASAP7_75t_L g887 ( 
.A(n_694),
.B(n_721),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_721),
.B(n_722),
.Y(n_888)
);

OAI22x1_ASAP7_75t_L g889 ( 
.A1(n_770),
.A2(n_813),
.B1(n_814),
.B2(n_805),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_732),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_691),
.B(n_690),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_771),
.B(n_772),
.Y(n_892)
);

O2A1O1Ixp5_ASAP7_75t_L g893 ( 
.A1(n_706),
.A2(n_759),
.B(n_709),
.C(n_720),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_L g894 ( 
.A(n_771),
.B(n_762),
.C(n_774),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_759),
.A2(n_803),
.B(n_767),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_826),
.A2(n_824),
.B(n_689),
.C(n_796),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_704),
.B(n_779),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_704),
.B(n_781),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_713),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_694),
.A2(n_710),
.B(n_793),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_SL g901 ( 
.A1(n_769),
.A2(n_722),
.B(n_714),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_692),
.A2(n_801),
.B(n_774),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_763),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_692),
.B(n_801),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_713),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_703),
.A2(n_712),
.B(n_756),
.Y(n_906)
);

OAI21x1_ASAP7_75t_L g907 ( 
.A1(n_714),
.A2(n_764),
.B(n_760),
.Y(n_907)
);

OAI21x1_ASAP7_75t_SL g908 ( 
.A1(n_698),
.A2(n_727),
.B(n_772),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_681),
.A2(n_778),
.B(n_771),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_693),
.B(n_776),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_693),
.B(n_776),
.Y(n_911)
);

OAI21x1_ASAP7_75t_L g912 ( 
.A1(n_685),
.A2(n_696),
.B(n_708),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_780),
.A2(n_802),
.B(n_775),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_680),
.B(n_773),
.Y(n_914)
);

OAI21x1_ASAP7_75t_SL g915 ( 
.A1(n_767),
.A2(n_723),
.B(n_753),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_831),
.A2(n_653),
.B1(n_802),
.B2(n_775),
.Y(n_916)
);

AO31x2_ASAP7_75t_L g917 ( 
.A1(n_749),
.A2(n_831),
.A3(n_707),
.B(n_802),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_693),
.B(n_776),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_780),
.A2(n_802),
.B(n_775),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_721),
.B(n_714),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_693),
.B(n_776),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_765),
.A2(n_750),
.B(n_746),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_765),
.A2(n_750),
.B(n_746),
.Y(n_923)
);

NAND3xp33_ASAP7_75t_L g924 ( 
.A(n_780),
.B(n_819),
.C(n_576),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_693),
.B(n_776),
.Y(n_925)
);

OAI21x1_ASAP7_75t_L g926 ( 
.A1(n_685),
.A2(n_696),
.B(n_708),
.Y(n_926)
);

OR2x6_ASAP7_75t_L g927 ( 
.A(n_767),
.B(n_657),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_693),
.B(n_776),
.Y(n_928)
);

OAI21x1_ASAP7_75t_L g929 ( 
.A1(n_685),
.A2(n_696),
.B(n_708),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_819),
.A2(n_780),
.B1(n_725),
.B2(n_726),
.Y(n_930)
);

OAI21x1_ASAP7_75t_L g931 ( 
.A1(n_685),
.A2(n_696),
.B(n_708),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_765),
.A2(n_750),
.B(n_746),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_765),
.A2(n_750),
.B(n_746),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_831),
.A2(n_653),
.B1(n_802),
.B2(n_775),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_829),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_693),
.B(n_776),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_719),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_834),
.Y(n_938)
);

AOI221xp5_ASAP7_75t_L g939 ( 
.A1(n_831),
.A2(n_819),
.B1(n_745),
.B2(n_726),
.C(n_748),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_783),
.B(n_818),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_685),
.A2(n_696),
.B(n_708),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_693),
.B(n_776),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_680),
.B(n_417),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_693),
.B(n_776),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_831),
.A2(n_653),
.B1(n_802),
.B2(n_775),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_685),
.A2(n_696),
.B(n_708),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_693),
.B(n_776),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_743),
.Y(n_948)
);

INVx5_ASAP7_75t_L g949 ( 
.A(n_834),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_834),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_734),
.Y(n_951)
);

OR2x6_ASAP7_75t_L g952 ( 
.A(n_767),
.B(n_657),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_765),
.A2(n_750),
.B(n_746),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_743),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_765),
.A2(n_750),
.B(n_746),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_853),
.A2(n_939),
.B(n_839),
.C(n_924),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_860),
.B(n_914),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_859),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_847),
.A2(n_939),
.B1(n_872),
.B2(n_868),
.Y(n_959)
);

NAND3xp33_ASAP7_75t_L g960 ( 
.A(n_835),
.B(n_930),
.C(n_839),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_837),
.B(n_840),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_861),
.A2(n_852),
.B(n_878),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_836),
.A2(n_919),
.B(n_913),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_888),
.B(n_920),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_836),
.A2(n_875),
.B1(n_906),
.B2(n_876),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_935),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_843),
.B(n_940),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_851),
.B(n_868),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_879),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_949),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_848),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_903),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_887),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_837),
.B(n_840),
.Y(n_974)
);

BUFx10_ASAP7_75t_L g975 ( 
.A(n_888),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_943),
.B(n_892),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_872),
.B(n_851),
.Y(n_977)
);

NAND2x1p5_ASAP7_75t_L g978 ( 
.A(n_949),
.B(n_920),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_850),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_862),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_863),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_841),
.A2(n_933),
.B(n_932),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_910),
.B(n_911),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_951),
.B(n_890),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_842),
.A2(n_912),
.B(n_931),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_870),
.Y(n_986)
);

BUFx2_ASAP7_75t_R g987 ( 
.A(n_918),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_918),
.A2(n_928),
.B1(n_925),
.B2(n_921),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_846),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_921),
.B(n_925),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_928),
.B(n_936),
.Y(n_991)
);

OA21x2_ASAP7_75t_L g992 ( 
.A1(n_874),
.A2(n_893),
.B(n_873),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_854),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_899),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_883),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_902),
.B(n_877),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_894),
.A2(n_869),
.B1(n_916),
.B2(n_945),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_904),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_916),
.A2(n_945),
.B(n_934),
.C(n_936),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_934),
.A2(n_955),
.B(n_953),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_854),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_904),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_838),
.B(n_942),
.Y(n_1003)
);

NAND2x1p5_ASAP7_75t_L g1004 ( 
.A(n_949),
.B(n_854),
.Y(n_1004)
);

INVx5_ASAP7_75t_L g1005 ( 
.A(n_950),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_948),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_907),
.B(n_905),
.Y(n_1007)
);

AOI222xp33_ASAP7_75t_L g1008 ( 
.A1(n_942),
.A2(n_944),
.B1(n_947),
.B2(n_881),
.C1(n_885),
.C2(n_889),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_883),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_922),
.A2(n_955),
.B(n_953),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_909),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_947),
.A2(n_891),
.B1(n_954),
.B2(n_923),
.Y(n_1012)
);

AOI222xp33_ASAP7_75t_L g1013 ( 
.A1(n_908),
.A2(n_891),
.B1(n_898),
.B2(n_897),
.C1(n_886),
.C2(n_937),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_923),
.A2(n_895),
.B(n_900),
.C(n_896),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_858),
.B(n_884),
.Y(n_1015)
);

AOI222xp33_ASAP7_75t_L g1016 ( 
.A1(n_898),
.A2(n_882),
.B1(n_880),
.B2(n_915),
.C1(n_865),
.C2(n_867),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_950),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_901),
.B(n_938),
.Y(n_1018)
);

OR2x2_ASAP7_75t_SL g1019 ( 
.A(n_927),
.B(n_952),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_917),
.B(n_844),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_927),
.B(n_952),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_927),
.B(n_952),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_849),
.B(n_855),
.Y(n_1023)
);

AND2x6_ASAP7_75t_L g1024 ( 
.A(n_917),
.B(n_866),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_900),
.B(n_864),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_917),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_866),
.B(n_856),
.Y(n_1027)
);

BUFx12f_ASAP7_75t_L g1028 ( 
.A(n_857),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_845),
.Y(n_1029)
);

BUFx10_ASAP7_75t_L g1030 ( 
.A(n_871),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_926),
.A2(n_929),
.B(n_941),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_946),
.B(n_860),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_860),
.B(n_783),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_860),
.A2(n_819),
.B1(n_780),
.B2(n_725),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_L g1035 ( 
.A(n_939),
.B(n_780),
.C(n_819),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_SL g1036 ( 
.A(n_859),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_839),
.A2(n_819),
.B(n_775),
.C(n_806),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_836),
.A2(n_780),
.B(n_839),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_847),
.B(n_837),
.Y(n_1039)
);

INVx3_ASAP7_75t_SL g1040 ( 
.A(n_903),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_888),
.B(n_920),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_879),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_847),
.B(n_837),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_861),
.A2(n_852),
.B(n_878),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_847),
.B(n_837),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_847),
.B(n_837),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_847),
.B(n_837),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_860),
.B(n_783),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_939),
.A2(n_819),
.B1(n_780),
.B2(n_726),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_859),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_887),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_847),
.B(n_837),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_939),
.A2(n_819),
.B1(n_780),
.B2(n_726),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_861),
.A2(n_852),
.B(n_878),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_847),
.A2(n_831),
.B1(n_653),
.B2(n_776),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_887),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_879),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_860),
.B(n_783),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_854),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_860),
.B(n_783),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_860),
.B(n_914),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_862),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_839),
.A2(n_819),
.B(n_775),
.C(n_806),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_879),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_853),
.A2(n_819),
.B(n_780),
.C(n_802),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_847),
.B(n_837),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_847),
.B(n_837),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_860),
.B(n_783),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_853),
.A2(n_819),
.B(n_780),
.C(n_802),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_860),
.B(n_783),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_862),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_887),
.Y(n_1072)
);

NAND2x1p5_ASAP7_75t_L g1073 ( 
.A(n_949),
.B(n_888),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_981),
.Y(n_1074)
);

BUFx8_ASAP7_75t_L g1075 ( 
.A(n_1036),
.Y(n_1075)
);

CKINVDCx11_ASAP7_75t_R g1076 ( 
.A(n_972),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_958),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_986),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1006),
.Y(n_1079)
);

OAI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_1034),
.A2(n_1035),
.B1(n_977),
.B2(n_960),
.Y(n_1080)
);

OR2x6_ASAP7_75t_L g1081 ( 
.A(n_1022),
.B(n_1021),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_957),
.B(n_1061),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_967),
.B(n_976),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1062),
.Y(n_1084)
);

BUFx2_ASAP7_75t_R g1085 ( 
.A(n_1040),
.Y(n_1085)
);

NAND2x1p5_ASAP7_75t_L g1086 ( 
.A(n_1022),
.B(n_970),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1071),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_971),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1033),
.B(n_1048),
.Y(n_1089)
);

INVxp67_ASAP7_75t_SL g1090 ( 
.A(n_969),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_979),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1058),
.B(n_1060),
.Y(n_1092)
);

INVx6_ASAP7_75t_L g1093 ( 
.A(n_975),
.Y(n_1093)
);

OA21x2_ASAP7_75t_L g1094 ( 
.A1(n_962),
.A2(n_1044),
.B(n_1054),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_1005),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_966),
.Y(n_1096)
);

INVxp33_ASAP7_75t_L g1097 ( 
.A(n_984),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_968),
.B(n_1039),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_998),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_1007),
.B(n_964),
.Y(n_1100)
);

BUFx10_ASAP7_75t_L g1101 ( 
.A(n_1036),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_1005),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_1050),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1068),
.B(n_1070),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_SL g1105 ( 
.A1(n_1038),
.A2(n_959),
.B1(n_1055),
.B2(n_995),
.Y(n_1105)
);

BUFx12f_ASAP7_75t_L g1106 ( 
.A(n_1042),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1015),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_1057),
.Y(n_1108)
);

CKINVDCx11_ASAP7_75t_R g1109 ( 
.A(n_975),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1015),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_1064),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1049),
.A2(n_1053),
.B1(n_965),
.B2(n_1038),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_989),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_SL g1114 ( 
.A1(n_959),
.A2(n_1055),
.B1(n_963),
.B2(n_1009),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1007),
.B(n_964),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1041),
.B(n_996),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_992),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1002),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_SL g1119 ( 
.A1(n_987),
.A2(n_1046),
.B1(n_1067),
.B2(n_1066),
.Y(n_1119)
);

OAI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1043),
.A2(n_1052),
.B1(n_1066),
.B2(n_1067),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1002),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_992),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1045),
.A2(n_1052),
.B1(n_1047),
.B2(n_1046),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1041),
.B(n_1003),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1027),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1065),
.A2(n_1069),
.B(n_956),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_1019),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_994),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1012),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1012),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1026),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1045),
.A2(n_1047),
.B1(n_997),
.B2(n_1008),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_961),
.B(n_991),
.Y(n_1133)
);

BUFx10_ASAP7_75t_L g1134 ( 
.A(n_1018),
.Y(n_1134)
);

CKINVDCx8_ASAP7_75t_R g1135 ( 
.A(n_993),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_993),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_SL g1137 ( 
.A1(n_1000),
.A2(n_988),
.B1(n_982),
.B2(n_1032),
.Y(n_1137)
);

CKINVDCx11_ASAP7_75t_R g1138 ( 
.A(n_1001),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_SL g1139 ( 
.A1(n_988),
.A2(n_1011),
.B1(n_983),
.B2(n_974),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1008),
.A2(n_1013),
.B1(n_990),
.B2(n_974),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1025),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1001),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1025),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1029),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1020),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1013),
.A2(n_991),
.B1(n_1024),
.B2(n_1016),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1023),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1017),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_973),
.B(n_1056),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1017),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_978),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1073),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1004),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1004),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_999),
.B(n_1063),
.Y(n_1155)
);

CKINVDCx11_ASAP7_75t_R g1156 ( 
.A(n_1028),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_1059),
.Y(n_1157)
);

AO21x1_ASAP7_75t_L g1158 ( 
.A1(n_1037),
.A2(n_1010),
.B(n_1073),
.Y(n_1158)
);

BUFx12f_ASAP7_75t_L g1159 ( 
.A(n_1059),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1014),
.A2(n_1051),
.B1(n_1072),
.B2(n_1016),
.Y(n_1160)
);

OR2x6_ASAP7_75t_L g1161 ( 
.A(n_1072),
.B(n_1024),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_1030),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1030),
.A2(n_1031),
.B(n_985),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1024),
.Y(n_1164)
);

OAI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1034),
.A2(n_847),
.B1(n_726),
.B2(n_831),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_980),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1131),
.Y(n_1167)
);

AO21x1_ASAP7_75t_L g1168 ( 
.A1(n_1126),
.A2(n_1080),
.B(n_1165),
.Y(n_1168)
);

AO31x2_ASAP7_75t_L g1169 ( 
.A1(n_1158),
.A2(n_1122),
.A3(n_1117),
.B(n_1129),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1098),
.B(n_1082),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1145),
.B(n_1130),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1125),
.B(n_1114),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1105),
.B(n_1130),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1134),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1110),
.B(n_1123),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1144),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1144),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1141),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1081),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1110),
.B(n_1123),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1118),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_1081),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1094),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1164),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1143),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1143),
.Y(n_1186)
);

OR2x6_ASAP7_75t_L g1187 ( 
.A(n_1161),
.B(n_1147),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1107),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1121),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1134),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1094),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1081),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_1155),
.B(n_1120),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1137),
.B(n_1098),
.Y(n_1194)
);

BUFx5_ASAP7_75t_L g1195 ( 
.A(n_1134),
.Y(n_1195)
);

OA21x2_ASAP7_75t_L g1196 ( 
.A1(n_1146),
.A2(n_1163),
.B(n_1140),
.Y(n_1196)
);

AO21x2_ASAP7_75t_L g1197 ( 
.A1(n_1165),
.A2(n_1160),
.B(n_1120),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_1093),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1088),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1091),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1099),
.B(n_1080),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1161),
.B(n_1100),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1166),
.B(n_1083),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1082),
.B(n_1133),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1090),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1112),
.A2(n_1132),
.B(n_1140),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1108),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1108),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1074),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1078),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1162),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1115),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1079),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1084),
.Y(n_1214)
);

NAND2x1p5_ASAP7_75t_L g1215 ( 
.A(n_1115),
.B(n_1124),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1087),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1093),
.Y(n_1217)
);

OR2x6_ASAP7_75t_L g1218 ( 
.A(n_1086),
.B(n_1115),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1146),
.A2(n_1132),
.B(n_1112),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_1111),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1089),
.B(n_1092),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1139),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1104),
.B(n_1097),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1111),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1149),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1149),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1116),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1153),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1154),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1175),
.B(n_1119),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1169),
.B(n_1127),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1169),
.Y(n_1232)
);

OAI211xp5_ASAP7_75t_L g1233 ( 
.A1(n_1206),
.A2(n_1170),
.B(n_1194),
.C(n_1219),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1169),
.B(n_1127),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1169),
.B(n_1150),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1183),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1169),
.B(n_1148),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1169),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1194),
.B(n_1156),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1176),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1176),
.Y(n_1241)
);

INVxp67_ASAP7_75t_SL g1242 ( 
.A(n_1205),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1177),
.Y(n_1243)
);

AND2x6_ASAP7_75t_SL g1244 ( 
.A(n_1218),
.B(n_1085),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1168),
.A2(n_1106),
.B1(n_1152),
.B2(n_1151),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1191),
.B(n_1142),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1197),
.B(n_1113),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1201),
.B(n_1157),
.Y(n_1248)
);

INVx2_ASAP7_75t_R g1249 ( 
.A(n_1167),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1177),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1197),
.B(n_1136),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1197),
.B(n_1101),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1168),
.A2(n_1106),
.B1(n_1076),
.B2(n_1075),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1178),
.B(n_1101),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1180),
.B(n_1193),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1195),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1219),
.A2(n_1076),
.B1(n_1075),
.B2(n_1109),
.Y(n_1257)
);

NOR3xp33_ASAP7_75t_L g1258 ( 
.A(n_1222),
.B(n_1109),
.C(n_1128),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1187),
.Y(n_1259)
);

AOI21xp33_ASAP7_75t_L g1260 ( 
.A1(n_1219),
.A2(n_1075),
.B(n_1159),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1255),
.B(n_1242),
.Y(n_1261)
);

OAI211xp5_ASAP7_75t_L g1262 ( 
.A1(n_1233),
.A2(n_1222),
.B(n_1204),
.C(n_1193),
.Y(n_1262)
);

OAI221xp5_ASAP7_75t_L g1263 ( 
.A1(n_1253),
.A2(n_1224),
.B1(n_1223),
.B2(n_1220),
.C(n_1179),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1233),
.A2(n_1173),
.B(n_1196),
.Y(n_1264)
);

AND2x2_ASAP7_75t_SL g1265 ( 
.A(n_1231),
.B(n_1196),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1258),
.A2(n_1173),
.B1(n_1227),
.B2(n_1224),
.Y(n_1266)
);

NOR3xp33_ASAP7_75t_L g1267 ( 
.A(n_1260),
.B(n_1179),
.C(n_1192),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1255),
.B(n_1181),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1255),
.B(n_1189),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1242),
.B(n_1223),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1247),
.B(n_1171),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1247),
.B(n_1171),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1253),
.A2(n_1196),
.B1(n_1208),
.B2(n_1207),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1247),
.B(n_1188),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1247),
.B(n_1172),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1231),
.B(n_1185),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1230),
.A2(n_1196),
.B1(n_1172),
.B2(n_1221),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1258),
.B(n_1174),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1234),
.B(n_1185),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1257),
.A2(n_1227),
.B1(n_1192),
.B2(n_1182),
.Y(n_1280)
);

NAND3xp33_ASAP7_75t_L g1281 ( 
.A(n_1257),
.B(n_1229),
.C(n_1228),
.Y(n_1281)
);

AND2x2_ASAP7_75t_SL g1282 ( 
.A(n_1234),
.B(n_1202),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1234),
.B(n_1186),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1234),
.B(n_1186),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1230),
.A2(n_1221),
.B1(n_1188),
.B2(n_1203),
.Y(n_1285)
);

OAI221xp5_ASAP7_75t_SL g1286 ( 
.A1(n_1245),
.A2(n_1187),
.B1(n_1218),
.B2(n_1226),
.C(n_1225),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1246),
.B(n_1184),
.Y(n_1287)
);

NAND3xp33_ASAP7_75t_L g1288 ( 
.A(n_1245),
.B(n_1229),
.C(n_1228),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1240),
.B(n_1199),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1239),
.B(n_1198),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1239),
.A2(n_1182),
.B1(n_1202),
.B2(n_1212),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1245),
.A2(n_1202),
.B(n_1215),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1240),
.B(n_1199),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1241),
.B(n_1200),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1241),
.B(n_1243),
.Y(n_1295)
);

OR2x2_ASAP7_75t_SL g1296 ( 
.A(n_1248),
.B(n_1211),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1236),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1243),
.B(n_1200),
.Y(n_1298)
);

AOI221xp5_ASAP7_75t_L g1299 ( 
.A1(n_1252),
.A2(n_1209),
.B1(n_1210),
.B2(n_1213),
.C(n_1214),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1250),
.B(n_1252),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1246),
.B(n_1184),
.Y(n_1301)
);

NAND3xp33_ASAP7_75t_L g1302 ( 
.A(n_1252),
.B(n_1210),
.C(n_1216),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1297),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1297),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1261),
.B(n_1235),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1274),
.B(n_1232),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1289),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1265),
.B(n_1249),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1302),
.B(n_1256),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1293),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1268),
.B(n_1237),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1265),
.B(n_1249),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1300),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1296),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1265),
.B(n_1249),
.Y(n_1315)
);

INVxp67_ASAP7_75t_L g1316 ( 
.A(n_1302),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1267),
.B(n_1256),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1296),
.B(n_1232),
.Y(n_1318)
);

OR2x6_ASAP7_75t_L g1319 ( 
.A(n_1292),
.B(n_1259),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1295),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1276),
.B(n_1256),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1276),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1294),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1282),
.B(n_1238),
.Y(n_1324)
);

NOR2xp67_ASAP7_75t_L g1325 ( 
.A(n_1288),
.B(n_1252),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1298),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1271),
.B(n_1250),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1282),
.B(n_1237),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1269),
.B(n_1237),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1282),
.B(n_1279),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1271),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1283),
.B(n_1237),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1272),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1307),
.B(n_1275),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1319),
.B(n_1288),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1330),
.B(n_1283),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1307),
.B(n_1285),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1310),
.B(n_1285),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1327),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1310),
.B(n_1270),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1327),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1303),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1323),
.B(n_1326),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1306),
.B(n_1272),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1327),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1322),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1330),
.B(n_1284),
.Y(n_1347)
);

NAND2x1_ASAP7_75t_L g1348 ( 
.A(n_1319),
.B(n_1259),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1319),
.B(n_1284),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1319),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1319),
.B(n_1254),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1323),
.B(n_1251),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1320),
.Y(n_1353)
);

AOI32xp33_ASAP7_75t_L g1354 ( 
.A1(n_1308),
.A2(n_1273),
.A3(n_1277),
.B1(n_1278),
.B2(n_1263),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1330),
.B(n_1292),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1322),
.Y(n_1356)
);

INVxp67_ASAP7_75t_SL g1357 ( 
.A(n_1325),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1320),
.Y(n_1358)
);

NAND2x1p5_ASAP7_75t_L g1359 ( 
.A(n_1325),
.B(n_1256),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1306),
.B(n_1277),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1303),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_L g1362 ( 
.A(n_1316),
.B(n_1262),
.C(n_1273),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1328),
.B(n_1287),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1328),
.B(n_1301),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1303),
.Y(n_1365)
);

NOR2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1314),
.B(n_1281),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1304),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1328),
.B(n_1301),
.Y(n_1368)
);

INVxp33_ASAP7_75t_SL g1369 ( 
.A(n_1324),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1304),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1355),
.B(n_1314),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1353),
.Y(n_1372)
);

OAI221xp5_ASAP7_75t_L g1373 ( 
.A1(n_1354),
.A2(n_1316),
.B1(n_1266),
.B2(n_1314),
.C(n_1291),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1337),
.B(n_1311),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1350),
.B(n_1319),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1338),
.B(n_1311),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1355),
.B(n_1336),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1362),
.B(n_1313),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1357),
.B(n_1308),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1358),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1339),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1369),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1369),
.B(n_1290),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1339),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1366),
.B(n_1313),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1340),
.B(n_1329),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1341),
.B(n_1329),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1349),
.B(n_1308),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1350),
.B(n_1309),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1345),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1348),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1334),
.B(n_1345),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1343),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1360),
.B(n_1305),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1361),
.Y(n_1395)
);

OAI31xp33_ASAP7_75t_L g1396 ( 
.A1(n_1335),
.A2(n_1315),
.A3(n_1312),
.B(n_1317),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1335),
.A2(n_1264),
.B1(n_1281),
.B2(n_1317),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1370),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1363),
.B(n_1331),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1349),
.B(n_1312),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1361),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1360),
.B(n_1305),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1365),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1349),
.B(n_1312),
.Y(n_1404)
);

OAI21xp33_ASAP7_75t_L g1405 ( 
.A1(n_1335),
.A2(n_1264),
.B(n_1315),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1365),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_SL g1407 ( 
.A(n_1350),
.B(n_1286),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1336),
.B(n_1321),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1363),
.B(n_1331),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1344),
.B(n_1333),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1342),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1344),
.B(n_1333),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1382),
.B(n_1364),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1378),
.B(n_1364),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1377),
.B(n_1359),
.Y(n_1415)
);

NOR3xp33_ASAP7_75t_L g1416 ( 
.A(n_1373),
.B(n_1260),
.C(n_1348),
.Y(n_1416)
);

NAND3xp33_ASAP7_75t_L g1417 ( 
.A(n_1407),
.B(n_1315),
.C(n_1299),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1385),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1381),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1371),
.B(n_1375),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1371),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1383),
.B(n_1368),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1375),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1395),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1394),
.B(n_1352),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1383),
.B(n_1372),
.Y(n_1426)
);

NOR2x1_ASAP7_75t_L g1427 ( 
.A(n_1391),
.B(n_1318),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1397),
.B(n_1359),
.Y(n_1428)
);

CKINVDCx16_ASAP7_75t_R g1429 ( 
.A(n_1375),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1384),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1390),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1401),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1389),
.B(n_1359),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1403),
.Y(n_1434)
);

NAND3x1_ASAP7_75t_L g1435 ( 
.A(n_1396),
.B(n_1324),
.C(n_1347),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1380),
.B(n_1368),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1386),
.B(n_1347),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1406),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1389),
.B(n_1351),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1411),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1389),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1379),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1379),
.B(n_1351),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1408),
.B(n_1351),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1388),
.B(n_1332),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1391),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1388),
.B(n_1332),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1421),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1441),
.Y(n_1449)
);

OAI32xp33_ASAP7_75t_L g1450 ( 
.A1(n_1418),
.A2(n_1405),
.A3(n_1318),
.B1(n_1374),
.B2(n_1376),
.Y(n_1450)
);

NOR2x1_ASAP7_75t_L g1451 ( 
.A(n_1423),
.B(n_1391),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1418),
.B(n_1386),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1424),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1428),
.A2(n_1392),
.B(n_1393),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1442),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1420),
.B(n_1400),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1426),
.B(n_1402),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1432),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1422),
.B(n_1399),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1423),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1432),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1434),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1441),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1424),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1434),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1420),
.B(n_1400),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1442),
.B(n_1404),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1433),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1438),
.Y(n_1469)
);

AOI21xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1429),
.A2(n_1387),
.B(n_1096),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1438),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1419),
.Y(n_1472)
);

NAND2x1_ASAP7_75t_L g1473 ( 
.A(n_1451),
.B(n_1427),
.Y(n_1473)
);

NOR3xp33_ASAP7_75t_L g1474 ( 
.A(n_1449),
.B(n_1429),
.C(n_1417),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1455),
.Y(n_1475)
);

INVxp67_ASAP7_75t_L g1476 ( 
.A(n_1460),
.Y(n_1476)
);

NAND2x1_ASAP7_75t_L g1477 ( 
.A(n_1467),
.B(n_1427),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1463),
.B(n_1413),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1452),
.B(n_1414),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1460),
.B(n_1442),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1453),
.Y(n_1481)
);

INVxp67_ASAP7_75t_L g1482 ( 
.A(n_1448),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1453),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_SL g1484 ( 
.A(n_1470),
.B(n_1417),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1456),
.B(n_1439),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1448),
.B(n_1437),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1468),
.B(n_1436),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1468),
.B(n_1445),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1457),
.B(n_1439),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1456),
.B(n_1443),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1464),
.Y(n_1491)
);

NOR3xp33_ASAP7_75t_L g1492 ( 
.A(n_1474),
.B(n_1450),
.C(n_1458),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1473),
.A2(n_1477),
.B(n_1484),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1479),
.A2(n_1450),
.B(n_1454),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1476),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1478),
.A2(n_1459),
.B(n_1416),
.Y(n_1496)
);

AOI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1482),
.A2(n_1472),
.B1(n_1471),
.B2(n_1469),
.C(n_1461),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1482),
.A2(n_1446),
.B(n_1467),
.Y(n_1498)
);

OAI221xp5_ASAP7_75t_L g1499 ( 
.A1(n_1489),
.A2(n_1446),
.B1(n_1465),
.B2(n_1462),
.C(n_1466),
.Y(n_1499)
);

OAI21xp5_ASAP7_75t_SL g1500 ( 
.A1(n_1486),
.A2(n_1466),
.B(n_1467),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1476),
.A2(n_1464),
.B(n_1430),
.Y(n_1501)
);

O2A1O1Ixp5_ASAP7_75t_L g1502 ( 
.A1(n_1475),
.A2(n_1433),
.B(n_1424),
.C(n_1440),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1498),
.B(n_1490),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1495),
.B(n_1103),
.Y(n_1504)
);

OAI322xp33_ASAP7_75t_L g1505 ( 
.A1(n_1494),
.A2(n_1480),
.A3(n_1487),
.B1(n_1488),
.B2(n_1481),
.C1(n_1483),
.C2(n_1491),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1493),
.B(n_1485),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1501),
.Y(n_1507)
);

AOI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1492),
.A2(n_1430),
.B1(n_1431),
.B2(n_1419),
.C(n_1440),
.Y(n_1508)
);

NOR3xp33_ASAP7_75t_L g1509 ( 
.A(n_1499),
.B(n_1431),
.C(n_1077),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1502),
.Y(n_1510)
);

NAND4xp25_ASAP7_75t_SL g1511 ( 
.A(n_1496),
.B(n_1415),
.C(n_1443),
.D(n_1435),
.Y(n_1511)
);

O2A1O1Ixp5_ASAP7_75t_L g1512 ( 
.A1(n_1510),
.A2(n_1415),
.B(n_1500),
.C(n_1497),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_SL g1513 ( 
.A(n_1503),
.B(n_1435),
.C(n_1135),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1506),
.B(n_1444),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1507),
.B(n_1445),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1508),
.B(n_1447),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1513),
.A2(n_1511),
.B1(n_1509),
.B2(n_1504),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1515),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1516),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1514),
.A2(n_1444),
.B1(n_1447),
.B2(n_1404),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1512),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1515),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1521),
.B(n_1505),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_L g1524 ( 
.A(n_1518),
.B(n_1103),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1519),
.B(n_1425),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1522),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1517),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1525),
.B(n_1520),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1524),
.B(n_1523),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1527),
.A2(n_1425),
.B1(n_1317),
.B2(n_1174),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1528),
.Y(n_1531)
);

AOI222xp33_ASAP7_75t_L g1532 ( 
.A1(n_1531),
.A2(n_1529),
.B1(n_1526),
.B2(n_1530),
.C1(n_1398),
.C2(n_1409),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1532),
.A2(n_1398),
.B1(n_1317),
.B2(n_1190),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1533),
.A2(n_1138),
.B1(n_1317),
.B2(n_1198),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1534),
.A2(n_1412),
.B1(n_1410),
.B2(n_1346),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1535),
.A2(n_1370),
.B(n_1342),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1536),
.A2(n_1138),
.B1(n_1159),
.B2(n_1217),
.Y(n_1537)
);

OAI221xp5_ASAP7_75t_R g1538 ( 
.A1(n_1536),
.A2(n_1280),
.B1(n_1244),
.B2(n_1217),
.C(n_1367),
.Y(n_1538)
);

OAI221xp5_ASAP7_75t_R g1539 ( 
.A1(n_1537),
.A2(n_1244),
.B1(n_1356),
.B2(n_1346),
.C(n_1318),
.Y(n_1539)
);

AOI211xp5_ASAP7_75t_L g1540 ( 
.A1(n_1539),
.A2(n_1538),
.B(n_1095),
.C(n_1102),
.Y(n_1540)
);


endmodule