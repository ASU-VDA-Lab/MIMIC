module fake_netlist_6_3421_n_1770 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1770);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1770;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g174 ( 
.A(n_49),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_11),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_83),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_11),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_25),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_100),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_110),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_173),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_35),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_74),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_40),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_6),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_65),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_9),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_73),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_151),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_95),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_52),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_75),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_21),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_133),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_165),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_118),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_94),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_62),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_116),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_124),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_120),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_15),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_86),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_36),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_111),
.Y(n_212)
);

BUFx8_ASAP7_75t_SL g213 ( 
.A(n_171),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_2),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_33),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_54),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_14),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_168),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_82),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_127),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_59),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_7),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_15),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_64),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_50),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_122),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_76),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_49),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_45),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_48),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_32),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_67),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_125),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_0),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_88),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_42),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_108),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_138),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_163),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_147),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_105),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_155),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_54),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_109),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_129),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_167),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_2),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_101),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_140),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_31),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_141),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_42),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_121),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_164),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_66),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_4),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_166),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_80),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_10),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_91),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_106),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_17),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_14),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_40),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_21),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_135),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_56),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_58),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_99),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_19),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_35),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_63),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_104),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_136),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_37),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_37),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_47),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_10),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_160),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_154),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_117),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_20),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_7),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_46),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_38),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_68),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_32),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_29),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_5),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_34),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_8),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_96),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_169),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_162),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_69),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_170),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_33),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_8),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_12),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_70),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_150),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_27),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_128),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_58),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_9),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_158),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_1),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_153),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_43),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_51),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_103),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_28),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_93),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_77),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_3),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_34),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_46),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_134),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_172),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_148),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_29),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_72),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_102),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_6),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_152),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_45),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_22),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_92),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_18),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_44),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_30),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_85),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_38),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_20),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_131),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_145),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_149),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_98),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_139),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_25),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_52),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_5),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_81),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_3),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_115),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_17),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_87),
.Y(n_348)
);

BUFx10_ASAP7_75t_L g349 ( 
.A(n_84),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_71),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_19),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_114),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_107),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_328),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_174),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_263),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_222),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_221),
.B(n_0),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_261),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_235),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_176),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_235),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_263),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_300),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_312),
.B(n_1),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_263),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_177),
.B(n_4),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_226),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_263),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_229),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_302),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_333),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_213),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_263),
.Y(n_374)
);

BUFx6f_ASAP7_75t_SL g375 ( 
.A(n_202),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_259),
.B(n_12),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_232),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_348),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_253),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_265),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_268),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_248),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_178),
.Y(n_383)
);

INVxp33_ASAP7_75t_L g384 ( 
.A(n_185),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_209),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_211),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_214),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_223),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_297),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_309),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_269),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_309),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_248),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_186),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_199),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_272),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_230),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_231),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_220),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_244),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_251),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_271),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_284),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_272),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_260),
.Y(n_406)
);

INVxp33_ASAP7_75t_SL g407 ( 
.A(n_186),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_190),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_277),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_228),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_283),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_236),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_286),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_325),
.B(n_13),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_R g415 ( 
.A(n_239),
.B(n_161),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_334),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_285),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_240),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_202),
.Y(n_419)
);

BUFx2_ASAP7_75t_SL g420 ( 
.A(n_259),
.Y(n_420)
);

INVxp33_ASAP7_75t_L g421 ( 
.A(n_341),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_288),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_242),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_179),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_181),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_243),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_184),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_245),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_187),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_188),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_289),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_247),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_290),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_279),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_279),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_193),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_195),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_249),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_291),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_197),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_292),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_219),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_190),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_305),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_305),
.Y(n_445)
);

NOR2xp67_ASAP7_75t_L g446 ( 
.A(n_276),
.B(n_13),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_254),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_356),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_363),
.B(n_321),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_356),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_374),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_395),
.Y(n_454)
);

OA21x2_ASAP7_75t_L g455 ( 
.A1(n_366),
.A2(n_203),
.B(n_191),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_369),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_394),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_358),
.B(n_202),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_394),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_397),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_427),
.B(n_321),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_397),
.Y(n_462)
);

INVxp33_ASAP7_75t_SL g463 ( 
.A(n_354),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_382),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_424),
.B(n_344),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_382),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_405),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_405),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_425),
.B(n_344),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_376),
.B(n_294),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_443),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_434),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_365),
.B(n_294),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_434),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_435),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_435),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_385),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_SL g478 ( 
.A(n_375),
.B(n_237),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_444),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_420),
.B(n_252),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_444),
.Y(n_481)
);

AND2x6_ASAP7_75t_L g482 ( 
.A(n_429),
.B(n_294),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_430),
.B(n_436),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_445),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_419),
.B(n_233),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_437),
.B(n_180),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_445),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_440),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_442),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_383),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_386),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_387),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_388),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_373),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_390),
.B(n_180),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_391),
.B(n_182),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_393),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_420),
.B(n_182),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_389),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_360),
.B(n_189),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_400),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_398),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_399),
.Y(n_504)
);

OA21x2_ASAP7_75t_L g505 ( 
.A1(n_401),
.A2(n_203),
.B(n_191),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_402),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_362),
.B(n_189),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_406),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_413),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_372),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_354),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_416),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_364),
.Y(n_514)
);

OA21x2_ASAP7_75t_L g515 ( 
.A1(n_355),
.A2(n_352),
.B(n_205),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_396),
.B(n_237),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_367),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_357),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_357),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_367),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_414),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_414),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_411),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_446),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_384),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_492),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_477),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_520),
.A2(n_361),
.B1(n_410),
.B2(n_428),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_456),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_525),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_458),
.B(n_205),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_450),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_456),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_492),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_477),
.B(n_224),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_491),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_470),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_491),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_477),
.B(n_225),
.Y(n_539)
);

OR2x6_ASAP7_75t_L g540 ( 
.A(n_520),
.B(n_266),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_456),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_449),
.B(n_227),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_473),
.A2(n_521),
.B1(n_522),
.B2(n_520),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_458),
.B(n_352),
.Y(n_544)
);

AND2x6_ASAP7_75t_L g545 ( 
.A(n_521),
.B(n_294),
.Y(n_545)
);

NAND2x1p5_ASAP7_75t_L g546 ( 
.A(n_483),
.B(n_234),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_449),
.B(n_238),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_449),
.B(n_241),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_483),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_450),
.Y(n_550)
);

AO22x2_ASAP7_75t_L g551 ( 
.A1(n_486),
.A2(n_266),
.B1(n_198),
.B2(n_216),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_493),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_525),
.B(n_421),
.Y(n_553)
);

BUFx4f_ASAP7_75t_L g554 ( 
.A(n_473),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_504),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_506),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_521),
.B(n_368),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_506),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_522),
.B(n_368),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_522),
.B(n_370),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_460),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_508),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_449),
.B(n_250),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_473),
.A2(n_516),
.B1(n_461),
.B2(n_470),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_523),
.B(n_370),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_483),
.Y(n_566)
);

INVx3_ASAP7_75t_R g567 ( 
.A(n_512),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_449),
.B(n_255),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_523),
.B(n_377),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_508),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_509),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_480),
.B(n_294),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_498),
.B(n_407),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_509),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_510),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_483),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_523),
.B(n_377),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_475),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_498),
.B(n_407),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_460),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_492),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_492),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_511),
.A2(n_447),
.B1(n_412),
.B2(n_418),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_480),
.B(n_378),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_499),
.B(n_379),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_473),
.A2(n_408),
.B1(n_375),
.B2(n_281),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_510),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_473),
.A2(n_408),
.B1(n_375),
.B2(n_273),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_492),
.Y(n_589)
);

CKINVDCx8_ASAP7_75t_R g590 ( 
.A(n_502),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_499),
.B(n_379),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_511),
.B(n_423),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_514),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_514),
.Y(n_594)
);

AND2x6_ASAP7_75t_L g595 ( 
.A(n_517),
.B(n_262),
.Y(n_595)
);

AND2x6_ASAP7_75t_L g596 ( 
.A(n_517),
.B(n_267),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_471),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_483),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_496),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_483),
.Y(n_600)
);

BUFx4_ASAP7_75t_L g601 ( 
.A(n_496),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_454),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_463),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_448),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_454),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_451),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_497),
.B(n_426),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_473),
.B(n_380),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_497),
.B(n_380),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_483),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_483),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_492),
.Y(n_612)
);

AND2x2_ASAP7_75t_SL g613 ( 
.A(n_518),
.B(n_293),
.Y(n_613)
);

AND2x2_ASAP7_75t_SL g614 ( 
.A(n_518),
.B(n_304),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_494),
.B(n_323),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_512),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_452),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_475),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_452),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_461),
.B(n_381),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_453),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_515),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_515),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_513),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_494),
.B(n_336),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_471),
.B(n_432),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_519),
.B(n_438),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_524),
.B(n_392),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_519),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_475),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_487),
.B(n_403),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_475),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_501),
.B(n_403),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_473),
.B(n_404),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_501),
.Y(n_635)
);

AO22x2_ASAP7_75t_L g636 ( 
.A1(n_486),
.A2(n_257),
.B1(n_346),
.B2(n_340),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_475),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_475),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_513),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_507),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_513),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_513),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_505),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_516),
.B(n_404),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_494),
.B(n_353),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_507),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_487),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_495),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_L g649 ( 
.A(n_473),
.B(n_417),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_468),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_468),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_489),
.B(n_417),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_489),
.B(n_422),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_489),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_515),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_468),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_490),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_470),
.B(n_422),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_527),
.B(n_500),
.Y(n_659)
);

BUFx6f_ASAP7_75t_SL g660 ( 
.A(n_613),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_599),
.A2(n_470),
.B1(n_515),
.B2(n_175),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_536),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_538),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_527),
.B(n_500),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_599),
.A2(n_470),
.B1(n_515),
.B2(n_183),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_643),
.B(n_505),
.Y(n_666)
);

OAI221xp5_ASAP7_75t_L g667 ( 
.A1(n_640),
.A2(n_465),
.B1(n_469),
.B2(n_484),
.C(n_503),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_552),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_635),
.B(n_431),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_646),
.B(n_431),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_555),
.Y(n_671)
);

NOR2xp67_ASAP7_75t_L g672 ( 
.A(n_583),
.B(n_433),
.Y(n_672)
);

OR2x6_ASAP7_75t_L g673 ( 
.A(n_616),
.B(n_484),
.Y(n_673)
);

AO22x2_ASAP7_75t_L g674 ( 
.A1(n_644),
.A2(n_469),
.B1(n_465),
.B2(n_264),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_553),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_556),
.Y(n_676)
);

OAI221xp5_ASAP7_75t_L g677 ( 
.A1(n_640),
.A2(n_503),
.B1(n_490),
.B2(n_466),
.C(n_488),
.Y(n_677)
);

NAND2x1p5_ASAP7_75t_L g678 ( 
.A(n_554),
.B(n_537),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_558),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_SL g680 ( 
.A1(n_627),
.A2(n_278),
.B1(n_359),
.B2(n_371),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_543),
.B(n_505),
.Y(n_681)
);

NAND2x1p5_ASAP7_75t_L g682 ( 
.A(n_554),
.B(n_505),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_532),
.Y(n_683)
);

NAND2x1p5_ASAP7_75t_L g684 ( 
.A(n_554),
.B(n_505),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_562),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_570),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_622),
.B(n_470),
.Y(n_687)
);

AO22x2_ASAP7_75t_L g688 ( 
.A1(n_644),
.A2(n_478),
.B1(n_18),
.B2(n_22),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_532),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_629),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_636),
.A2(n_470),
.B1(n_490),
.B2(n_441),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_571),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_605),
.Y(n_693)
);

OAI221xp5_ASAP7_75t_L g694 ( 
.A1(n_531),
.A2(n_503),
.B1(n_488),
.B2(n_485),
.C(n_466),
.Y(n_694)
);

AO22x2_ASAP7_75t_L g695 ( 
.A1(n_531),
.A2(n_544),
.B1(n_620),
.B2(n_560),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_574),
.Y(n_696)
);

AO22x2_ASAP7_75t_L g697 ( 
.A1(n_544),
.A2(n_16),
.B1(n_23),
.B2(n_24),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_532),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_575),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_587),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_595),
.A2(n_470),
.B1(n_455),
.B2(n_482),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_553),
.B(n_433),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_622),
.B(n_470),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_550),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_604),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_623),
.B(n_455),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_623),
.B(n_455),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_636),
.A2(n_318),
.B1(n_217),
.B2(n_215),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_606),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_617),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_619),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_621),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_655),
.B(n_455),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_631),
.B(n_530),
.Y(n_714)
);

OAI221xp5_ASAP7_75t_L g715 ( 
.A1(n_564),
.A2(n_485),
.B1(n_474),
.B2(n_479),
.C(n_299),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_648),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_636),
.A2(n_439),
.B1(n_441),
.B2(n_287),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_573),
.Y(n_718)
);

AO22x2_ASAP7_75t_L g719 ( 
.A1(n_620),
.A2(n_16),
.B1(n_23),
.B2(n_24),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_590),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_590),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_565),
.B(n_439),
.Y(n_722)
);

AO22x2_ASAP7_75t_L g723 ( 
.A1(n_560),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_605),
.Y(n_724)
);

NAND2x1p5_ASAP7_75t_L g725 ( 
.A(n_537),
.B(n_655),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_565),
.B(n_474),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_607),
.B(n_192),
.Y(n_727)
);

AO22x2_ASAP7_75t_L g728 ( 
.A1(n_528),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_728)
);

OAI221xp5_ASAP7_75t_L g729 ( 
.A1(n_530),
.A2(n_479),
.B1(n_313),
.B2(n_298),
.C(n_311),
.Y(n_729)
);

AO22x2_ASAP7_75t_L g730 ( 
.A1(n_551),
.A2(n_36),
.B1(n_39),
.B2(n_41),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_650),
.Y(n_731)
);

OAI221xp5_ASAP7_75t_L g732 ( 
.A1(n_647),
.A2(n_310),
.B1(n_308),
.B2(n_306),
.C(n_303),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_585),
.B(n_464),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_650),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_651),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_602),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_550),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_535),
.B(n_457),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_591),
.B(n_192),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_633),
.B(n_194),
.Y(n_740)
);

AO22x2_ASAP7_75t_L g741 ( 
.A1(n_551),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_597),
.Y(n_742)
);

AO22x2_ASAP7_75t_L g743 ( 
.A1(n_551),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_550),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_603),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_656),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_656),
.Y(n_747)
);

OR2x6_ASAP7_75t_L g748 ( 
.A(n_540),
.B(n_464),
.Y(n_748)
);

AO21x2_ASAP7_75t_L g749 ( 
.A1(n_608),
.A2(n_415),
.B(n_457),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_655),
.B(n_464),
.Y(n_750)
);

AO22x2_ASAP7_75t_L g751 ( 
.A1(n_551),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_579),
.B(n_194),
.Y(n_752)
);

OR2x6_ASAP7_75t_L g753 ( 
.A(n_540),
.B(n_557),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_593),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_569),
.B(n_459),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_594),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_654),
.Y(n_757)
);

AO22x2_ASAP7_75t_L g758 ( 
.A1(n_633),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_569),
.B(n_459),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_557),
.B(n_467),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_657),
.Y(n_761)
);

AO22x2_ASAP7_75t_L g762 ( 
.A1(n_609),
.A2(n_55),
.B1(n_57),
.B2(n_316),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_559),
.B(n_467),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_615),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_615),
.Y(n_765)
);

OAI221xp5_ASAP7_75t_L g766 ( 
.A1(n_586),
.A2(n_322),
.B1(n_318),
.B2(n_317),
.C(n_316),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_615),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_625),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_559),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_636),
.A2(n_275),
.B1(n_307),
.B2(n_295),
.Y(n_770)
);

INVxp33_ASAP7_75t_SL g771 ( 
.A(n_603),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_577),
.B(n_462),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_625),
.Y(n_773)
);

NAND2x1p5_ASAP7_75t_L g774 ( 
.A(n_537),
.B(n_462),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_577),
.B(n_467),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_625),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_628),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_628),
.B(n_472),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_626),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_592),
.B(n_472),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_645),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_595),
.B(n_476),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_561),
.Y(n_783)
);

OAI221xp5_ASAP7_75t_L g784 ( 
.A1(n_588),
.A2(n_317),
.B1(n_217),
.B2(n_215),
.C(n_351),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_561),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_609),
.B(n_200),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_535),
.B(n_476),
.Y(n_787)
);

OAI221xp5_ASAP7_75t_L g788 ( 
.A1(n_540),
.A2(n_196),
.B1(n_322),
.B2(n_351),
.C(n_327),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_540),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_613),
.A2(n_256),
.B1(n_282),
.B2(n_280),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_535),
.B(n_481),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_584),
.B(n_200),
.Y(n_792)
);

OAI221xp5_ASAP7_75t_L g793 ( 
.A1(n_572),
.A2(n_196),
.B1(n_327),
.B2(n_330),
.C(n_331),
.Y(n_793)
);

BUFx8_ASAP7_75t_L g794 ( 
.A(n_567),
.Y(n_794)
);

AO22x2_ASAP7_75t_L g795 ( 
.A1(n_572),
.A2(n_57),
.B1(n_347),
.B2(n_345),
.Y(n_795)
);

OAI221xp5_ASAP7_75t_L g796 ( 
.A1(n_652),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.C(n_335),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_777),
.B(n_614),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_780),
.B(n_634),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_775),
.B(n_760),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_669),
.B(n_539),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_670),
.B(n_539),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_SL g802 ( 
.A(n_660),
.B(n_567),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_722),
.B(n_539),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_702),
.B(n_652),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_714),
.B(n_658),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_726),
.B(n_653),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_675),
.B(n_542),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_727),
.B(n_547),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_778),
.B(n_739),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_769),
.B(n_547),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_790),
.B(n_547),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_790),
.B(n_548),
.Y(n_812)
);

NAND2xp33_ASAP7_75t_SL g813 ( 
.A(n_660),
.B(n_601),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_760),
.B(n_595),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_755),
.B(n_548),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_759),
.B(n_548),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_772),
.B(n_563),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_763),
.B(n_779),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_763),
.B(n_563),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_786),
.B(n_563),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_752),
.B(n_649),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_792),
.B(n_568),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_690),
.B(n_568),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_659),
.B(n_568),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_659),
.B(n_201),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_SL g826 ( 
.A(n_720),
.B(n_204),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_664),
.B(n_204),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_664),
.B(n_206),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_738),
.B(n_742),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_SL g830 ( 
.A(n_721),
.B(n_206),
.Y(n_830)
);

NAND2xp33_ASAP7_75t_SL g831 ( 
.A(n_789),
.B(n_207),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_733),
.B(n_717),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_717),
.B(n_208),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_770),
.B(n_208),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_770),
.B(n_787),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_787),
.B(n_210),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_705),
.B(n_595),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_791),
.B(n_210),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_791),
.B(n_662),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_663),
.B(n_212),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_748),
.B(n_595),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_709),
.B(n_595),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_SL g843 ( 
.A(n_681),
.B(n_218),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_693),
.B(n_649),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_668),
.B(n_218),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_671),
.B(n_270),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_SL g847 ( 
.A(n_681),
.B(n_270),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_676),
.B(n_314),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_710),
.B(n_596),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_679),
.B(n_315),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_685),
.B(n_315),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_711),
.B(n_596),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_712),
.B(n_596),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_686),
.B(n_596),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_692),
.B(n_319),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_696),
.B(n_319),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_699),
.B(n_596),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_700),
.B(n_320),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_736),
.B(n_320),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_672),
.B(n_324),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_724),
.B(n_324),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_673),
.B(n_740),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_691),
.B(n_326),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_695),
.B(n_639),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_691),
.B(n_326),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_716),
.B(n_329),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_661),
.B(n_665),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_661),
.B(n_337),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_665),
.B(n_337),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_695),
.B(n_666),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_771),
.B(n_338),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_764),
.B(n_338),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_748),
.B(n_630),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_765),
.B(n_339),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_666),
.B(n_639),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_767),
.B(n_339),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_768),
.B(n_350),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_773),
.B(n_776),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_781),
.B(n_350),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_673),
.B(n_332),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_673),
.B(n_680),
.Y(n_881)
);

NAND2xp33_ASAP7_75t_L g882 ( 
.A(n_678),
.B(n_545),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_SL g883 ( 
.A(n_687),
.B(n_526),
.Y(n_883)
);

NAND2xp33_ASAP7_75t_SL g884 ( 
.A(n_687),
.B(n_534),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_678),
.B(n_534),
.Y(n_885)
);

NAND2xp33_ASAP7_75t_SL g886 ( 
.A(n_703),
.B(n_581),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_706),
.B(n_642),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_706),
.B(n_642),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_SL g889 ( 
.A(n_703),
.B(n_582),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_SL g890 ( 
.A(n_707),
.B(n_582),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_732),
.B(n_335),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_680),
.B(n_582),
.Y(n_892)
);

NAND2xp33_ASAP7_75t_SL g893 ( 
.A(n_707),
.B(n_589),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_753),
.B(n_674),
.Y(n_894)
);

NAND2xp33_ASAP7_75t_SL g895 ( 
.A(n_701),
.B(n_589),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_754),
.B(n_612),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_756),
.B(n_612),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_757),
.B(n_612),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_761),
.B(n_258),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_782),
.B(n_274),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_796),
.B(n_345),
.Y(n_901)
);

NAND2xp33_ASAP7_75t_SL g902 ( 
.A(n_708),
.B(n_343),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_750),
.B(n_545),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_725),
.B(n_301),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_667),
.B(n_545),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_683),
.B(n_349),
.Y(n_906)
);

NAND2xp33_ASAP7_75t_SL g907 ( 
.A(n_745),
.B(n_342),
.Y(n_907)
);

NAND2xp33_ASAP7_75t_SL g908 ( 
.A(n_708),
.B(n_342),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_713),
.B(n_545),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_713),
.B(n_545),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_689),
.B(n_233),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_731),
.B(n_545),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_698),
.B(n_246),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_734),
.B(n_735),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_704),
.B(n_246),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_737),
.B(n_246),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_744),
.B(n_296),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_SL g918 ( 
.A(n_749),
.B(n_347),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_748),
.B(n_753),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_682),
.B(n_296),
.Y(n_920)
);

NAND2xp33_ASAP7_75t_SL g921 ( 
.A(n_749),
.B(n_630),
.Y(n_921)
);

NAND2xp33_ASAP7_75t_SL g922 ( 
.A(n_794),
.B(n_632),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_682),
.B(n_296),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_684),
.B(n_638),
.Y(n_924)
);

NAND2xp33_ASAP7_75t_SL g925 ( 
.A(n_746),
.B(n_637),
.Y(n_925)
);

NAND2xp33_ASAP7_75t_SL g926 ( 
.A(n_747),
.B(n_637),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_774),
.B(n_578),
.Y(n_927)
);

NAND2xp33_ASAP7_75t_SL g928 ( 
.A(n_783),
.B(n_641),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_753),
.B(n_618),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_774),
.B(n_794),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_785),
.B(n_578),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_729),
.B(n_624),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_793),
.B(n_580),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_788),
.B(n_481),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_766),
.B(n_529),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_SL g936 ( 
.A(n_795),
.B(n_541),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_715),
.B(n_529),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_674),
.B(n_541),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_784),
.B(n_533),
.Y(n_939)
);

NAND2xp33_ASAP7_75t_SL g940 ( 
.A(n_795),
.B(n_730),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_688),
.B(n_533),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_688),
.B(n_546),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_730),
.B(n_546),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_741),
.B(n_598),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_799),
.B(n_762),
.Y(n_945)
);

NOR4xp25_ASAP7_75t_L g946 ( 
.A(n_832),
.B(n_741),
.C(n_751),
.D(n_743),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_875),
.A2(n_576),
.B(n_598),
.Y(n_947)
);

NOR2x1_ASAP7_75t_SL g948 ( 
.A(n_885),
.B(n_566),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_862),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_804),
.B(n_694),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_821),
.A2(n_576),
.B(n_598),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_798),
.A2(n_576),
.B(n_610),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_901),
.A2(n_677),
.B(n_751),
.C(n_743),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_914),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_887),
.A2(n_610),
.B(n_566),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_810),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_829),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_797),
.B(n_60),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_839),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_878),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_880),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_818),
.B(n_61),
.Y(n_962)
);

AOI21x1_ASAP7_75t_SL g963 ( 
.A1(n_864),
.A2(n_697),
.B(n_719),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_870),
.B(n_762),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_919),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_813),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_895),
.A2(n_610),
.B(n_611),
.Y(n_967)
);

AOI21xp33_ASAP7_75t_L g968 ( 
.A1(n_867),
.A2(n_719),
.B(n_723),
.Y(n_968)
);

OAI22x1_ASAP7_75t_L g969 ( 
.A1(n_891),
.A2(n_833),
.B1(n_881),
.B2(n_894),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_809),
.B(n_723),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_800),
.A2(n_758),
.B1(n_728),
.B2(n_482),
.Y(n_971)
);

AO31x2_ASAP7_75t_L g972 ( 
.A1(n_905),
.A2(n_758),
.A3(n_728),
.B(n_482),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_895),
.A2(n_611),
.B(n_600),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_SL g974 ( 
.A1(n_814),
.A2(n_600),
.B(n_549),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_806),
.B(n_482),
.Y(n_975)
);

AO31x2_ASAP7_75t_L g976 ( 
.A1(n_937),
.A2(n_482),
.A3(n_79),
.B(n_89),
.Y(n_976)
);

AO31x2_ASAP7_75t_L g977 ( 
.A1(n_903),
.A2(n_482),
.A3(n_90),
.B(n_97),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_803),
.B(n_78),
.Y(n_978)
);

OA21x2_ASAP7_75t_L g979 ( 
.A1(n_909),
.A2(n_482),
.B(n_123),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_820),
.A2(n_549),
.B(n_126),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_801),
.B(n_113),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_819),
.A2(n_549),
.B(n_132),
.Y(n_982)
);

OR2x6_ASAP7_75t_L g983 ( 
.A(n_919),
.B(n_130),
.Y(n_983)
);

AO31x2_ASAP7_75t_L g984 ( 
.A1(n_910),
.A2(n_482),
.A3(n_142),
.B(n_156),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_873),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_929),
.Y(n_986)
);

NAND2x1p5_ASAP7_75t_L g987 ( 
.A(n_841),
.B(n_919),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_935),
.A2(n_939),
.B(n_847),
.Y(n_988)
);

AO21x1_ASAP7_75t_L g989 ( 
.A1(n_940),
.A2(n_918),
.B(n_921),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_844),
.B(n_815),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_841),
.B(n_929),
.Y(n_991)
);

AO31x2_ASAP7_75t_L g992 ( 
.A1(n_837),
.A2(n_849),
.A3(n_852),
.B(n_857),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_823),
.B(n_938),
.Y(n_993)
);

AND3x4_ASAP7_75t_L g994 ( 
.A(n_929),
.B(n_841),
.C(n_907),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_816),
.B(n_817),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_859),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_811),
.A2(n_812),
.B1(n_835),
.B2(n_943),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_807),
.B(n_930),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_940),
.A2(n_936),
.B(n_853),
.C(n_842),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_808),
.B(n_822),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_936),
.A2(n_869),
.B1(n_868),
.B2(n_863),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_802),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_941),
.B(n_854),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_861),
.Y(n_1004)
);

AO31x2_ASAP7_75t_L g1005 ( 
.A1(n_912),
.A2(n_931),
.A3(n_847),
.B(n_843),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_942),
.B(n_892),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_SL g1007 ( 
.A1(n_944),
.A2(n_923),
.B(n_920),
.C(n_865),
.Y(n_1007)
);

NAND2xp33_ASAP7_75t_R g1008 ( 
.A(n_826),
.B(n_830),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_866),
.B(n_871),
.Y(n_1009)
);

NOR2xp67_ASAP7_75t_L g1010 ( 
.A(n_860),
.B(n_906),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_831),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_802),
.Y(n_1012)
);

AOI211x1_ASAP7_75t_L g1013 ( 
.A1(n_834),
.A2(n_934),
.B(n_845),
.C(n_846),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_843),
.A2(n_908),
.B(n_902),
.C(n_889),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_933),
.A2(n_893),
.B(n_890),
.Y(n_1015)
);

NAND2x1p5_ASAP7_75t_L g1016 ( 
.A(n_824),
.B(n_927),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_932),
.B(n_900),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_872),
.B(n_874),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_882),
.A2(n_890),
.B(n_893),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_876),
.B(n_879),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_883),
.A2(n_884),
.B(n_886),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_SL g1022 ( 
.A1(n_840),
.A2(n_855),
.B(n_858),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_883),
.A2(n_886),
.B(n_884),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_889),
.A2(n_925),
.B(n_926),
.Y(n_1024)
);

OAI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_836),
.A2(n_838),
.B1(n_827),
.B2(n_828),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_896),
.Y(n_1026)
);

BUFx4f_ASAP7_75t_L g1027 ( 
.A(n_922),
.Y(n_1027)
);

AO21x2_ASAP7_75t_L g1028 ( 
.A1(n_897),
.A2(n_898),
.B(n_904),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_877),
.A2(n_848),
.B(n_850),
.C(n_851),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_899),
.A2(n_825),
.B(n_856),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_928),
.A2(n_911),
.B(n_913),
.Y(n_1031)
);

AO31x2_ASAP7_75t_L g1032 ( 
.A1(n_928),
.A2(n_915),
.A3(n_916),
.B(n_917),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_799),
.B(n_821),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_799),
.B(n_599),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_810),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_914),
.Y(n_1036)
);

AO32x2_ASAP7_75t_L g1037 ( 
.A1(n_940),
.A2(n_708),
.A3(n_599),
.B1(n_640),
.B2(n_936),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_914),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_799),
.B(n_821),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_799),
.B(n_821),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_862),
.Y(n_1041)
);

NOR2xp67_ASAP7_75t_L g1042 ( 
.A(n_804),
.B(n_690),
.Y(n_1042)
);

BUFx12f_ASAP7_75t_L g1043 ( 
.A(n_919),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_867),
.A2(n_821),
.B1(n_799),
.B2(n_543),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_914),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_813),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_799),
.B(n_821),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_799),
.B(n_821),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_SL g1049 ( 
.A1(n_864),
.A2(n_870),
.B(n_799),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_870),
.A2(n_867),
.B(n_821),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_799),
.B(n_821),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_862),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_799),
.B(n_821),
.Y(n_1053)
);

AND2x2_ASAP7_75t_SL g1054 ( 
.A(n_881),
.B(n_613),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_799),
.B(n_821),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_799),
.B(n_821),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_799),
.B(n_821),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_813),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_797),
.B(n_718),
.Y(n_1059)
);

AOI31xp67_ASAP7_75t_L g1060 ( 
.A1(n_805),
.A2(n_832),
.A3(n_798),
.B(n_864),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_799),
.B(n_821),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_799),
.B(n_821),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_804),
.B(n_629),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_887),
.A2(n_888),
.B(n_924),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_870),
.A2(n_867),
.B(n_821),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_862),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_799),
.B(n_821),
.Y(n_1067)
);

O2A1O1Ixp5_ASAP7_75t_L g1068 ( 
.A1(n_821),
.A2(n_727),
.B(n_832),
.C(n_920),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_914),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_914),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_SL g1071 ( 
.A1(n_867),
.A2(n_943),
.B(n_944),
.C(n_864),
.Y(n_1071)
);

INVx6_ASAP7_75t_L g1072 ( 
.A(n_965),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1034),
.B(n_1033),
.Y(n_1073)
);

AO21x1_ASAP7_75t_L g1074 ( 
.A1(n_997),
.A2(n_1024),
.B(n_988),
.Y(n_1074)
);

OA21x2_ASAP7_75t_L g1075 ( 
.A1(n_988),
.A2(n_1015),
.B(n_1050),
.Y(n_1075)
);

OA21x2_ASAP7_75t_L g1076 ( 
.A1(n_1015),
.A2(n_1065),
.B(n_1050),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_954),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_1059),
.B(n_1063),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_956),
.Y(n_1079)
);

AOI22x1_ASAP7_75t_L g1080 ( 
.A1(n_969),
.A2(n_1049),
.B1(n_1024),
.B2(n_1016),
.Y(n_1080)
);

OA21x2_ASAP7_75t_L g1081 ( 
.A1(n_1065),
.A2(n_1064),
.B(n_1068),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_960),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_986),
.B(n_991),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1033),
.B(n_1039),
.Y(n_1084)
);

OR2x6_ASAP7_75t_L g1085 ( 
.A(n_983),
.B(n_987),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_SL g1086 ( 
.A1(n_1054),
.A2(n_946),
.B1(n_994),
.B2(n_1058),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_966),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1038),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1039),
.B(n_1040),
.Y(n_1089)
);

AO21x2_ASAP7_75t_L g1090 ( 
.A1(n_997),
.A2(n_989),
.B(n_1014),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1040),
.B(n_1047),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_959),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1047),
.B(n_1048),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_953),
.A2(n_1025),
.B(n_1029),
.C(n_1011),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_968),
.A2(n_1044),
.B1(n_1053),
.B2(n_1056),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_968),
.A2(n_1044),
.B1(n_1048),
.B2(n_1051),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1035),
.B(n_949),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1051),
.A2(n_1055),
.B(n_1057),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_985),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1053),
.B(n_1055),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_965),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_987),
.Y(n_1102)
);

OA21x2_ASAP7_75t_L g1103 ( 
.A1(n_1017),
.A2(n_999),
.B(n_1062),
.Y(n_1103)
);

CKINVDCx9p33_ASAP7_75t_R g1104 ( 
.A(n_1012),
.Y(n_1104)
);

CKINVDCx6p67_ASAP7_75t_R g1105 ( 
.A(n_1043),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1036),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_1022),
.A2(n_1071),
.B(n_970),
.C(n_1018),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1045),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1056),
.A2(n_1067),
.B1(n_1062),
.B2(n_1061),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_961),
.A2(n_1042),
.B1(n_1009),
.B2(n_996),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_990),
.A2(n_1057),
.B(n_1067),
.Y(n_1111)
);

AO21x2_ASAP7_75t_L g1112 ( 
.A1(n_1007),
.A2(n_1017),
.B(n_1061),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_990),
.B(n_1041),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_1052),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_974),
.A2(n_1000),
.B(n_951),
.Y(n_1115)
);

INVxp67_ASAP7_75t_L g1116 ( 
.A(n_1066),
.Y(n_1116)
);

AO21x1_ASAP7_75t_L g1117 ( 
.A1(n_958),
.A2(n_945),
.B(n_962),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1069),
.A2(n_1070),
.B1(n_1001),
.B2(n_945),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1000),
.A2(n_967),
.B(n_973),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_993),
.B(n_957),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_1027),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_950),
.A2(n_971),
.B(n_970),
.C(n_964),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_955),
.A2(n_952),
.B(n_982),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1003),
.A2(n_1060),
.B(n_995),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_995),
.B(n_1020),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_947),
.A2(n_980),
.B(n_1003),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_998),
.B(n_1004),
.Y(n_1127)
);

BUFx10_ASAP7_75t_L g1128 ( 
.A(n_1046),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_964),
.B(n_1020),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1018),
.B(n_1006),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_SL g1131 ( 
.A1(n_978),
.A2(n_1006),
.B1(n_1027),
.B2(n_983),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_981),
.A2(n_948),
.B(n_1031),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_1002),
.Y(n_1133)
);

AO21x2_ASAP7_75t_L g1134 ( 
.A1(n_1031),
.A2(n_1028),
.B(n_946),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_983),
.B(n_1006),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_979),
.A2(n_963),
.B(n_1016),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1137)
);

NAND3xp33_ASAP7_75t_L g1138 ( 
.A(n_1008),
.B(n_975),
.C(n_1026),
.Y(n_1138)
);

OAI211xp5_ASAP7_75t_L g1139 ( 
.A1(n_1030),
.A2(n_979),
.B(n_972),
.C(n_1037),
.Y(n_1139)
);

OA21x2_ASAP7_75t_L g1140 ( 
.A1(n_1037),
.A2(n_1005),
.B(n_976),
.Y(n_1140)
);

OAI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_972),
.A2(n_1037),
.B1(n_1032),
.B2(n_1028),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_972),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1032),
.Y(n_1143)
);

INVx6_ASAP7_75t_L g1144 ( 
.A(n_1032),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_992),
.A2(n_984),
.B(n_977),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_976),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_977),
.A2(n_1068),
.B(n_821),
.Y(n_1147)
);

AO21x2_ASAP7_75t_L g1148 ( 
.A1(n_984),
.A2(n_988),
.B(n_1015),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_965),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_986),
.B(n_991),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1059),
.B(n_718),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_949),
.Y(n_1152)
);

OR2x6_ASAP7_75t_L g1153 ( 
.A(n_983),
.B(n_987),
.Y(n_1153)
);

OA21x2_ASAP7_75t_L g1154 ( 
.A1(n_988),
.A2(n_1015),
.B(n_1050),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_983),
.B(n_987),
.Y(n_1155)
);

AOI221xp5_ASAP7_75t_L g1156 ( 
.A1(n_968),
.A2(n_901),
.B1(n_891),
.B2(n_551),
.C(n_674),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_954),
.Y(n_1157)
);

OA21x2_ASAP7_75t_L g1158 ( 
.A1(n_988),
.A2(n_1015),
.B(n_1050),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_990),
.B(n_1033),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1034),
.B(n_1033),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1034),
.B(n_1033),
.Y(n_1161)
);

AO21x2_ASAP7_75t_L g1162 ( 
.A1(n_988),
.A2(n_1015),
.B(n_1024),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_986),
.B(n_991),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1034),
.B(n_1033),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_949),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1068),
.A2(n_821),
.B(n_990),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_949),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_966),
.Y(n_1168)
);

OA21x2_ASAP7_75t_L g1169 ( 
.A1(n_988),
.A2(n_1015),
.B(n_1050),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1035),
.B(n_777),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_956),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_966),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_968),
.A2(n_940),
.B1(n_730),
.B2(n_743),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_954),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_988),
.A2(n_1015),
.B(n_1050),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_986),
.B(n_991),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_965),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1059),
.B(n_718),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_954),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1033),
.A2(n_821),
.B(n_867),
.C(n_1039),
.Y(n_1180)
);

OA21x2_ASAP7_75t_L g1181 ( 
.A1(n_988),
.A2(n_1015),
.B(n_1050),
.Y(n_1181)
);

AOI221x1_ASAP7_75t_L g1182 ( 
.A1(n_968),
.A2(n_940),
.B1(n_953),
.B2(n_969),
.C(n_918),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_965),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_985),
.B(n_986),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_949),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1033),
.A2(n_1040),
.B1(n_1047),
.B2(n_1039),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_968),
.A2(n_940),
.B1(n_730),
.B2(n_743),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1035),
.B(n_777),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1034),
.B(n_1033),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_966),
.Y(n_1190)
);

AO21x1_ASAP7_75t_L g1191 ( 
.A1(n_997),
.A2(n_821),
.B(n_940),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1019),
.A2(n_1023),
.B(n_1021),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1019),
.A2(n_1023),
.B(n_1021),
.Y(n_1193)
);

BUFx8_ASAP7_75t_L g1194 ( 
.A(n_949),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_965),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_983),
.B(n_987),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_1114),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1170),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1142),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1194),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1085),
.B(n_1153),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1087),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1077),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1152),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_1165),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1121),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1088),
.Y(n_1207)
);

BUFx2_ASAP7_75t_SL g1208 ( 
.A(n_1121),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1167),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1102),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1088),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1125),
.B(n_1111),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1188),
.Y(n_1213)
);

INVx6_ASAP7_75t_L g1214 ( 
.A(n_1194),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1102),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1143),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1072),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1097),
.Y(n_1218)
);

INVx5_ASAP7_75t_L g1219 ( 
.A(n_1085),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1098),
.A2(n_1180),
.B(n_1115),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_1147),
.A2(n_1145),
.B(n_1124),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1194),
.Y(n_1222)
);

INVx6_ASAP7_75t_L g1223 ( 
.A(n_1195),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1185),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1144),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1144),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_1127),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1101),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1144),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1074),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_1087),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1134),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1134),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1090),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1156),
.A2(n_1117),
.B1(n_1130),
.B2(n_1178),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1129),
.B(n_1122),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1090),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1104),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1157),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1174),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1179),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1102),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1106),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1108),
.Y(n_1244)
);

INVx5_ASAP7_75t_L g1245 ( 
.A(n_1085),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1079),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1122),
.B(n_1159),
.Y(n_1247)
);

AO21x2_ASAP7_75t_L g1248 ( 
.A1(n_1141),
.A2(n_1119),
.B(n_1145),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_SL g1249 ( 
.A1(n_1151),
.A2(n_1130),
.B1(n_1135),
.B2(n_1078),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1101),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1153),
.B(n_1155),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1078),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1084),
.A2(n_1100),
.B1(n_1091),
.B2(n_1093),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1153),
.B(n_1155),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1149),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1103),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1103),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1125),
.B(n_1109),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1177),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1162),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1116),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1109),
.B(n_1095),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1095),
.B(n_1096),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1072),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1082),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1072),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1171),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1104),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1076),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1076),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1092),
.Y(n_1271)
);

INVx4_ASAP7_75t_SL g1272 ( 
.A(n_1155),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1076),
.Y(n_1273)
);

OR2x6_ASAP7_75t_L g1274 ( 
.A(n_1196),
.B(n_1132),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1075),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1120),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1075),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1166),
.A2(n_1139),
.B(n_1146),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1075),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1154),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1073),
.B(n_1160),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1161),
.B(n_1164),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1196),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1149),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1099),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1099),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1096),
.B(n_1089),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1099),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1196),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1083),
.B(n_1150),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_R g1291 ( 
.A(n_1168),
.B(n_1190),
.Y(n_1291)
);

NOR2x1_ASAP7_75t_SL g1292 ( 
.A(n_1112),
.B(n_1148),
.Y(n_1292)
);

CKINVDCx14_ASAP7_75t_R g1293 ( 
.A(n_1105),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1158),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1189),
.B(n_1181),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1169),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1180),
.A2(n_1094),
.B(n_1186),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1177),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1192),
.A2(n_1193),
.B(n_1123),
.Y(n_1299)
);

XNOR2xp5_ASAP7_75t_L g1300 ( 
.A(n_1231),
.B(n_1168),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1281),
.B(n_1113),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1282),
.B(n_1118),
.Y(n_1302)
);

NAND2xp33_ASAP7_75t_R g1303 ( 
.A(n_1291),
.B(n_1190),
.Y(n_1303)
);

CKINVDCx12_ASAP7_75t_R g1304 ( 
.A(n_1249),
.Y(n_1304)
);

NAND2xp33_ASAP7_75t_R g1305 ( 
.A(n_1202),
.B(n_1172),
.Y(n_1305)
);

OR2x6_ASAP7_75t_L g1306 ( 
.A(n_1208),
.B(n_1133),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1253),
.B(n_1107),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1272),
.B(n_1201),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_R g1309 ( 
.A(n_1202),
.B(n_1172),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_R g1310 ( 
.A(n_1293),
.B(n_1105),
.Y(n_1310)
);

OR2x6_ASAP7_75t_L g1311 ( 
.A(n_1208),
.B(n_1086),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_1254),
.B(n_1195),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1218),
.Y(n_1313)
);

XNOR2xp5_ASAP7_75t_L g1314 ( 
.A(n_1200),
.B(n_1110),
.Y(n_1314)
);

NAND2xp33_ASAP7_75t_R g1315 ( 
.A(n_1238),
.B(n_1268),
.Y(n_1315)
);

OR2x6_ASAP7_75t_L g1316 ( 
.A(n_1254),
.B(n_1195),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_R g1317 ( 
.A(n_1206),
.B(n_1128),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1212),
.B(n_1137),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_R g1319 ( 
.A(n_1206),
.B(n_1128),
.Y(n_1319)
);

NAND2xp33_ASAP7_75t_R g1320 ( 
.A(n_1238),
.B(n_1268),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1265),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1204),
.Y(n_1322)
);

INVx8_ASAP7_75t_L g1323 ( 
.A(n_1259),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1228),
.Y(n_1324)
);

BUFx10_ASAP7_75t_L g1325 ( 
.A(n_1214),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1201),
.B(n_1177),
.Y(n_1326)
);

XOR2xp5_ASAP7_75t_L g1327 ( 
.A(n_1276),
.B(n_1131),
.Y(n_1327)
);

XOR2x2_ASAP7_75t_L g1328 ( 
.A(n_1224),
.B(n_1138),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1251),
.B(n_1177),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1261),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1251),
.B(n_1183),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1290),
.B(n_1183),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1204),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1198),
.B(n_1173),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_R g1335 ( 
.A(n_1214),
.B(n_1128),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1213),
.B(n_1252),
.Y(n_1336)
);

CKINVDCx12_ASAP7_75t_R g1337 ( 
.A(n_1254),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1205),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1205),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1290),
.B(n_1183),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1227),
.B(n_1258),
.Y(n_1341)
);

NAND2xp33_ASAP7_75t_R g1342 ( 
.A(n_1209),
.B(n_1163),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1258),
.B(n_1173),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_R g1344 ( 
.A(n_1214),
.B(n_1150),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_R g1345 ( 
.A(n_1214),
.B(n_1150),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1199),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_R g1347 ( 
.A(n_1210),
.B(n_1176),
.Y(n_1347)
);

XOR2xp5_ASAP7_75t_L g1348 ( 
.A(n_1222),
.B(n_1080),
.Y(n_1348)
);

XNOR2xp5_ASAP7_75t_L g1349 ( 
.A(n_1222),
.B(n_1163),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1235),
.B(n_1163),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_R g1351 ( 
.A(n_1210),
.B(n_1083),
.Y(n_1351)
);

NAND2xp33_ASAP7_75t_R g1352 ( 
.A(n_1209),
.B(n_1176),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1287),
.B(n_1187),
.Y(n_1353)
);

INVxp67_ASAP7_75t_L g1354 ( 
.A(n_1197),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1236),
.B(n_1112),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1254),
.B(n_1083),
.Y(n_1356)
);

XNOR2xp5_ASAP7_75t_L g1357 ( 
.A(n_1283),
.B(n_1182),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1289),
.B(n_1136),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1228),
.Y(n_1359)
);

NAND2xp33_ASAP7_75t_R g1360 ( 
.A(n_1289),
.B(n_1181),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1236),
.B(n_1191),
.Y(n_1361)
);

CKINVDCx8_ASAP7_75t_R g1362 ( 
.A(n_1259),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_1250),
.Y(n_1363)
);

INVxp67_ASAP7_75t_L g1364 ( 
.A(n_1250),
.Y(n_1364)
);

NAND2xp33_ASAP7_75t_R g1365 ( 
.A(n_1215),
.B(n_1181),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1216),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1219),
.B(n_1136),
.Y(n_1367)
);

BUFx10_ASAP7_75t_L g1368 ( 
.A(n_1217),
.Y(n_1368)
);

XOR2xp5_ASAP7_75t_L g1369 ( 
.A(n_1247),
.B(n_1184),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1262),
.B(n_1175),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1219),
.B(n_1192),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1262),
.B(n_1297),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1219),
.B(n_1148),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_R g1374 ( 
.A(n_1242),
.B(n_1169),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1255),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1219),
.B(n_1245),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1247),
.B(n_1175),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_R g1378 ( 
.A(n_1242),
.B(n_1081),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1219),
.B(n_1126),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1245),
.B(n_1123),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_1255),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1271),
.Y(n_1382)
);

NAND2xp33_ASAP7_75t_SL g1383 ( 
.A(n_1263),
.B(n_1243),
.Y(n_1383)
);

OR2x6_ASAP7_75t_L g1384 ( 
.A(n_1274),
.B(n_1081),
.Y(n_1384)
);

NAND2xp33_ASAP7_75t_R g1385 ( 
.A(n_1274),
.B(n_1263),
.Y(n_1385)
);

NAND2xp33_ASAP7_75t_R g1386 ( 
.A(n_1274),
.B(n_1140),
.Y(n_1386)
);

OR2x6_ASAP7_75t_L g1387 ( 
.A(n_1274),
.B(n_1140),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_R g1388 ( 
.A(n_1223),
.B(n_1284),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1217),
.B(n_1264),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_R g1390 ( 
.A(n_1223),
.B(n_1284),
.Y(n_1390)
);

XOR2xp5_ASAP7_75t_L g1391 ( 
.A(n_1295),
.B(n_1230),
.Y(n_1391)
);

XNOR2xp5_ASAP7_75t_L g1392 ( 
.A(n_1264),
.B(n_1266),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1298),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_SL g1394 ( 
.A(n_1245),
.B(n_1223),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1298),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1244),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_R g1397 ( 
.A(n_1223),
.B(n_1266),
.Y(n_1397)
);

NAND2xp33_ASAP7_75t_R g1398 ( 
.A(n_1295),
.B(n_1288),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_R g1399 ( 
.A(n_1288),
.B(n_1259),
.Y(n_1399)
);

XOR2xp5_ASAP7_75t_L g1400 ( 
.A(n_1230),
.B(n_1225),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1246),
.Y(n_1401)
);

CKINVDCx6p67_ASAP7_75t_R g1402 ( 
.A(n_1245),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1245),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_R g1404 ( 
.A(n_1288),
.B(n_1267),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1240),
.B(n_1241),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1377),
.B(n_1260),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1370),
.B(n_1260),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1346),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1366),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1358),
.B(n_1256),
.Y(n_1410)
);

NOR2x1_ASAP7_75t_SL g1411 ( 
.A(n_1387),
.B(n_1278),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1355),
.B(n_1387),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1338),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1321),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1378),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1307),
.A2(n_1220),
.B(n_1299),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1396),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1341),
.B(n_1275),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1309),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1372),
.B(n_1275),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1382),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1313),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1358),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1365),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1391),
.B(n_1277),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1301),
.B(n_1354),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1318),
.B(n_1203),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1401),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1384),
.B(n_1232),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1384),
.B(n_1277),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1361),
.B(n_1279),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1373),
.B(n_1279),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1302),
.B(n_1207),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1373),
.B(n_1280),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1336),
.B(n_1211),
.Y(n_1435)
);

OAI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1348),
.A2(n_1229),
.B1(n_1226),
.B2(n_1234),
.C(n_1237),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1371),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1405),
.Y(n_1438)
);

NAND2x1_ASAP7_75t_L g1439 ( 
.A(n_1376),
.B(n_1256),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1371),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1367),
.B(n_1257),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1404),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1339),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1330),
.B(n_1239),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1367),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1350),
.A2(n_1229),
.B1(n_1226),
.B2(n_1278),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1380),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1374),
.Y(n_1448)
);

AND2x4_ASAP7_75t_SL g1449 ( 
.A(n_1402),
.B(n_1257),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1308),
.B(n_1356),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1379),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1344),
.B(n_1239),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1383),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1333),
.B(n_1328),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1311),
.A2(n_1327),
.B1(n_1400),
.B2(n_1322),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1357),
.B(n_1296),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1389),
.Y(n_1457)
);

BUFx2_ASAP7_75t_SL g1458 ( 
.A(n_1362),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1311),
.A2(n_1278),
.B1(n_1286),
.B2(n_1285),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1337),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_1398),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1353),
.B(n_1343),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1315),
.Y(n_1463)
);

AND2x2_ASAP7_75t_SL g1464 ( 
.A(n_1446),
.B(n_1394),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_SL g1465 ( 
.A(n_1453),
.B(n_1312),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1408),
.Y(n_1466)
);

NAND4xp25_ASAP7_75t_L g1467 ( 
.A(n_1426),
.B(n_1334),
.C(n_1320),
.D(n_1303),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1449),
.Y(n_1468)
);

NAND4xp25_ASAP7_75t_L g1469 ( 
.A(n_1454),
.B(n_1305),
.C(n_1385),
.D(n_1342),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1408),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1409),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1449),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1432),
.B(n_1221),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1439),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1407),
.B(n_1233),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1432),
.B(n_1248),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1429),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1437),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1414),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1421),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1414),
.Y(n_1481)
);

AND2x2_ASAP7_75t_SL g1482 ( 
.A(n_1448),
.B(n_1403),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_1406),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1428),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1434),
.B(n_1248),
.Y(n_1485)
);

AOI211xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1436),
.A2(n_1304),
.B(n_1364),
.C(n_1381),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_1429),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_L g1488 ( 
.A(n_1416),
.B(n_1352),
.C(n_1314),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1441),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1416),
.A2(n_1292),
.B(n_1248),
.Y(n_1490)
);

OAI211xp5_ASAP7_75t_L g1491 ( 
.A1(n_1455),
.A2(n_1317),
.B(n_1319),
.C(n_1335),
.Y(n_1491)
);

NAND4xp25_ASAP7_75t_SL g1492 ( 
.A(n_1442),
.B(n_1393),
.C(n_1360),
.D(n_1310),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1407),
.B(n_1269),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1437),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1434),
.B(n_1269),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1430),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1417),
.Y(n_1497)
);

AOI33xp33_ASAP7_75t_L g1498 ( 
.A1(n_1456),
.A2(n_1326),
.A3(n_1329),
.B1(n_1331),
.B2(n_1340),
.B3(n_1332),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1431),
.B(n_1270),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1417),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1421),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1430),
.B(n_1273),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1449),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_SL g1504 ( 
.A(n_1452),
.B(n_1425),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1441),
.B(n_1294),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1483),
.B(n_1431),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1496),
.B(n_1424),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1496),
.B(n_1425),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1483),
.B(n_1420),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1480),
.B(n_1420),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1496),
.B(n_1423),
.Y(n_1511)
);

NAND2x1p5_ASAP7_75t_L g1512 ( 
.A(n_1472),
.B(n_1448),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1473),
.B(n_1423),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1480),
.B(n_1456),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1501),
.B(n_1413),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1477),
.B(n_1406),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1501),
.B(n_1418),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1484),
.Y(n_1518)
);

NOR2x1p5_ASAP7_75t_L g1519 ( 
.A(n_1469),
.B(n_1461),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1479),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1474),
.B(n_1411),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1473),
.B(n_1423),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1473),
.B(n_1411),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1477),
.B(n_1445),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1493),
.Y(n_1525)
);

NOR2xp67_ASAP7_75t_L g1526 ( 
.A(n_1474),
.B(n_1463),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1477),
.B(n_1412),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1466),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1487),
.B(n_1445),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1487),
.B(n_1412),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1487),
.B(n_1440),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1466),
.Y(n_1532)
);

INVx4_ASAP7_75t_L g1533 ( 
.A(n_1472),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1470),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1489),
.B(n_1440),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1489),
.B(n_1447),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1470),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1499),
.B(n_1443),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1499),
.B(n_1447),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1471),
.Y(n_1540)
);

AND2x2_ASAP7_75t_SL g1541 ( 
.A(n_1464),
.B(n_1415),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1471),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1475),
.B(n_1418),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1476),
.B(n_1410),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1476),
.B(n_1410),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1481),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1494),
.B(n_1410),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1541),
.B(n_1526),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1518),
.B(n_1467),
.Y(n_1549)
);

NAND2xp33_ASAP7_75t_R g1550 ( 
.A(n_1507),
.B(n_1419),
.Y(n_1550)
);

AO221x2_ASAP7_75t_L g1551 ( 
.A1(n_1514),
.A2(n_1488),
.B1(n_1486),
.B2(n_1460),
.C(n_1467),
.Y(n_1551)
);

NAND2xp33_ASAP7_75t_SL g1552 ( 
.A(n_1519),
.B(n_1498),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1515),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1541),
.A2(n_1464),
.B1(n_1488),
.B2(n_1492),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1541),
.A2(n_1464),
.B1(n_1492),
.B2(n_1469),
.Y(n_1555)
);

AO221x2_ASAP7_75t_L g1556 ( 
.A1(n_1514),
.A2(n_1486),
.B1(n_1460),
.B2(n_1504),
.C(n_1464),
.Y(n_1556)
);

OAI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1526),
.A2(n_1491),
.B1(n_1484),
.B2(n_1457),
.C(n_1442),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1538),
.B(n_1422),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1527),
.B(n_1504),
.Y(n_1559)
);

NAND2xp33_ASAP7_75t_SL g1560 ( 
.A(n_1519),
.B(n_1498),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1533),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_R g1562 ( 
.A(n_1533),
.B(n_1300),
.Y(n_1562)
);

OAI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1509),
.A2(n_1453),
.B1(n_1415),
.B2(n_1312),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1525),
.B(n_1497),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1510),
.B(n_1506),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1538),
.B(n_1505),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1508),
.B(n_1505),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_SL g1568 ( 
.A(n_1508),
.B(n_1345),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1515),
.B(n_1505),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1509),
.B(n_1502),
.Y(n_1570)
);

AO221x2_ASAP7_75t_L g1571 ( 
.A1(n_1506),
.A2(n_1504),
.B1(n_1369),
.B2(n_1462),
.C(n_1497),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1544),
.B(n_1502),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1510),
.B(n_1502),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1543),
.B(n_1495),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1512),
.B(n_1482),
.Y(n_1575)
);

NOR2x1_ASAP7_75t_L g1576 ( 
.A(n_1533),
.B(n_1491),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1543),
.B(n_1495),
.Y(n_1577)
);

OAI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1512),
.A2(n_1316),
.B1(n_1451),
.B2(n_1472),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1533),
.B(n_1465),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1544),
.B(n_1482),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1539),
.B(n_1507),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1539),
.B(n_1495),
.Y(n_1582)
);

NAND2xp33_ASAP7_75t_SL g1583 ( 
.A(n_1511),
.B(n_1388),
.Y(n_1583)
);

INVxp67_ASAP7_75t_SL g1584 ( 
.A(n_1516),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_SL g1585 ( 
.A(n_1512),
.B(n_1482),
.Y(n_1585)
);

NAND2xp33_ASAP7_75t_SL g1586 ( 
.A(n_1511),
.B(n_1390),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1517),
.B(n_1500),
.Y(n_1587)
);

CKINVDCx16_ASAP7_75t_R g1588 ( 
.A(n_1550),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1549),
.B(n_1527),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1564),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1562),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1552),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1581),
.B(n_1530),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1556),
.A2(n_1482),
.B1(n_1451),
.B2(n_1523),
.Y(n_1594)
);

OAI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1554),
.A2(n_1386),
.B1(n_1504),
.B2(n_1306),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1556),
.A2(n_1523),
.B1(n_1450),
.B2(n_1485),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1564),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1565),
.B(n_1530),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1565),
.B(n_1516),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1566),
.B(n_1517),
.Y(n_1600)
);

INVxp67_ASAP7_75t_SL g1601 ( 
.A(n_1548),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1555),
.A2(n_1459),
.B1(n_1458),
.B2(n_1547),
.Y(n_1602)
);

CKINVDCx16_ASAP7_75t_R g1603 ( 
.A(n_1560),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1558),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1557),
.B(n_1375),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1580),
.B(n_1545),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1553),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1561),
.B(n_1563),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1567),
.B(n_1545),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1551),
.B(n_1524),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1587),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1551),
.B(n_1524),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1569),
.B(n_1559),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1576),
.B(n_1547),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1570),
.B(n_1529),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1582),
.B(n_1529),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1572),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1587),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1584),
.B(n_1531),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_SL g1620 ( 
.A(n_1585),
.B(n_1472),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1571),
.A2(n_1490),
.B1(n_1306),
.B2(n_1316),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1573),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1574),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1577),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1583),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1579),
.B(n_1465),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1586),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1579),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1575),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1578),
.A2(n_1458),
.B1(n_1472),
.B2(n_1503),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1571),
.B(n_1513),
.Y(n_1631)
);

AOI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1592),
.A2(n_1568),
.B1(n_1521),
.B2(n_1531),
.C(n_1535),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1607),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1604),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1614),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1590),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1589),
.B(n_1535),
.Y(n_1637)
);

NAND3xp33_ASAP7_75t_SL g1638 ( 
.A(n_1625),
.B(n_1397),
.C(n_1399),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1603),
.A2(n_1490),
.B1(n_1349),
.B2(n_1329),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1588),
.A2(n_1601),
.B1(n_1608),
.B2(n_1595),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1597),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1589),
.B(n_1536),
.Y(n_1642)
);

AOI222xp33_ASAP7_75t_L g1643 ( 
.A1(n_1610),
.A2(n_1485),
.B1(n_1476),
.B2(n_1521),
.C1(n_1444),
.C2(n_1536),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1627),
.B(n_1513),
.Y(n_1644)
);

OAI31xp33_ASAP7_75t_L g1645 ( 
.A1(n_1595),
.A2(n_1521),
.A3(n_1474),
.B(n_1468),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1628),
.B(n_1521),
.Y(n_1646)
);

O2A1O1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1601),
.A2(n_1612),
.B(n_1602),
.C(n_1605),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1614),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1608),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

OAI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1621),
.A2(n_1435),
.B1(n_1392),
.B2(n_1542),
.C(n_1540),
.Y(n_1651)
);

OAI32xp33_ASAP7_75t_L g1652 ( 
.A1(n_1629),
.A2(n_1475),
.A3(n_1468),
.B1(n_1503),
.B2(n_1493),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1631),
.B(n_1522),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1617),
.Y(n_1654)
);

OAI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1621),
.A2(n_1532),
.B1(n_1528),
.B2(n_1542),
.C(n_1540),
.Y(n_1655)
);

AND2x4_ASAP7_75t_SL g1656 ( 
.A(n_1626),
.B(n_1325),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1617),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1606),
.B(n_1522),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1591),
.B(n_1528),
.Y(n_1659)
);

AOI21xp33_ASAP7_75t_L g1660 ( 
.A1(n_1605),
.A2(n_1433),
.B(n_1427),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1594),
.B(n_1532),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_SL g1662 ( 
.A(n_1596),
.B(n_1351),
.C(n_1347),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1626),
.B(n_1485),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1619),
.B(n_1438),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1623),
.B(n_1534),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1618),
.Y(n_1666)
);

INVxp67_ASAP7_75t_SL g1667 ( 
.A(n_1618),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1635),
.B(n_1624),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1635),
.B(n_1598),
.Y(n_1669)
);

NAND3x1_ASAP7_75t_L g1670 ( 
.A(n_1640),
.B(n_1620),
.C(n_1609),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1648),
.B(n_1624),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1644),
.B(n_1622),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1648),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1649),
.B(n_1593),
.Y(n_1674)
);

O2A1O1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1649),
.A2(n_1630),
.B(n_1613),
.C(n_1622),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1634),
.B(n_1599),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1667),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1659),
.B(n_1600),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1662),
.A2(n_1616),
.B1(n_1490),
.B2(n_1615),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1633),
.B(n_1534),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1667),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1656),
.B(n_1546),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1666),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1654),
.B(n_1537),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1656),
.B(n_1537),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1646),
.B(n_1520),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1657),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1646),
.B(n_1520),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1637),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1663),
.B(n_1520),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1653),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1658),
.B(n_1546),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1636),
.B(n_1478),
.Y(n_1693)
);

INVxp33_ASAP7_75t_SL g1694 ( 
.A(n_1673),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1677),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1677),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1681),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1670),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1681),
.Y(n_1699)
);

BUFx12f_ASAP7_75t_L g1700 ( 
.A(n_1669),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1669),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1691),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1672),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1687),
.Y(n_1704)
);

NAND2x1_ASAP7_75t_SL g1705 ( 
.A(n_1674),
.B(n_1641),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1687),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1672),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1683),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1689),
.B(n_1647),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1683),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1671),
.B(n_1642),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1668),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1680),
.Y(n_1713)
);

NAND4xp25_ASAP7_75t_L g1714 ( 
.A(n_1709),
.B(n_1679),
.C(n_1675),
.D(n_1645),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1694),
.B(n_1676),
.Y(n_1715)
);

AND3x2_ASAP7_75t_L g1716 ( 
.A(n_1701),
.B(n_1685),
.C(n_1632),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1703),
.B(n_1678),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1694),
.B(n_1651),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1700),
.B(n_1660),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1698),
.B(n_1638),
.Y(n_1720)
);

O2A1O1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1698),
.A2(n_1661),
.B(n_1652),
.C(n_1655),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1707),
.B(n_1685),
.Y(n_1722)
);

NOR3xp33_ASAP7_75t_SL g1723 ( 
.A(n_1712),
.B(n_1670),
.C(n_1650),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1698),
.A2(n_1639),
.B1(n_1685),
.B2(n_1684),
.C(n_1688),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1700),
.B(n_1702),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1723),
.A2(n_1639),
.B1(n_1707),
.B2(n_1711),
.Y(n_1726)
);

OAI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1721),
.A2(n_1705),
.B1(n_1712),
.B2(n_1713),
.C(n_1697),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1722),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1717),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1720),
.Y(n_1730)
);

AO22x2_ASAP7_75t_L g1731 ( 
.A1(n_1715),
.A2(n_1695),
.B1(n_1696),
.B2(n_1699),
.Y(n_1731)
);

OAI211xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1725),
.A2(n_1695),
.B(n_1696),
.C(n_1699),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1718),
.B(n_1705),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1716),
.Y(n_1734)
);

INVxp33_ASAP7_75t_L g1735 ( 
.A(n_1719),
.Y(n_1735)
);

AOI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1714),
.A2(n_1708),
.B1(n_1706),
.B2(n_1704),
.C(n_1710),
.Y(n_1736)
);

OAI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1724),
.A2(n_1685),
.B(n_1643),
.Y(n_1737)
);

OAI31xp33_ASAP7_75t_L g1738 ( 
.A1(n_1727),
.A2(n_1682),
.A3(n_1688),
.B(n_1686),
.Y(n_1738)
);

NOR2xp67_ASAP7_75t_L g1739 ( 
.A(n_1729),
.B(n_1682),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1731),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1731),
.Y(n_1741)
);

NOR2xp67_ASAP7_75t_L g1742 ( 
.A(n_1728),
.B(n_1686),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1730),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1734),
.B(n_1692),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_R g1745 ( 
.A(n_1743),
.B(n_1733),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1739),
.B(n_1726),
.Y(n_1746)
);

NAND2xp33_ASAP7_75t_SL g1747 ( 
.A(n_1740),
.B(n_1735),
.Y(n_1747)
);

NAND2xp33_ASAP7_75t_SL g1748 ( 
.A(n_1741),
.B(n_1737),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_R g1749 ( 
.A(n_1744),
.B(n_1732),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1738),
.B(n_1736),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1742),
.B(n_1693),
.Y(n_1751)
);

AOI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1748),
.A2(n_1744),
.B1(n_1692),
.B2(n_1690),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1747),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1746),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1751),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1749),
.B(n_1690),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1745),
.Y(n_1757)
);

OAI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1752),
.A2(n_1750),
.B(n_1665),
.Y(n_1758)
);

XNOR2xp5_ASAP7_75t_L g1759 ( 
.A(n_1757),
.B(n_1664),
.Y(n_1759)
);

AO22x2_ASAP7_75t_L g1760 ( 
.A1(n_1753),
.A2(n_1359),
.B1(n_1363),
.B2(n_1546),
.Y(n_1760)
);

INVx2_ASAP7_75t_SL g1761 ( 
.A(n_1760),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1754),
.B1(n_1757),
.B2(n_1755),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1762),
.A2(n_1758),
.B(n_1756),
.Y(n_1763)
);

O2A1O1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1762),
.A2(n_1759),
.B(n_1503),
.C(n_1468),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1763),
.Y(n_1765)
);

INVx2_ASAP7_75t_SL g1766 ( 
.A(n_1764),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1765),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1766),
.Y(n_1768)
);

OAI221xp5_ASAP7_75t_R g1769 ( 
.A1(n_1767),
.A2(n_1323),
.B1(n_1368),
.B2(n_1325),
.C(n_1324),
.Y(n_1769)
);

AOI211xp5_ASAP7_75t_L g1770 ( 
.A1(n_1769),
.A2(n_1768),
.B(n_1324),
.C(n_1395),
.Y(n_1770)
);


endmodule