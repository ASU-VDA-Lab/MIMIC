module fake_jpeg_21869_n_282 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_282);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_24),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_26),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_34),
.B1(n_27),
.B2(n_25),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_50),
.B(n_58),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_34),
.B1(n_28),
.B2(n_27),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_41),
.C(n_37),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_34),
.B1(n_27),
.B2(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_56),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_20),
.B1(n_28),
.B2(n_19),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_53),
.A2(n_41),
.B1(n_37),
.B2(n_31),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_20),
.B1(n_23),
.B2(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_29),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_60),
.A2(n_18),
.B1(n_21),
.B2(n_17),
.Y(n_97)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVxp67_ASAP7_75t_SL g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_64),
.B(n_83),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_43),
.B1(n_26),
.B2(n_39),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_67),
.A2(n_46),
.B1(n_56),
.B2(n_51),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_72),
.Y(n_100)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_76),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_41),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_90),
.Y(n_113)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_82),
.Y(n_119)
);

CKINVDCx12_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_36),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_89),
.Y(n_117)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_48),
.B(n_35),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_85),
.B(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_29),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_91),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_36),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_41),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_58),
.B(n_41),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_67),
.CI(n_81),
.CON(n_109),
.SN(n_109)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_49),
.B(n_18),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_10),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_37),
.B1(n_61),
.B2(n_46),
.Y(n_106)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_98),
.B1(n_30),
.B2(n_56),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_49),
.A2(n_21),
.B1(n_30),
.B2(n_31),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_37),
.C(n_41),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_89),
.C(n_87),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_50),
.B1(n_45),
.B2(n_51),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_101),
.A2(n_103),
.B1(n_115),
.B2(n_79),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_116),
.B1(n_96),
.B2(n_71),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_76),
.B(n_64),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_68),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_84),
.A2(n_44),
.B1(n_37),
.B2(n_61),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_32),
.B1(n_61),
.B2(n_43),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_26),
.B1(n_32),
.B2(n_36),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_118),
.A2(n_65),
.B1(n_88),
.B2(n_72),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_74),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_70),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_36),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_70),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_128),
.B(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_131),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_12),
.Y(n_179)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_133),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_155),
.C(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_66),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_126),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_144),
.B1(n_103),
.B2(n_124),
.Y(n_172)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_142),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_92),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_143),
.A2(n_149),
.B(n_156),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_147),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_115),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_83),
.Y(n_148)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_107),
.B1(n_122),
.B2(n_118),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_90),
.Y(n_153)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_112),
.B(n_90),
.Y(n_154)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_73),
.C(n_80),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_32),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_69),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_172),
.B1(n_180),
.B2(n_181),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_155),
.C(n_143),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_122),
.B(n_109),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_175),
.B(n_178),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_152),
.A2(n_101),
.B1(n_109),
.B2(n_99),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_167),
.A2(n_174),
.B1(n_168),
.B2(n_134),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_179),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_99),
.B1(n_95),
.B2(n_78),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_114),
.B(n_104),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_104),
.B(n_108),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_124),
.B1(n_96),
.B2(n_91),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_128),
.A2(n_82),
.B1(n_111),
.B2(n_69),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_197),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_189),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_194),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_203),
.B1(n_206),
.B2(n_174),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_140),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_196),
.C(n_199),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_145),
.C(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

OAI22x1_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_143),
.B1(n_150),
.B2(n_156),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_202),
.B1(n_184),
.B2(n_176),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_138),
.C(n_146),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_131),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_201),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_149),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_129),
.B(n_135),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_136),
.B1(n_111),
.B2(n_1),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_159),
.B(n_9),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_205),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_9),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_9),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_167),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_212),
.B1(n_219),
.B2(n_226),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_178),
.B(n_175),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_221),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_166),
.B1(n_170),
.B2(n_184),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_200),
.B(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_217),
.A2(n_224),
.B1(n_187),
.B2(n_190),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_191),
.B(n_170),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_226),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_166),
.B1(n_158),
.B2(n_173),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_203),
.C(n_186),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_185),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_179),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_10),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_173),
.B1(n_183),
.B2(n_1),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_202),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_195),
.C(n_196),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_229),
.C(n_230),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_199),
.C(n_207),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_187),
.C(n_188),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_237),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_16),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

BUFx12_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_2),
.C(n_4),
.Y(n_238)
);

NOR2xp67_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_4),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_239),
.B(n_240),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_16),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_225),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_235),
.A2(n_217),
.B1(n_215),
.B2(n_222),
.Y(n_242)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_236),
.A2(n_209),
.B1(n_213),
.B2(n_211),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_251),
.B1(n_5),
.B2(n_7),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_236),
.B(n_233),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_247),
.B(n_229),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_215),
.B1(n_222),
.B2(n_210),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_238),
.A2(n_223),
.B1(n_225),
.B2(n_7),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_234),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_259),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_228),
.C(n_237),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_257),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_234),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_258),
.B(n_262),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_5),
.B(n_6),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_262),
.B1(n_251),
.B2(n_247),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_8),
.C(n_10),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_244),
.B1(n_242),
.B2(n_252),
.Y(n_263)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_243),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_267),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_261),
.B(n_248),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_265),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_243),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_272),
.Y(n_276)
);

AOI21x1_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_254),
.B(n_12),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_266),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_11),
.B1(n_15),
.B2(n_276),
.Y(n_279)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_270),
.A2(n_264),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_16),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_273),
.C(n_14),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_279),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_15),
.Y(n_282)
);


endmodule