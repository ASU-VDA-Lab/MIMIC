module fake_netlist_1_348_n_1081 (n_120, n_136, n_260, n_155, n_107, n_103, n_157, n_52, n_162, n_114, n_156, n_154, n_50, n_7, n_239, n_222, n_253, n_3, n_34, n_142, n_273, n_231, n_25, n_9, n_163, n_96, n_204, n_72, n_77, n_90, n_169, n_178, n_214, n_227, n_180, n_250, n_99, n_43, n_73, n_190, n_62, n_167, n_97, n_229, n_133, n_199, n_268, n_33, n_192, n_4, n_59, n_76, n_6, n_74, n_8, n_61, n_44, n_189, n_216, n_153, n_187, n_226, n_66, n_88, n_46, n_121, n_174, n_240, n_188, n_108, n_161, n_37, n_122, n_165, n_224, n_18, n_247, n_65, n_87, n_207, n_5, n_197, n_81, n_211, n_85, n_112, n_215, n_264, n_102, n_172, n_47, n_109, n_198, n_1, n_201, n_16, n_78, n_95, n_217, n_40, n_68, n_105, n_210, n_251, n_36, n_228, n_259, n_11, n_244, n_115, n_270, n_225, n_179, n_208, n_237, n_252, n_15, n_168, n_271, n_139, n_152, n_151, n_71, n_117, n_238, n_176, n_70, n_256, n_94, n_2, n_194, n_17, n_221, n_58, n_195, n_113, n_242, n_209, n_241, n_20, n_84, n_130, n_266, n_12, n_56, n_80, n_223, n_67, n_116, n_22, n_118, n_19, n_233, n_257, n_202, n_26, n_203, n_261, n_274, n_243, n_39, n_101, n_98, n_150, n_220, n_235, n_38, n_230, n_245, n_104, n_272, n_100, n_159, n_24, n_141, n_35, n_91, n_146, n_160, n_32, n_148, n_149, n_246, n_263, n_93, n_191, n_143, n_134, n_48, n_63, n_255, n_54, n_193, n_232, n_125, n_41, n_147, n_55, n_145, n_185, n_29, n_166, n_218, n_267, n_173, n_181, n_123, n_171, n_219, n_60, n_135, n_138, n_140, n_111, n_10, n_212, n_30, n_13, n_254, n_92, n_75, n_82, n_53, n_183, n_64, n_132, n_69, n_196, n_213, n_175, n_248, n_127, n_128, n_170, n_83, n_200, n_158, n_205, n_23, n_0, n_126, n_258, n_110, n_249, n_262, n_234, n_184, n_182, n_269, n_119, n_265, n_57, n_51, n_144, n_106, n_186, n_45, n_42, n_21, n_137, n_236, n_131, n_86, n_27, n_124, n_89, n_177, n_28, n_79, n_129, n_164, n_49, n_206, n_14, n_31, n_1081, n_1082);
input n_120;
input n_136;
input n_260;
input n_155;
input n_107;
input n_103;
input n_157;
input n_52;
input n_162;
input n_114;
input n_156;
input n_154;
input n_50;
input n_7;
input n_239;
input n_222;
input n_253;
input n_3;
input n_34;
input n_142;
input n_273;
input n_231;
input n_25;
input n_9;
input n_163;
input n_96;
input n_204;
input n_72;
input n_77;
input n_90;
input n_169;
input n_178;
input n_214;
input n_227;
input n_180;
input n_250;
input n_99;
input n_43;
input n_73;
input n_190;
input n_62;
input n_167;
input n_97;
input n_229;
input n_133;
input n_199;
input n_268;
input n_33;
input n_192;
input n_4;
input n_59;
input n_76;
input n_6;
input n_74;
input n_8;
input n_61;
input n_44;
input n_189;
input n_216;
input n_153;
input n_187;
input n_226;
input n_66;
input n_88;
input n_46;
input n_121;
input n_174;
input n_240;
input n_188;
input n_108;
input n_161;
input n_37;
input n_122;
input n_165;
input n_224;
input n_18;
input n_247;
input n_65;
input n_87;
input n_207;
input n_5;
input n_197;
input n_81;
input n_211;
input n_85;
input n_112;
input n_215;
input n_264;
input n_102;
input n_172;
input n_47;
input n_109;
input n_198;
input n_1;
input n_201;
input n_16;
input n_78;
input n_95;
input n_217;
input n_40;
input n_68;
input n_105;
input n_210;
input n_251;
input n_36;
input n_228;
input n_259;
input n_11;
input n_244;
input n_115;
input n_270;
input n_225;
input n_179;
input n_208;
input n_237;
input n_252;
input n_15;
input n_168;
input n_271;
input n_139;
input n_152;
input n_151;
input n_71;
input n_117;
input n_238;
input n_176;
input n_70;
input n_256;
input n_94;
input n_2;
input n_194;
input n_17;
input n_221;
input n_58;
input n_195;
input n_113;
input n_242;
input n_209;
input n_241;
input n_20;
input n_84;
input n_130;
input n_266;
input n_12;
input n_56;
input n_80;
input n_223;
input n_67;
input n_116;
input n_22;
input n_118;
input n_19;
input n_233;
input n_257;
input n_202;
input n_26;
input n_203;
input n_261;
input n_274;
input n_243;
input n_39;
input n_101;
input n_98;
input n_150;
input n_220;
input n_235;
input n_38;
input n_230;
input n_245;
input n_104;
input n_272;
input n_100;
input n_159;
input n_24;
input n_141;
input n_35;
input n_91;
input n_146;
input n_160;
input n_32;
input n_148;
input n_149;
input n_246;
input n_263;
input n_93;
input n_191;
input n_143;
input n_134;
input n_48;
input n_63;
input n_255;
input n_54;
input n_193;
input n_232;
input n_125;
input n_41;
input n_147;
input n_55;
input n_145;
input n_185;
input n_29;
input n_166;
input n_218;
input n_267;
input n_173;
input n_181;
input n_123;
input n_171;
input n_219;
input n_60;
input n_135;
input n_138;
input n_140;
input n_111;
input n_10;
input n_212;
input n_30;
input n_13;
input n_254;
input n_92;
input n_75;
input n_82;
input n_53;
input n_183;
input n_64;
input n_132;
input n_69;
input n_196;
input n_213;
input n_175;
input n_248;
input n_127;
input n_128;
input n_170;
input n_83;
input n_200;
input n_158;
input n_205;
input n_23;
input n_0;
input n_126;
input n_258;
input n_110;
input n_249;
input n_262;
input n_234;
input n_184;
input n_182;
input n_269;
input n_119;
input n_265;
input n_57;
input n_51;
input n_144;
input n_106;
input n_186;
input n_45;
input n_42;
input n_21;
input n_137;
input n_236;
input n_131;
input n_86;
input n_27;
input n_124;
input n_89;
input n_177;
input n_28;
input n_79;
input n_129;
input n_164;
input n_49;
input n_206;
input n_14;
input n_31;
output n_1081;
output n_1082;
wire n_890;
wire n_107;
wire n_646;
wire n_759;
wire n_987;
wire n_658;
wire n_673;
wire n_156;
wire n_154;
wire n_239;
wire n_7;
wire n_309;
wire n_944;
wire n_356;
wire n_895;
wire n_1029;
wire n_327;
wire n_25;
wire n_1014;
wire n_994;
wire n_204;
wire n_592;
wire n_769;
wire n_929;
wire n_1041;
wire n_370;
wire n_384;
wire n_439;
wire n_545;
wire n_169;
wire n_959;
wire n_180;
wire n_604;
wire n_1015;
wire n_99;
wire n_43;
wire n_73;
wire n_440;
wire n_199;
wire n_279;
wire n_786;
wire n_831;
wire n_357;
wire n_74;
wire n_729;
wire n_308;
wire n_518;
wire n_394;
wire n_44;
wire n_189;
wire n_681;
wire n_226;
wire n_447;
wire n_352;
wire n_66;
wire n_379;
wire n_903;
wire n_535;
wire n_689;
wire n_886;
wire n_595;
wire n_875;
wire n_626;
wire n_316;
wire n_285;
wire n_952;
wire n_564;
wire n_586;
wire n_1047;
wire n_471;
wire n_47;
wire n_766;
wire n_1049;
wire n_475;
wire n_744;
wire n_949;
wire n_850;
wire n_281;
wire n_645;
wire n_497;
wire n_399;
wire n_11;
wire n_1035;
wire n_942;
wire n_295;
wire n_371;
wire n_579;
wire n_516;
wire n_608;
wire n_368;
wire n_805;
wire n_373;
wire n_1020;
wire n_139;
wire n_342;
wire n_151;
wire n_71;
wire n_288;
wire n_557;
wire n_753;
wire n_176;
wire n_859;
wire n_436;
wire n_438;
wire n_900;
wire n_869;
wire n_935;
wire n_931;
wire n_359;
wire n_195;
wire n_300;
wire n_487;
wire n_461;
wire n_723;
wire n_223;
wire n_833;
wire n_405;
wire n_830;
wire n_562;
wire n_19;
wire n_409;
wire n_971;
wire n_482;
wire n_838;
wire n_967;
wire n_1050;
wire n_534;
wire n_569;
wire n_707;
wire n_526;
wire n_261;
wire n_423;
wire n_483;
wire n_220;
wire n_353;
wire n_410;
wire n_104;
wire n_709;
wire n_303;
wire n_502;
wire n_821;
wire n_468;
wire n_159;
wire n_566;
wire n_91;
wire n_301;
wire n_340;
wire n_963;
wire n_148;
wire n_149;
wire n_567;
wire n_378;
wire n_752;
wire n_246;
wire n_676;
wire n_823;
wire n_191;
wire n_143;
wire n_780;
wire n_864;
wire n_629;
wire n_446;
wire n_63;
wire n_402;
wire n_54;
wire n_876;
wire n_387;
wire n_125;
wire n_145;
wire n_961;
wire n_166;
wire n_558;
wire n_596;
wire n_1046;
wire n_492;
wire n_181;
wire n_123;
wire n_219;
wire n_494;
wire n_553;
wire n_555;
wire n_343;
wire n_1059;
wire n_135;
wire n_481;
wire n_621;
wire n_817;
wire n_776;
wire n_315;
wire n_397;
wire n_53;
wire n_880;
wire n_981;
wire n_213;
wire n_196;
wire n_293;
wire n_797;
wire n_836;
wire n_127;
wire n_312;
wire n_1058;
wire n_1045;
wire n_742;
wire n_424;
wire n_23;
wire n_110;
wire n_1028;
wire n_990;
wire n_1048;
wire n_663;
wire n_269;
wire n_182;
wire n_1019;
wire n_529;
wire n_656;
wire n_751;
wire n_887;
wire n_186;
wire n_137;
wire n_507;
wire n_334;
wire n_1062;
wire n_993;
wire n_164;
wire n_1024;
wire n_433;
wire n_660;
wire n_120;
wire n_392;
wire n_650;
wire n_806;
wire n_155;
wire n_1053;
wire n_162;
wire n_114;
wire n_977;
wire n_772;
wire n_50;
wire n_816;
wire n_789;
wire n_3;
wire n_331;
wire n_651;
wire n_574;
wire n_882;
wire n_999;
wire n_636;
wire n_330;
wire n_614;
wire n_231;
wire n_884;
wire n_9;
wire n_737;
wire n_428;
wire n_178;
wire n_478;
wire n_814;
wire n_652;
wire n_678;
wire n_708;
wire n_229;
wire n_97;
wire n_982;
wire n_133;
wire n_442;
wire n_324;
wire n_991;
wire n_422;
wire n_192;
wire n_699;
wire n_857;
wire n_329;
wire n_6;
wire n_8;
wire n_998;
wire n_578;
wire n_928;
wire n_883;
wire n_187;
wire n_548;
wire n_188;
wire n_443;
wire n_304;
wire n_18;
wire n_682;
wire n_801;
wire n_441;
wire n_868;
wire n_628;
wire n_425;
wire n_920;
wire n_912;
wire n_314;
wire n_824;
wire n_601;
wire n_307;
wire n_517;
wire n_215;
wire n_736;
wire n_172;
wire n_905;
wire n_109;
wire n_332;
wire n_198;
wire n_386;
wire n_934;
wire n_653;
wire n_351;
wire n_1;
wire n_979;
wire n_670;
wire n_16;
wire n_95;
wire n_40;
wire n_210;
wire n_426;
wire n_755;
wire n_716;
wire n_228;
wire n_863;
wire n_671;
wire n_892;
wire n_278;
wire n_115;
wire n_270;
wire n_476;
wire n_989;
wire n_765;
wire n_829;
wire n_599;
wire n_715;
wire n_849;
wire n_1077;
wire n_984;
wire n_404;
wire n_289;
wire n_179;
wire n_366;
wire n_721;
wire n_362;
wire n_617;
wire n_688;
wire n_837;
wire n_485;
wire n_396;
wire n_549;
wire n_354;
wire n_720;
wire n_152;
wire n_851;
wire n_980;
wire n_70;
wire n_588;
wire n_458;
wire n_375;
wire n_855;
wire n_17;
wire n_322;
wire n_911;
wire n_506;
wire n_317;
wire n_328;
wire n_711;
wire n_221;
wire n_491;
wire n_800;
wire n_973;
wire n_388;
wire n_773;
wire n_266;
wire n_763;
wire n_80;
wire n_632;
wire n_793;
wire n_906;
wire n_679;
wire n_522;
wire n_1055;
wire n_546;
wire n_615;
wire n_684;
wire n_701;
wire n_326;
wire n_532;
wire n_756;
wire n_635;
wire n_544;
wire n_888;
wire n_879;
wire n_576;
wire n_992;
wire n_275;
wire n_691;
wire n_622;
wire n_661;
wire n_909;
wire n_493;
wire n_274;
wire n_910;
wire n_972;
wire n_235;
wire n_150;
wire n_690;
wire n_38;
wire n_533;
wire n_272;
wire n_686;
wire n_965;
wire n_299;
wire n_100;
wire n_561;
wire n_1023;
wire n_1057;
wire n_1072;
wire n_581;
wire n_280;
wire n_141;
wire n_1068;
wire n_509;
wire n_160;
wire n_499;
wire n_377;
wire n_1043;
wire n_1044;
wire n_263;
wire n_757;
wire n_844;
wire n_1013;
wire n_1060;
wire n_695;
wire n_193;
wire n_232;
wire n_344;
wire n_878;
wire n_783;
wire n_812;
wire n_147;
wire n_1065;
wire n_185;
wire n_367;
wire n_955;
wire n_795;
wire n_267;
wire n_1007;
wire n_687;
wire n_950;
wire n_638;
wire n_171;
wire n_873;
wire n_899;
wire n_450;
wire n_585;
wire n_644;
wire n_140;
wire n_111;
wire n_746;
wire n_212;
wire n_779;
wire n_978;
wire n_1064;
wire n_30;
wire n_634;
wire n_13;
wire n_254;
wire n_559;
wire n_728;
wire n_435;
wire n_704;
wire n_583;
wire n_841;
wire n_64;
wire n_69;
wire n_248;
wire n_866;
wire n_407;
wire n_970;
wire n_527;
wire n_1021;
wire n_83;
wire n_200;
wire n_603;
wire n_986;
wire n_262;
wire n_1032;
wire n_921;
wire n_119;
wire n_667;
wire n_503;
wire n_969;
wire n_856;
wire n_1076;
wire n_1081;
wire n_927;
wire n_1012;
wire n_339;
wire n_347;
wire n_124;
wire n_696;
wire n_748;
wire n_1018;
wire n_79;
wire n_129;
wire n_904;
wire n_611;
wire n_1016;
wire n_521;
wire n_157;
wire n_774;
wire n_103;
wire n_808;
wire n_421;
wire n_1080;
wire n_52;
wire n_253;
wire n_1038;
wire n_434;
wire n_677;
wire n_624;
wire n_273;
wire n_325;
wire n_571;
wire n_524;
wire n_692;
wire n_530;
wire n_743;
wire n_951;
wire n_163;
wire n_348;
wire n_96;
wire n_669;
wire n_685;
wire n_90;
wire n_72;
wire n_77;
wire n_594;
wire n_762;
wire n_740;
wire n_214;
wire n_787;
wire n_1030;
wire n_1074;
wire n_770;
wire n_167;
wire n_861;
wire n_809;
wire n_364;
wire n_33;
wire n_908;
wire n_464;
wire n_76;
wire n_470;
wire n_590;
wire n_61;
wire n_1022;
wire n_463;
wire n_216;
wire n_609;
wire n_355;
wire n_153;
wire n_946;
wire n_1066;
wire n_121;
wire n_286;
wire n_408;
wire n_1003;
wire n_247;
wire n_484;
wire n_224;
wire n_161;
wire n_431;
wire n_165;
wire n_860;
wire n_413;
wire n_65;
wire n_537;
wire n_710;
wire n_525;
wire n_560;
wire n_5;
wire n_496;
wire n_393;
wire n_843;
wire n_211;
wire n_85;
wire n_320;
wire n_264;
wire n_102;
wire n_283;
wire n_733;
wire n_846;
wire n_290;
wire n_217;
wire n_201;
wire n_1031;
wire n_791;
wire n_792;
wire n_277;
wire n_932;
wire n_259;
wire n_885;
wire n_612;
wire n_244;
wire n_666;
wire n_771;
wire n_827;
wire n_1061;
wire n_276;
wire n_297;
wire n_225;
wire n_1037;
wire n_631;
wire n_350;
wire n_747;
wire n_616;
wire n_208;
wire n_815;
wire n_523;
wire n_854;
wire n_901;
wire n_528;
wire n_419;
wire n_985;
wire n_252;
wire n_922;
wire n_519;
wire n_168;
wire n_839;
wire n_271;
wire n_966;
wire n_693;
wire n_1011;
wire n_785;
wire n_896;
wire n_739;
wire n_1056;
wire n_94;
wire n_997;
wire n_194;
wire n_858;
wire n_758;
wire n_825;
wire n_282;
wire n_58;
wire n_775;
wire n_113;
wire n_242;
wire n_498;
wire n_501;
wire n_284;
wire n_538;
wire n_302;
wire n_321;
wire n_703;
wire n_811;
wire n_116;
wire n_734;
wire n_292;
wire n_547;
wire n_593;
wire n_118;
wire n_587;
wire n_233;
wire n_554;
wire n_597;
wire n_741;
wire n_705;
wire n_257;
wire n_698;
wire n_828;
wire n_722;
wire n_988;
wire n_26;
wire n_203;
wire n_477;
wire n_996;
wire n_460;
wire n_243;
wire n_318;
wire n_346;
wire n_98;
wire n_345;
wire n_230;
wire n_452;
wire n_714;
wire n_146;
wire n_337;
wire n_32;
wire n_637;
wire n_641;
wire n_726;
wire n_531;
wire n_957;
wire n_872;
wire n_93;
wire n_539;
wire n_847;
wire n_406;
wire n_372;
wire n_842;
wire n_820;
wire n_713;
wire n_467;
wire n_923;
wire n_702;
wire n_41;
wire n_760;
wire n_826;
wire n_918;
wire n_1009;
wire n_623;
wire n_417;
wire n_451;
wire n_665;
wire n_898;
wire n_647;
wire n_445;
wire n_500;
wire n_948;
wire n_732;
wire n_926;
wire n_1026;
wire n_845;
wire n_575;
wire n_390;
wire n_600;
wire n_10;
wire n_1001;
wire n_1036;
wire n_818;
wire n_75;
wire n_82;
wire n_183;
wire n_731;
wire n_550;
wire n_132;
wire n_643;
wire n_761;
wire n_1006;
wire n_778;
wire n_582;
wire n_784;
wire n_170;
wire n_925;
wire n_1075;
wire n_205;
wire n_158;
wire n_915;
wire n_126;
wire n_473;
wire n_249;
wire n_389;
wire n_834;
wire n_510;
wire n_360;
wire n_363;
wire n_749;
wire n_1069;
wire n_427;
wire n_1078;
wire n_724;
wire n_1040;
wire n_1067;
wire n_106;
wire n_296;
wire n_605;
wire n_42;
wire n_21;
wire n_835;
wire n_437;
wire n_871;
wire n_620;
wire n_975;
wire n_89;
wire n_480;
wire n_1073;
wire n_1039;
wire n_939;
wire n_940;
wire n_130;
wire n_310;
wire n_341;
wire n_700;
wire n_640;
wire n_14;
wire n_236;
wire n_639;
wire n_1033;
wire n_727;
wire n_260;
wire n_136;
wire n_891;
wire n_1004;
wire n_1002;
wire n_580;
wire n_976;
wire n_610;
wire n_938;
wire n_1008;
wire n_222;
wire n_657;
wire n_822;
wire n_381;
wire n_964;
wire n_34;
wire n_142;
wire n_853;
wire n_754;
wire n_385;
wire n_798;
wire n_227;
wire n_395;
wire n_454;
wire n_943;
wire n_453;
wire n_250;
wire n_551;
wire n_268;
wire n_190;
wire n_606;
wire n_62;
wire n_712;
wire n_777;
wire n_4;
wire n_565;
wire n_323;
wire n_59;
wire n_956;
wire n_781;
wire n_954;
wire n_914;
wire n_1071;
wire n_945;
wire n_852;
wire n_376;
wire n_902;
wire n_694;
wire n_459;
wire n_768;
wire n_240;
wire n_568;
wire n_88;
wire n_46;
wire n_174;
wire n_717;
wire n_807;
wire n_108;
wire n_335;
wire n_37;
wire n_122;
wire n_374;
wire n_613;
wire n_380;
wire n_515;
wire n_802;
wire n_865;
wire n_1042;
wire n_672;
wire n_867;
wire n_466;
wire n_87;
wire n_349;
wire n_207;
wire n_1027;
wire n_197;
wire n_541;
wire n_572;
wire n_81;
wire n_298;
wire n_112;
wire n_630;
wire n_735;
wire n_649;
wire n_983;
wire n_1052;
wire n_602;
wire n_78;
wire n_552;
wire n_68;
wire n_919;
wire n_444;
wire n_105;
wire n_598;
wire n_251;
wire n_810;
wire n_416;
wire n_36;
wire n_962;
wire n_916;
wire n_889;
wire n_870;
wire n_432;
wire n_913;
wire n_917;
wire n_465;
wire n_414;
wire n_680;
wire n_730;
wire n_369;
wire n_469;
wire n_361;
wire n_767;
wire n_237;
wire n_1034;
wire n_881;
wire n_654;
wire n_520;
wire n_633;
wire n_15;
wire n_429;
wire n_803;
wire n_960;
wire n_398;
wire n_668;
wire n_256;
wire n_117;
wire n_238;
wire n_365;
wire n_577;
wire n_796;
wire n_804;
wire n_294;
wire n_2;
wire n_338;
wire n_662;
wire n_907;
wire n_591;
wire n_391;
wire n_1025;
wire n_209;
wire n_241;
wire n_874;
wire n_84;
wire n_20;
wire n_782;
wire n_449;
wire n_832;
wire n_1070;
wire n_412;
wire n_12;
wire n_618;
wire n_455;
wire n_504;
wire n_56;
wire n_67;
wire n_790;
wire n_456;
wire n_22;
wire n_683;
wire n_479;
wire n_584;
wire n_311;
wire n_401;
wire n_877;
wire n_383;
wire n_813;
wire n_202;
wire n_319;
wire n_542;
wire n_725;
wire n_819;
wire n_862;
wire n_930;
wire n_39;
wire n_101;
wire n_953;
wire n_941;
wire n_1063;
wire n_291;
wire n_489;
wire n_245;
wire n_664;
wire n_933;
wire n_508;
wire n_764;
wire n_719;
wire n_486;
wire n_788;
wire n_24;
wire n_35;
wire n_655;
wire n_472;
wire n_490;
wire n_540;
wire n_947;
wire n_840;
wire n_1010;
wire n_400;
wire n_794;
wire n_457;
wire n_659;
wire n_134;
wire n_48;
wire n_255;
wire n_968;
wire n_563;
wire n_1017;
wire n_513;
wire n_55;
wire n_718;
wire n_543;
wire n_336;
wire n_29;
wire n_218;
wire n_893;
wire n_173;
wire n_488;
wire n_556;
wire n_648;
wire n_382;
wire n_799;
wire n_894;
wire n_138;
wire n_60;
wire n_936;
wire n_937;
wire n_462;
wire n_536;
wire n_573;
wire n_474;
wire n_924;
wire n_745;
wire n_305;
wire n_505;
wire n_430;
wire n_418;
wire n_495;
wire n_92;
wire n_313;
wire n_333;
wire n_358;
wire n_627;
wire n_750;
wire n_706;
wire n_589;
wire n_175;
wire n_897;
wire n_128;
wire n_306;
wire n_31;
wire n_697;
wire n_958;
wire n_0;
wire n_512;
wire n_675;
wire n_619;
wire n_642;
wire n_258;
wire n_974;
wire n_234;
wire n_607;
wire n_848;
wire n_184;
wire n_1000;
wire n_1005;
wire n_265;
wire n_57;
wire n_674;
wire n_51;
wire n_570;
wire n_411;
wire n_514;
wire n_287;
wire n_625;
wire n_403;
wire n_144;
wire n_995;
wire n_45;
wire n_420;
wire n_131;
wire n_86;
wire n_27;
wire n_738;
wire n_177;
wire n_28;
wire n_511;
wire n_1054;
wire n_448;
wire n_49;
wire n_206;
wire n_1051;
wire n_415;
CKINVDCx16_ASAP7_75t_R g275 ( .A(n_254), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_246), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_18), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_200), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_18), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_211), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_191), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_247), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_34), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_228), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_238), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_235), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_86), .Y(n_287) );
BUFx2_ASAP7_75t_SL g288 ( .A(n_17), .Y(n_288) );
INVxp33_ASAP7_75t_SL g289 ( .A(n_99), .Y(n_289) );
INVxp33_ASAP7_75t_SL g290 ( .A(n_255), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_23), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_248), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_231), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_212), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_257), .Y(n_295) );
INVxp33_ASAP7_75t_SL g296 ( .A(n_38), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_236), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g298 ( .A(n_180), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_250), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_46), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_227), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_165), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_259), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_201), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_69), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_123), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_119), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_156), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_135), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_125), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_137), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_26), .Y(n_312) );
CKINVDCx14_ASAP7_75t_R g313 ( .A(n_159), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_224), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_166), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_55), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_132), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_142), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_242), .Y(n_319) );
CKINVDCx16_ASAP7_75t_R g320 ( .A(n_103), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_207), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_203), .Y(n_322) );
BUFx10_ASAP7_75t_L g323 ( .A(n_109), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_215), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_190), .Y(n_325) );
INVxp33_ASAP7_75t_SL g326 ( .A(n_168), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_110), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_139), .Y(n_328) );
INVx1_ASAP7_75t_SL g329 ( .A(n_155), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_233), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_91), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_204), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_84), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_198), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_197), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_225), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_53), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g338 ( .A(n_244), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_85), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_63), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_243), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_92), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_219), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_210), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_138), .Y(n_345) );
INVxp67_ASAP7_75t_SL g346 ( .A(n_7), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_267), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_175), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_196), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_188), .Y(n_350) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_6), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_264), .Y(n_352) );
INVxp67_ASAP7_75t_L g353 ( .A(n_70), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_65), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_265), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_193), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_273), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_27), .Y(n_358) );
INVxp33_ASAP7_75t_SL g359 ( .A(n_32), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_245), .Y(n_360) );
INVxp33_ASAP7_75t_L g361 ( .A(n_13), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_90), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_41), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_216), .B(n_237), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_114), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_220), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_91), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_40), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_19), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_61), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_167), .Y(n_371) );
INVx2_ASAP7_75t_SL g372 ( .A(n_234), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_161), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_145), .B(n_19), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_120), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_66), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_111), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_232), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_45), .B(n_32), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_158), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_152), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_108), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_173), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_151), .Y(n_384) );
INVxp33_ASAP7_75t_L g385 ( .A(n_226), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_41), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_206), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_101), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_9), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_112), .Y(n_390) );
BUFx2_ASAP7_75t_L g391 ( .A(n_178), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_160), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_129), .Y(n_393) );
CKINVDCx16_ASAP7_75t_R g394 ( .A(n_72), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_54), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_28), .Y(n_396) );
CKINVDCx14_ASAP7_75t_R g397 ( .A(n_28), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_146), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_202), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_58), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_260), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_5), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_107), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_83), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_157), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_127), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_77), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_133), .Y(n_408) );
NOR2xp67_ASAP7_75t_L g409 ( .A(n_274), .B(n_205), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_266), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_71), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_23), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_162), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_268), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_116), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_189), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_136), .Y(n_417) );
INVxp33_ASAP7_75t_SL g418 ( .A(n_40), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_263), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_163), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_128), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_64), .Y(n_422) );
INVx3_ASAP7_75t_L g423 ( .A(n_411), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_282), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_411), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_282), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_315), .B(n_0), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_282), .Y(n_429) );
OA21x2_ASAP7_75t_L g430 ( .A1(n_276), .A2(n_94), .B(n_93), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_282), .Y(n_431) );
AND2x2_ASAP7_75t_SL g432 ( .A(n_383), .B(n_95), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_362), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_391), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_361), .B(n_0), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_278), .Y(n_436) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_278), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_407), .B(n_1), .Y(n_438) );
CKINVDCx8_ASAP7_75t_R g439 ( .A(n_275), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_323), .Y(n_440) );
INVx4_ASAP7_75t_L g441 ( .A(n_323), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_361), .B(n_1), .Y(n_442) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_285), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_372), .B(n_2), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_323), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_407), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_369), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_369), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_376), .Y(n_449) );
NOR2xp33_ASAP7_75t_SL g450 ( .A(n_320), .B(n_272), .Y(n_450) );
AND2x6_ASAP7_75t_L g451 ( .A(n_285), .B(n_96), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_276), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_284), .B(n_2), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_386), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_394), .Y(n_455) );
OAI21x1_ASAP7_75t_L g456 ( .A1(n_307), .A2(n_98), .B(n_97), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_429), .Y(n_457) );
BUFx8_ASAP7_75t_SL g458 ( .A(n_455), .Y(n_458) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_429), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_452), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_452), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_428), .B(n_353), .Y(n_462) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_429), .Y(n_463) );
INVx4_ASAP7_75t_L g464 ( .A(n_451), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_434), .B(n_441), .Y(n_465) );
INVx4_ASAP7_75t_L g466 ( .A(n_451), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_441), .B(n_385), .Y(n_467) );
AND2x2_ASAP7_75t_SL g468 ( .A(n_432), .B(n_450), .Y(n_468) );
BUFx3_ASAP7_75t_L g469 ( .A(n_451), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_429), .Y(n_470) );
BUFx3_ASAP7_75t_L g471 ( .A(n_451), .Y(n_471) );
NAND2xp33_ASAP7_75t_L g472 ( .A(n_451), .B(n_281), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_438), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_446), .B(n_313), .Y(n_474) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_429), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_429), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_440), .B(n_297), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_438), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_432), .A2(n_359), .B1(n_418), .B2(n_296), .Y(n_479) );
NAND2xp33_ASAP7_75t_L g480 ( .A(n_451), .B(n_293), .Y(n_480) );
INVx4_ASAP7_75t_SL g481 ( .A(n_451), .Y(n_481) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_435), .Y(n_482) );
INVx8_ASAP7_75t_L g483 ( .A(n_451), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_432), .A2(n_418), .B1(n_359), .B2(n_295), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_423), .B(n_376), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_434), .B(n_392), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_482), .Y(n_487) );
AND2x6_ASAP7_75t_SL g488 ( .A(n_458), .B(n_435), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_485), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_485), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_485), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_465), .B(n_440), .Y(n_492) );
INVx3_ASAP7_75t_L g493 ( .A(n_485), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_460), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_461), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_468), .A2(n_442), .B1(n_450), .B2(n_445), .Y(n_496) );
NAND2xp33_ASAP7_75t_SL g497 ( .A(n_465), .B(n_295), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_461), .Y(n_498) );
BUFx12f_ASAP7_75t_SL g499 ( .A(n_474), .Y(n_499) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_483), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_467), .B(n_440), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_473), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_477), .B(n_445), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_486), .B(n_427), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_462), .B(n_446), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_464), .B(n_438), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_464), .B(n_439), .Y(n_507) );
INVx5_ASAP7_75t_L g508 ( .A(n_478), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_468), .A2(n_439), .B1(n_298), .B2(n_338), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_473), .Y(n_510) );
OR2x6_ASAP7_75t_L g511 ( .A(n_484), .B(n_288), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_464), .B(n_439), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_462), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_478), .B(n_453), .Y(n_514) );
INVx4_ASAP7_75t_L g515 ( .A(n_483), .Y(n_515) );
INVx2_ASAP7_75t_SL g516 ( .A(n_478), .Y(n_516) );
NAND3xp33_ASAP7_75t_SL g517 ( .A(n_479), .B(n_312), .C(n_277), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_481), .B(n_425), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_466), .B(n_444), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_466), .B(n_423), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_466), .B(n_444), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_483), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_481), .B(n_423), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_481), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_483), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_472), .A2(n_324), .B1(n_338), .B2(n_298), .Y(n_526) );
BUFx3_ASAP7_75t_L g527 ( .A(n_469), .Y(n_527) );
NOR2xp33_ASAP7_75t_R g528 ( .A(n_480), .B(n_324), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_469), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_481), .Y(n_530) );
NAND3xp33_ASAP7_75t_SL g531 ( .A(n_457), .B(n_340), .C(n_337), .Y(n_531) );
NOR2x1p5_ASAP7_75t_L g532 ( .A(n_469), .B(n_346), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_471), .B(n_289), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_471), .B(n_313), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_471), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_481), .B(n_368), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_457), .Y(n_537) );
NAND2x1p5_ASAP7_75t_L g538 ( .A(n_459), .B(n_279), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_470), .B(n_400), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_508), .Y(n_540) );
INVx4_ASAP7_75t_L g541 ( .A(n_508), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_504), .B(n_290), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_513), .B(n_316), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_508), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_514), .B(n_290), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_506), .A2(n_456), .B(n_430), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_505), .B(n_316), .Y(n_547) );
INVx5_ASAP7_75t_L g548 ( .A(n_523), .Y(n_548) );
AOI21x1_ASAP7_75t_L g549 ( .A1(n_506), .A2(n_456), .B(n_430), .Y(n_549) );
INVx3_ASAP7_75t_L g550 ( .A(n_493), .Y(n_550) );
BUFx2_ASAP7_75t_L g551 ( .A(n_499), .Y(n_551) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_500), .Y(n_552) );
BUFx8_ASAP7_75t_L g553 ( .A(n_487), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_500), .B(n_326), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_SL g555 ( .A1(n_512), .A2(n_364), .B(n_286), .C(n_294), .Y(n_555) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_527), .Y(n_556) );
AND2x2_ASAP7_75t_SL g557 ( .A(n_526), .B(n_365), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_494), .Y(n_558) );
INVx5_ASAP7_75t_L g559 ( .A(n_523), .Y(n_559) );
INVx6_ASAP7_75t_L g560 ( .A(n_488), .Y(n_560) );
INVx3_ASAP7_75t_L g561 ( .A(n_493), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_532), .B(n_351), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_497), .Y(n_563) );
BUFx4f_ASAP7_75t_L g564 ( .A(n_511), .Y(n_564) );
BUFx3_ASAP7_75t_L g565 ( .A(n_489), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_515), .B(n_378), .Y(n_566) );
INVx4_ASAP7_75t_L g567 ( .A(n_518), .Y(n_567) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_528), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_520), .A2(n_456), .B(n_430), .Y(n_569) );
INVxp67_ASAP7_75t_L g570 ( .A(n_492), .Y(n_570) );
CKINVDCx16_ASAP7_75t_R g571 ( .A(n_528), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_492), .B(n_380), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_495), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_496), .A2(n_393), .B1(n_389), .B2(n_370), .Y(n_574) );
BUFx12f_ASAP7_75t_L g575 ( .A(n_518), .Y(n_575) );
BUFx2_ASAP7_75t_L g576 ( .A(n_509), .Y(n_576) );
OAI21x1_ASAP7_75t_L g577 ( .A1(n_538), .A2(n_430), .B(n_470), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_498), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_490), .B(n_393), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_521), .A2(n_430), .B(n_299), .Y(n_580) );
INVx3_ASAP7_75t_L g581 ( .A(n_515), .Y(n_581) );
NOR2x1_ASAP7_75t_L g582 ( .A(n_531), .B(n_374), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_516), .Y(n_583) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_529), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_501), .B(n_433), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_519), .A2(n_301), .B(n_292), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_519), .B(n_309), .Y(n_587) );
BUFx3_ASAP7_75t_L g588 ( .A(n_491), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_531), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_501), .A2(n_379), .B1(n_283), .B2(n_291), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_502), .A2(n_287), .B1(n_305), .B2(n_300), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_510), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_539), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_538), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_536), .Y(n_595) );
A2O1A1Ixp33_ASAP7_75t_L g596 ( .A1(n_503), .A2(n_379), .B(n_333), .C(n_339), .Y(n_596) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_535), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_533), .B(n_311), .Y(n_598) );
OR2x6_ASAP7_75t_L g599 ( .A(n_512), .B(n_395), .Y(n_599) );
NAND3xp33_ASAP7_75t_SL g600 ( .A(n_533), .B(n_329), .C(n_314), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_507), .B(n_331), .Y(n_601) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_522), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_534), .B(n_342), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_537), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_525), .A2(n_358), .B1(n_363), .B2(n_354), .Y(n_605) );
BUFx12f_ASAP7_75t_L g606 ( .A(n_525), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_524), .B(n_367), .Y(n_607) );
INVx5_ASAP7_75t_L g608 ( .A(n_530), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_494), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_506), .A2(n_303), .B(n_302), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_494), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_517), .A2(n_402), .B1(n_412), .B2(n_396), .Y(n_612) );
OAI21x1_ASAP7_75t_L g613 ( .A1(n_577), .A2(n_350), .B(n_307), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_592), .B(n_422), .Y(n_614) );
BUFx3_ASAP7_75t_L g615 ( .A(n_553), .Y(n_615) );
NAND3xp33_ASAP7_75t_SL g616 ( .A(n_589), .B(n_332), .C(n_330), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_SL g617 ( .A1(n_546), .A2(n_304), .B(n_308), .C(n_306), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_558), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_573), .Y(n_619) );
A2O1A1Ixp33_ASAP7_75t_L g620 ( .A1(n_592), .A2(n_448), .B(n_449), .C(n_447), .Y(n_620) );
BUFx12f_ASAP7_75t_L g621 ( .A(n_560), .Y(n_621) );
OAI21x1_ASAP7_75t_L g622 ( .A1(n_549), .A2(n_377), .B(n_350), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_573), .B(n_395), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_548), .B(n_448), .Y(n_624) );
OAI21x1_ASAP7_75t_L g625 ( .A1(n_569), .A2(n_415), .B(n_377), .Y(n_625) );
OAI21x1_ASAP7_75t_L g626 ( .A1(n_580), .A2(n_416), .B(n_415), .Y(n_626) );
BUFx8_ASAP7_75t_L g627 ( .A(n_551), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_570), .A2(n_317), .B(n_310), .Y(n_628) );
NAND2xp33_ASAP7_75t_SL g629 ( .A(n_576), .B(n_386), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_541), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_609), .Y(n_631) );
OA21x2_ASAP7_75t_L g632 ( .A1(n_603), .A2(n_319), .B(n_318), .Y(n_632) );
OR2x6_ASAP7_75t_L g633 ( .A(n_579), .B(n_404), .Y(n_633) );
AO31x2_ASAP7_75t_L g634 ( .A1(n_596), .A2(n_426), .A3(n_431), .B(n_424), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_547), .B(n_386), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_586), .A2(n_476), .B(n_322), .Y(n_636) );
AO21x2_ASAP7_75t_L g637 ( .A1(n_555), .A2(n_409), .B(n_325), .Y(n_637) );
OAI21x1_ASAP7_75t_L g638 ( .A1(n_611), .A2(n_327), .B(n_321), .Y(n_638) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_552), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_550), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_593), .B(n_328), .Y(n_641) );
A2O1A1Ixp33_ASAP7_75t_L g642 ( .A1(n_593), .A2(n_334), .B(n_341), .C(n_335), .Y(n_642) );
OA21x2_ASAP7_75t_L g643 ( .A1(n_610), .A2(n_344), .B(n_343), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_543), .B(n_3), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_557), .B(n_3), .Y(n_645) );
OAI21x1_ASAP7_75t_L g646 ( .A1(n_594), .A2(n_352), .B(n_349), .Y(n_646) );
NAND2x1p5_ASAP7_75t_L g647 ( .A(n_548), .B(n_388), .Y(n_647) );
INVx5_ASAP7_75t_L g648 ( .A(n_552), .Y(n_648) );
NOR2x1_ASAP7_75t_SL g649 ( .A(n_606), .B(n_575), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_SL g650 ( .A1(n_594), .A2(n_356), .B(n_360), .C(n_355), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_548), .B(n_366), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_578), .A2(n_373), .B(n_371), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_542), .B(n_280), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_571), .Y(n_654) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_564), .A2(n_417), .B1(n_388), .B2(n_382), .Y(n_655) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_552), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_572), .A2(n_413), .B1(n_384), .B2(n_387), .Y(n_657) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_582), .B(n_437), .C(n_436), .Y(n_658) );
AO21x2_ASAP7_75t_L g659 ( .A1(n_600), .A2(n_398), .B(n_381), .Y(n_659) );
NAND2x1p5_ASAP7_75t_L g660 ( .A(n_559), .B(n_399), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_612), .A2(n_405), .B(n_401), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_561), .Y(n_662) );
INVx3_ASAP7_75t_L g663 ( .A(n_567), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_604), .Y(n_664) );
INVx4_ASAP7_75t_L g665 ( .A(n_559), .Y(n_665) );
INVxp33_ASAP7_75t_L g666 ( .A(n_566), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_567), .B(n_408), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_585), .B(n_410), .Y(n_668) );
OAI21x1_ASAP7_75t_L g669 ( .A1(n_581), .A2(n_544), .B(n_540), .Y(n_669) );
OAI21x1_ASAP7_75t_SL g670 ( .A1(n_574), .A2(n_419), .B(n_414), .Y(n_670) );
OAI21x1_ASAP7_75t_L g671 ( .A1(n_607), .A2(n_421), .B(n_476), .Y(n_671) );
INVx2_ASAP7_75t_SL g672 ( .A(n_584), .Y(n_672) );
AND2x4_ASAP7_75t_L g673 ( .A(n_595), .B(n_4), .Y(n_673) );
OAI21x1_ASAP7_75t_L g674 ( .A1(n_583), .A2(n_476), .B(n_426), .Y(n_674) );
BUFx8_ASAP7_75t_L g675 ( .A(n_584), .Y(n_675) );
INVx5_ASAP7_75t_L g676 ( .A(n_602), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_565), .B(n_5), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_601), .A2(n_443), .B(n_437), .Y(n_678) );
INVx3_ASAP7_75t_L g679 ( .A(n_556), .Y(n_679) );
AOI21xp33_ASAP7_75t_L g680 ( .A1(n_599), .A2(n_443), .B(n_437), .Y(n_680) );
OAI21x1_ASAP7_75t_L g681 ( .A1(n_598), .A2(n_426), .B(n_424), .Y(n_681) );
BUFx3_ASAP7_75t_L g682 ( .A(n_556), .Y(n_682) );
INVx3_ASAP7_75t_L g683 ( .A(n_602), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_545), .A2(n_454), .B(n_345), .Y(n_684) );
OAI21x1_ASAP7_75t_L g685 ( .A1(n_554), .A2(n_454), .B(n_100), .Y(n_685) );
OA21x2_ASAP7_75t_L g686 ( .A1(n_590), .A2(n_347), .B(n_336), .Y(n_686) );
AO21x2_ASAP7_75t_L g687 ( .A1(n_605), .A2(n_463), .B(n_459), .Y(n_687) );
OA21x2_ASAP7_75t_L g688 ( .A1(n_591), .A2(n_587), .B(n_563), .Y(n_688) );
OAI21x1_ASAP7_75t_L g689 ( .A1(n_608), .A2(n_104), .B(n_102), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_562), .A2(n_357), .B1(n_375), .B2(n_348), .Y(n_690) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_602), .Y(n_691) );
BUFx2_ASAP7_75t_L g692 ( .A(n_568), .Y(n_692) );
AND2x4_ASAP7_75t_L g693 ( .A(n_588), .B(n_8), .Y(n_693) );
NOR2x1_ASAP7_75t_SL g694 ( .A(n_597), .B(n_8), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_673), .Y(n_695) );
INVx3_ASAP7_75t_L g696 ( .A(n_624), .Y(n_696) );
OR2x2_ASAP7_75t_L g697 ( .A(n_633), .B(n_597), .Y(n_697) );
OA21x2_ASAP7_75t_L g698 ( .A1(n_625), .A2(n_403), .B(n_390), .Y(n_698) );
OR2x6_ASAP7_75t_L g699 ( .A(n_615), .B(n_9), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_633), .A2(n_420), .B1(n_406), .B2(n_12), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_645), .A2(n_463), .B1(n_475), .B2(n_459), .Y(n_701) );
BUFx12f_ASAP7_75t_L g702 ( .A(n_621), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_673), .A2(n_463), .B1(n_475), .B2(n_459), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_666), .A2(n_475), .B1(n_463), .B2(n_12), .Y(n_704) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_639), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_666), .A2(n_475), .B1(n_463), .B2(n_13), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_664), .A2(n_14), .B1(n_10), .B2(n_11), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_629), .A2(n_475), .B1(n_463), .B2(n_15), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_629), .A2(n_475), .B1(n_15), .B2(n_11), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_670), .A2(n_17), .B1(n_14), .B2(n_16), .Y(n_710) );
INVx5_ASAP7_75t_L g711 ( .A(n_648), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_617), .A2(n_106), .B(n_105), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_622), .A2(n_626), .B(n_613), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_668), .A2(n_22), .B1(n_20), .B2(n_21), .Y(n_714) );
OAI211xp5_ASAP7_75t_L g715 ( .A1(n_657), .A2(n_26), .B(n_24), .C(n_25), .Y(n_715) );
BUFx5_ASAP7_75t_L g716 ( .A(n_682), .Y(n_716) );
BUFx3_ASAP7_75t_L g717 ( .A(n_675), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_677), .A2(n_31), .B1(n_29), .B2(n_30), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_693), .A2(n_35), .B1(n_33), .B2(n_34), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_644), .B(n_35), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_653), .A2(n_36), .B1(n_37), .B2(n_39), .C(n_42), .Y(n_721) );
OAI21xp5_ASAP7_75t_L g722 ( .A1(n_628), .A2(n_36), .B(n_37), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_693), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_635), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_660), .A2(n_44), .B1(n_42), .B2(n_43), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_636), .A2(n_115), .B(n_113), .Y(n_726) );
INVx3_ASAP7_75t_L g727 ( .A(n_624), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_618), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_620), .A2(n_46), .B(n_47), .C(n_48), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_628), .A2(n_47), .B(n_49), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_653), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_623), .Y(n_732) );
BUFx2_ASAP7_75t_L g733 ( .A(n_675), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_661), .B(n_50), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_627), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_655), .A2(n_56), .B1(n_57), .B2(n_58), .Y(n_736) );
OR2x6_ASAP7_75t_L g737 ( .A(n_672), .B(n_59), .Y(n_737) );
INVx3_ASAP7_75t_L g738 ( .A(n_676), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_686), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_739) );
OAI222xp33_ASAP7_75t_L g740 ( .A1(n_655), .A2(n_60), .B1(n_62), .B2(n_63), .C1(n_64), .C2(n_65), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_692), .B(n_66), .Y(n_741) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_678), .A2(n_681), .B(n_641), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_619), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_654), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_616), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_745) );
OAI22xp33_ASAP7_75t_L g746 ( .A1(n_616), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_746) );
OAI21x1_ASAP7_75t_L g747 ( .A1(n_669), .A2(n_118), .B(n_117), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_686), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_688), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_749) );
AO31x2_ASAP7_75t_L g750 ( .A1(n_620), .A2(n_76), .A3(n_78), .B(n_79), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_688), .A2(n_79), .B1(n_80), .B2(n_81), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_631), .Y(n_752) );
AO31x2_ASAP7_75t_L g753 ( .A1(n_642), .A2(n_80), .A3(n_81), .B(n_82), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_678), .A2(n_641), .B(n_674), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_614), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_690), .B(n_86), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_614), .Y(n_757) );
INVx5_ASAP7_75t_L g758 ( .A(n_648), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_667), .A2(n_87), .B1(n_88), .B2(n_89), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_634), .Y(n_760) );
BUFx8_ASAP7_75t_L g761 ( .A(n_651), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_687), .A2(n_122), .B(n_121), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_649), .B(n_652), .Y(n_763) );
NAND3xp33_ASAP7_75t_L g764 ( .A(n_658), .B(n_124), .C(n_126), .Y(n_764) );
AO31x2_ASAP7_75t_L g765 ( .A1(n_694), .A2(n_687), .A3(n_634), .B(n_662), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_634), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_652), .B(n_271), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_638), .Y(n_768) );
AOI21xp33_ASAP7_75t_L g769 ( .A1(n_658), .A2(n_270), .B(n_130), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_646), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_632), .B(n_131), .Y(n_771) );
OAI21xp5_ASAP7_75t_SL g772 ( .A1(n_647), .A2(n_134), .B(n_140), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_684), .A2(n_141), .B1(n_143), .B2(n_144), .C(n_147), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_659), .A2(n_684), .B1(n_637), .B2(n_665), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_650), .A2(n_148), .B1(n_149), .B2(n_150), .Y(n_775) );
AO21x2_ASAP7_75t_L g776 ( .A1(n_680), .A2(n_153), .B(n_154), .Y(n_776) );
BUFx3_ASAP7_75t_L g777 ( .A(n_711), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_743), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_728), .B(n_679), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_768), .Y(n_780) );
BUFx5_ASAP7_75t_L g781 ( .A(n_770), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_756), .A2(n_637), .B1(n_630), .B2(n_663), .Y(n_782) );
INVxp67_ASAP7_75t_L g783 ( .A(n_741), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_752), .B(n_734), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_760), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_755), .B(n_630), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_757), .B(n_640), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_766), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_705), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_705), .Y(n_790) );
OA21x2_ASAP7_75t_L g791 ( .A1(n_713), .A2(n_742), .B(n_754), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_732), .B(n_676), .Y(n_792) );
INVxp67_ASAP7_75t_SL g793 ( .A(n_723), .Y(n_793) );
INVx5_ASAP7_75t_SL g794 ( .A(n_699), .Y(n_794) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_737), .Y(n_795) );
BUFx3_ASAP7_75t_L g796 ( .A(n_711), .Y(n_796) );
BUFx6f_ASAP7_75t_L g797 ( .A(n_711), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_763), .B(n_676), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_722), .B(n_676), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_747), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_730), .B(n_691), .Y(n_801) );
OR2x2_ASAP7_75t_L g802 ( .A(n_697), .B(n_683), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_753), .B(n_691), .Y(n_803) );
INVx2_ASAP7_75t_SL g804 ( .A(n_758), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_753), .B(n_683), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_753), .B(n_643), .Y(n_806) );
INVx3_ASAP7_75t_L g807 ( .A(n_758), .Y(n_807) );
INVx1_ASAP7_75t_SL g808 ( .A(n_733), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_695), .B(n_648), .Y(n_809) );
INVxp67_ASAP7_75t_SL g810 ( .A(n_696), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_727), .B(n_656), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_750), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_750), .Y(n_813) );
INVxp67_ASAP7_75t_L g814 ( .A(n_699), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_738), .B(n_671), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_720), .B(n_685), .Y(n_816) );
AND2x4_ASAP7_75t_SL g817 ( .A(n_735), .B(n_689), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_765), .Y(n_818) );
INVx2_ASAP7_75t_SL g819 ( .A(n_717), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_765), .Y(n_820) );
BUFx3_ASAP7_75t_L g821 ( .A(n_761), .Y(n_821) );
INVx2_ASAP7_75t_SL g822 ( .A(n_716), .Y(n_822) );
INVx5_ASAP7_75t_L g823 ( .A(n_702), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_714), .Y(n_824) );
OA21x2_ASAP7_75t_L g825 ( .A1(n_762), .A2(n_712), .B(n_774), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_724), .B(n_164), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_765), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_771), .B(n_169), .Y(n_828) );
OR2x2_ASAP7_75t_L g829 ( .A(n_700), .B(n_170), .Y(n_829) );
AND2x4_ASAP7_75t_L g830 ( .A(n_701), .B(n_171), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_731), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_776), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_736), .B(n_172), .Y(n_833) );
INVx3_ASAP7_75t_L g834 ( .A(n_716), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_739), .B(n_174), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_698), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_698), .Y(n_837) );
AND2x2_ASAP7_75t_L g838 ( .A(n_748), .B(n_176), .Y(n_838) );
INVx1_ASAP7_75t_SL g839 ( .A(n_744), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_721), .B(n_269), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_718), .B(n_719), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_725), .Y(n_842) );
INVx3_ASAP7_75t_L g843 ( .A(n_716), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_729), .B(n_177), .Y(n_844) );
INVxp67_ASAP7_75t_SL g845 ( .A(n_709), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_716), .Y(n_846) );
AO21x2_ASAP7_75t_L g847 ( .A1(n_769), .A2(n_179), .B(n_181), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_749), .B(n_182), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_707), .Y(n_849) );
INVxp67_ASAP7_75t_L g850 ( .A(n_745), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_751), .B(n_183), .Y(n_851) );
OR2x2_ASAP7_75t_L g852 ( .A(n_767), .B(n_184), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_715), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_759), .B(n_185), .Y(n_854) );
INVxp67_ASAP7_75t_SL g855 ( .A(n_708), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_764), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_784), .B(n_710), .Y(n_857) );
NAND3xp33_ASAP7_75t_L g858 ( .A(n_782), .B(n_704), .C(n_706), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_805), .B(n_775), .Y(n_859) );
AND2x2_ASAP7_75t_L g860 ( .A(n_805), .B(n_703), .Y(n_860) );
AOI221xp5_ASAP7_75t_L g861 ( .A1(n_831), .A2(n_740), .B1(n_746), .B2(n_773), .C(n_772), .Y(n_861) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_795), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_850), .A2(n_841), .B1(n_783), .B2(n_842), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_780), .Y(n_864) );
AOI211xp5_ASAP7_75t_L g865 ( .A1(n_814), .A2(n_726), .B(n_186), .C(n_187), .Y(n_865) );
INVx3_ASAP7_75t_L g866 ( .A(n_834), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_778), .Y(n_867) );
OAI221xp5_ASAP7_75t_L g868 ( .A1(n_853), .A2(n_192), .B1(n_194), .B2(n_195), .C(n_199), .Y(n_868) );
INVx2_ASAP7_75t_L g869 ( .A(n_780), .Y(n_869) );
OAI211xp5_ASAP7_75t_SL g870 ( .A1(n_808), .A2(n_208), .B(n_209), .C(n_213), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_785), .B(n_214), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_829), .A2(n_217), .B1(n_218), .B2(n_221), .Y(n_872) );
NAND3xp33_ASAP7_75t_SL g873 ( .A(n_839), .B(n_222), .C(n_223), .Y(n_873) );
BUFx2_ASAP7_75t_L g874 ( .A(n_797), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_785), .B(n_229), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_788), .B(n_230), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_788), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_806), .B(n_239), .Y(n_878) );
AND2x2_ASAP7_75t_L g879 ( .A(n_806), .B(n_240), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_803), .B(n_241), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_787), .Y(n_881) );
OR2x2_ASAP7_75t_L g882 ( .A(n_793), .B(n_262), .Y(n_882) );
INVx2_ASAP7_75t_L g883 ( .A(n_818), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_803), .B(n_249), .Y(n_884) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_786), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_818), .Y(n_886) );
BUFx3_ASAP7_75t_L g887 ( .A(n_797), .Y(n_887) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_792), .Y(n_888) );
OR2x2_ASAP7_75t_L g889 ( .A(n_798), .B(n_251), .Y(n_889) );
INVxp67_ASAP7_75t_SL g890 ( .A(n_830), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_820), .Y(n_891) );
BUFx3_ASAP7_75t_L g892 ( .A(n_777), .Y(n_892) );
INVx2_ASAP7_75t_L g893 ( .A(n_827), .Y(n_893) );
A2O1A1Ixp33_ASAP7_75t_SL g894 ( .A1(n_836), .A2(n_252), .B(n_253), .C(n_256), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_781), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_812), .B(n_258), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_781), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_779), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_807), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_813), .B(n_261), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_807), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_807), .Y(n_902) );
INVx2_ASAP7_75t_L g903 ( .A(n_781), .Y(n_903) );
INVx5_ASAP7_75t_L g904 ( .A(n_794), .Y(n_904) );
BUFx6f_ASAP7_75t_L g905 ( .A(n_777), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_802), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_816), .B(n_815), .Y(n_907) );
INVx1_ASAP7_75t_SL g908 ( .A(n_821), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_815), .B(n_846), .Y(n_909) );
OR2x2_ASAP7_75t_L g910 ( .A(n_794), .B(n_819), .Y(n_910) );
BUFx2_ASAP7_75t_L g911 ( .A(n_796), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_781), .Y(n_912) );
OR2x2_ASAP7_75t_L g913 ( .A(n_819), .B(n_810), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g914 ( .A(n_824), .B(n_845), .Y(n_914) );
OAI21xp5_ASAP7_75t_L g915 ( .A1(n_855), .A2(n_849), .B(n_840), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_801), .B(n_837), .Y(n_916) );
INVx2_ASAP7_75t_L g917 ( .A(n_781), .Y(n_917) );
AND2x4_ASAP7_75t_L g918 ( .A(n_834), .B(n_843), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_801), .B(n_836), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_837), .B(n_789), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_804), .Y(n_921) );
INVx2_ASAP7_75t_L g922 ( .A(n_791), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_867), .Y(n_923) );
NOR2xp33_ASAP7_75t_SL g924 ( .A(n_890), .B(n_830), .Y(n_924) );
INVx2_ASAP7_75t_L g925 ( .A(n_877), .Y(n_925) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_863), .B(n_809), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_877), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_862), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_888), .B(n_811), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_907), .B(n_811), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_914), .B(n_799), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_914), .B(n_799), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_861), .A2(n_830), .B1(n_833), .B2(n_844), .Y(n_933) );
BUFx2_ASAP7_75t_L g934 ( .A(n_892), .Y(n_934) );
INVx2_ASAP7_75t_L g935 ( .A(n_864), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_885), .Y(n_936) );
INVx5_ASAP7_75t_SL g937 ( .A(n_905), .Y(n_937) );
HB1xp67_ASAP7_75t_L g938 ( .A(n_869), .Y(n_938) );
INVx1_ASAP7_75t_SL g939 ( .A(n_911), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_881), .Y(n_940) );
AND2x4_ASAP7_75t_L g941 ( .A(n_918), .B(n_822), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_898), .B(n_789), .Y(n_942) );
AOI31xp33_ASAP7_75t_L g943 ( .A1(n_908), .A2(n_828), .A3(n_854), .B(n_823), .Y(n_943) );
AND2x2_ASAP7_75t_L g944 ( .A(n_906), .B(n_790), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_921), .Y(n_945) );
OR2x6_ASAP7_75t_L g946 ( .A(n_895), .B(n_843), .Y(n_946) );
NOR3xp33_ASAP7_75t_SL g947 ( .A(n_873), .B(n_823), .C(n_817), .Y(n_947) );
INVx1_ASAP7_75t_SL g948 ( .A(n_892), .Y(n_948) );
XOR2xp5_ASAP7_75t_L g949 ( .A(n_910), .B(n_823), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_913), .Y(n_950) );
AND2x4_ASAP7_75t_L g951 ( .A(n_918), .B(n_834), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_909), .B(n_826), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_857), .B(n_916), .Y(n_953) );
NOR2x1_ASAP7_75t_L g954 ( .A(n_887), .B(n_826), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_899), .Y(n_955) );
OR2x2_ASAP7_75t_L g956 ( .A(n_916), .B(n_791), .Y(n_956) );
OR2x2_ASAP7_75t_L g957 ( .A(n_919), .B(n_823), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_874), .B(n_848), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_901), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_878), .B(n_851), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_878), .B(n_851), .Y(n_961) );
NOR2xp33_ASAP7_75t_L g962 ( .A(n_904), .B(n_852), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_879), .B(n_838), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_902), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_879), .B(n_838), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_860), .B(n_835), .Y(n_966) );
INVx1_ASAP7_75t_SL g967 ( .A(n_905), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_860), .B(n_835), .Y(n_968) );
OR2x2_ASAP7_75t_L g969 ( .A(n_880), .B(n_825), .Y(n_969) );
HB1xp67_ASAP7_75t_L g970 ( .A(n_883), .Y(n_970) );
INVx2_ASAP7_75t_L g971 ( .A(n_883), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_880), .B(n_817), .Y(n_972) );
NAND2x1p5_ASAP7_75t_L g973 ( .A(n_904), .B(n_800), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_884), .B(n_825), .Y(n_974) );
AND2x4_ASAP7_75t_L g975 ( .A(n_866), .B(n_832), .Y(n_975) );
OR2x2_ASAP7_75t_L g976 ( .A(n_884), .B(n_825), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_905), .B(n_856), .Y(n_977) );
HB1xp67_ASAP7_75t_L g978 ( .A(n_886), .Y(n_978) );
NAND2xp33_ASAP7_75t_SL g979 ( .A(n_905), .B(n_889), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_871), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_953), .B(n_920), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_923), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_925), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_930), .B(n_859), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_936), .B(n_915), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_940), .Y(n_986) );
NAND2x1_ASAP7_75t_L g987 ( .A(n_943), .B(n_897), .Y(n_987) );
INVx1_ASAP7_75t_SL g988 ( .A(n_948), .Y(n_988) );
OR2x2_ASAP7_75t_L g989 ( .A(n_950), .B(n_893), .Y(n_989) );
OR2x2_ASAP7_75t_L g990 ( .A(n_939), .B(n_891), .Y(n_990) );
INVx2_ASAP7_75t_L g991 ( .A(n_925), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_928), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_935), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_929), .B(n_897), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_956), .B(n_903), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_945), .Y(n_996) );
NAND2xp5_ASAP7_75t_SL g997 ( .A(n_924), .B(n_947), .Y(n_997) );
NOR2xp33_ASAP7_75t_L g998 ( .A(n_926), .B(n_904), .Y(n_998) );
INVx2_ASAP7_75t_SL g999 ( .A(n_934), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_955), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_959), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_931), .B(n_896), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_974), .B(n_895), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_952), .B(n_912), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_964), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_938), .B(n_970), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_932), .B(n_896), .Y(n_1007) );
INVx3_ASAP7_75t_L g1008 ( .A(n_946), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_944), .Y(n_1009) );
NOR2x1_ASAP7_75t_L g1010 ( .A(n_949), .B(n_882), .Y(n_1010) );
OAI21xp33_ASAP7_75t_L g1011 ( .A1(n_997), .A2(n_924), .B(n_933), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_984), .B(n_966), .Y(n_1012) );
INVxp67_ASAP7_75t_L g1013 ( .A(n_999), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_982), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_1009), .B(n_968), .Y(n_1015) );
OAI22xp33_ASAP7_75t_L g1016 ( .A1(n_987), .A2(n_957), .B1(n_948), .B2(n_904), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_981), .B(n_970), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_981), .B(n_978), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_1010), .A2(n_954), .B1(n_972), .B2(n_962), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_1003), .B(n_969), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_1004), .B(n_976), .Y(n_1021) );
NAND2xp5_ASAP7_75t_SL g1022 ( .A(n_997), .B(n_979), .Y(n_1022) );
BUFx2_ASAP7_75t_SL g1023 ( .A(n_999), .Y(n_1023) );
OAI31xp33_ASAP7_75t_SL g1024 ( .A1(n_998), .A2(n_960), .A3(n_965), .B(n_963), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_986), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_983), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_983), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_996), .Y(n_1028) );
AOI22xp5_ASAP7_75t_L g1029 ( .A1(n_998), .A2(n_979), .B1(n_961), .B2(n_958), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1000), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1001), .Y(n_1031) );
INVxp67_ASAP7_75t_L g1032 ( .A(n_988), .Y(n_1032) );
INVx2_ASAP7_75t_L g1033 ( .A(n_991), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_995), .B(n_971), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_985), .B(n_942), .Y(n_1035) );
NAND3xp33_ASAP7_75t_L g1036 ( .A(n_992), .B(n_977), .C(n_865), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_1017), .B(n_1006), .Y(n_1037) );
NOR3xp33_ASAP7_75t_SL g1038 ( .A(n_1011), .B(n_870), .C(n_858), .Y(n_1038) );
OAI22xp33_ASAP7_75t_L g1039 ( .A1(n_1019), .A2(n_1008), .B1(n_1007), .B2(n_1002), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1014), .Y(n_1040) );
INVx2_ASAP7_75t_L g1041 ( .A(n_1017), .Y(n_1041) );
INVx1_ASAP7_75t_SL g1042 ( .A(n_1023), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1025), .Y(n_1043) );
NOR3xp33_ASAP7_75t_SL g1044 ( .A(n_1022), .B(n_872), .C(n_868), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1018), .B(n_1006), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1028), .Y(n_1046) );
INVxp67_ASAP7_75t_L g1047 ( .A(n_1036), .Y(n_1047) );
NOR2xp33_ASAP7_75t_L g1048 ( .A(n_1032), .B(n_1005), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1030), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1031), .Y(n_1050) );
AOI21xp33_ASAP7_75t_L g1051 ( .A1(n_1016), .A2(n_990), .B(n_967), .Y(n_1051) );
O2A1O1Ixp33_ASAP7_75t_SL g1052 ( .A1(n_1042), .A2(n_1013), .B(n_1029), .C(n_1024), .Y(n_1052) );
AOI221x1_ASAP7_75t_SL g1053 ( .A1(n_1039), .A2(n_1012), .B1(n_1015), .B2(n_1035), .C(n_1027), .Y(n_1053) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1041), .Y(n_1054) );
NAND3xp33_ASAP7_75t_L g1055 ( .A(n_1038), .B(n_1027), .C(n_1033), .Y(n_1055) );
OAI21xp33_ASAP7_75t_L g1056 ( .A1(n_1047), .A2(n_1020), .B(n_1021), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1037), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1045), .Y(n_1058) );
BUFx2_ASAP7_75t_L g1059 ( .A(n_1040), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1043), .Y(n_1060) );
AOI221xp5_ASAP7_75t_L g1061 ( .A1(n_1052), .A2(n_1048), .B1(n_1050), .B2(n_1049), .C(n_1046), .Y(n_1061) );
AOI21xp5_ASAP7_75t_L g1062 ( .A1(n_1052), .A2(n_1051), .B(n_941), .Y(n_1062) );
A2O1A1Ixp33_ASAP7_75t_L g1063 ( .A1(n_1053), .A2(n_1044), .B(n_1034), .C(n_994), .Y(n_1063) );
NAND2x1_ASAP7_75t_L g1064 ( .A(n_1059), .B(n_1026), .Y(n_1064) );
OA211x2_ASAP7_75t_L g1065 ( .A1(n_1056), .A2(n_937), .B(n_973), .C(n_951), .Y(n_1065) );
NAND4xp25_ASAP7_75t_SL g1066 ( .A(n_1061), .B(n_1055), .C(n_1058), .D(n_1057), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1064), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1065), .Y(n_1068) );
OR2x2_ASAP7_75t_L g1069 ( .A(n_1063), .B(n_1060), .Y(n_1069) );
OAI21xp5_ASAP7_75t_L g1070 ( .A1(n_1062), .A2(n_1054), .B(n_973), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_1066), .A2(n_980), .B1(n_989), .B2(n_946), .Y(n_1071) );
NOR2xp33_ASAP7_75t_L g1072 ( .A(n_1068), .B(n_993), .Y(n_1072) );
INVx5_ASAP7_75t_L g1073 ( .A(n_1072), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_1071), .A2(n_1069), .B1(n_1070), .B2(n_1067), .Y(n_1074) );
BUFx6f_ASAP7_75t_L g1075 ( .A(n_1073), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1073), .Y(n_1076) );
XNOR2x1_ASAP7_75t_L g1077 ( .A(n_1076), .B(n_1074), .Y(n_1077) );
CKINVDCx20_ASAP7_75t_R g1078 ( .A(n_1075), .Y(n_1078) );
AOI22xp5_ASAP7_75t_L g1079 ( .A1(n_1078), .A2(n_975), .B1(n_876), .B2(n_875), .Y(n_1079) );
AOI21xp5_ASAP7_75t_L g1080 ( .A1(n_1077), .A2(n_894), .B(n_847), .Y(n_1080) );
UNKNOWN g1081 ( );
AOI222xp33_ASAP7_75t_L g1082 ( .A1(n_1081), .A2(n_1080), .B1(n_922), .B2(n_900), .C1(n_917), .C2(n_927), .Y(n_1082) );
endmodule