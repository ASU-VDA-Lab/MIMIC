module fake_jpeg_15054_n_110 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_31),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_17),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_11),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_48),
.B(n_30),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_33),
.B(n_35),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_58),
.B(n_62),
.Y(n_69)
);

BUFx24_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_61),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_2),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_33),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_17),
.B(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_23),
.B1(n_28),
.B2(n_14),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_46),
.B1(n_45),
.B2(n_39),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_14),
.B(n_25),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_19),
.B(n_24),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_24),
.B(n_15),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_46),
.B1(n_45),
.B2(n_42),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_72),
.B1(n_71),
.B2(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_67),
.B(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_64),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_75),
.C(n_19),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_41),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_58),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_60),
.B(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_82),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_56),
.C(n_53),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_80),
.C(n_85),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_84),
.Y(n_90)
);

XNOR2x1_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_63),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_62),
.B(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_72),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_19),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_7),
.Y(n_92)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_83),
.B(n_78),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_81),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_96),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_93),
.C(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_88),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_65),
.B(n_75),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_98),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_11),
.B(n_9),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_87),
.C(n_16),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_98),
.Y(n_103)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

AOI31xp67_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_9),
.A3(n_10),
.B(n_99),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_106),
.C(n_105),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_107),
.Y(n_110)
);


endmodule