module fake_jpeg_30141_n_440 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_440);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_440;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx8_ASAP7_75t_SL g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_48),
.Y(n_101)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_57),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_30),
.B(n_9),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_66),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx6f_ASAP7_75t_SL g69 ( 
.A(n_43),
.Y(n_69)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_76),
.Y(n_111)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_74),
.Y(n_107)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_35),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_41),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_83),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_30),
.B(n_9),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_88),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_24),
.B(n_8),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_25),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_36),
.B(n_10),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_90),
.B(n_31),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_120),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_49),
.A2(n_38),
.B1(n_36),
.B2(n_40),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_94),
.A2(n_122),
.B1(n_27),
.B2(n_25),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_38),
.B1(n_37),
.B2(n_20),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_98),
.A2(n_102),
.B1(n_58),
.B2(n_55),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_84),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g173 ( 
.A(n_100),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_48),
.A2(n_22),
.B1(n_20),
.B2(n_37),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_89),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_51),
.A2(n_38),
.B1(n_40),
.B2(n_39),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_67),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_125),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_134),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_72),
.B(n_39),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_135),
.B(n_138),
.Y(n_148)
);

AO22x1_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_62),
.B1(n_81),
.B2(n_79),
.Y(n_140)
);

AO22x1_ASAP7_75t_SL g202 ( 
.A1(n_140),
.A2(n_114),
.B1(n_63),
.B2(n_74),
.Y(n_202)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_143),
.A2(n_170),
.B1(n_175),
.B2(n_101),
.Y(n_176)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_145),
.Y(n_179)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_166),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_111),
.Y(n_151)
);

CKINVDCx9p33_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_152),
.Y(n_183)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_31),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_156),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_20),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_46),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_46),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_108),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_160),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_20),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_37),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_169),
.Y(n_198)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_163),
.Y(n_177)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_71),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_119),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_98),
.A2(n_102),
.B1(n_56),
.B2(n_47),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_107),
.B1(n_68),
.B2(n_101),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_97),
.A2(n_77),
.B1(n_53),
.B2(n_50),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_172),
.A2(n_92),
.B1(n_107),
.B2(n_97),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_37),
.Y(n_174)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_176),
.A2(n_184),
.B1(n_203),
.B2(n_183),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_148),
.B(n_149),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_199),
.B(n_147),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_44),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_116),
.C(n_127),
.Y(n_194)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_166),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_143),
.A2(n_100),
.B(n_125),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_202),
.B1(n_99),
.B2(n_114),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_171),
.A2(n_99),
.B1(n_88),
.B2(n_60),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_144),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_206),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_222),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_159),
.Y(n_206)
);

HAxp5_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_152),
.CON(n_207),
.SN(n_207)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_207),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_208),
.A2(n_92),
.B1(n_173),
.B2(n_96),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_209),
.A2(n_215),
.B(n_227),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_158),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_211),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_190),
.B(n_146),
.Y(n_211)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_212),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_173),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_225),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_215),
.B1(n_211),
.B2(n_225),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_140),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_219),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_218),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_177),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_223),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_226),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_170),
.C(n_169),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_203),
.B1(n_176),
.B2(n_190),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_228),
.A2(n_248),
.B1(n_251),
.B2(n_182),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_184),
.B(n_191),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_230),
.A2(n_223),
.B(n_219),
.Y(n_265)
);

OAI32xp33_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_202),
.A3(n_140),
.B1(n_193),
.B2(n_194),
.Y(n_233)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_202),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_240),
.C(n_243),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_200),
.B1(n_154),
.B2(n_165),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_216),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g268 ( 
.A1(n_238),
.A2(n_252),
.B1(n_226),
.B2(n_224),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_188),
.C(n_178),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_178),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_181),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_141),
.C(n_187),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_182),
.B1(n_154),
.B2(n_165),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_211),
.A2(n_130),
.B1(n_104),
.B2(n_132),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_253),
.A2(n_267),
.B1(n_186),
.B2(n_196),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_239),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_268),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_235),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_259),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_204),
.Y(n_257)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_235),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_227),
.Y(n_260)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_250),
.Y(n_261)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_261),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_206),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_271),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_236),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_263),
.Y(n_291)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_264),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_265),
.A2(n_269),
.B(n_232),
.Y(n_300)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_218),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_247),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_279),
.Y(n_306)
);

XOR2x2_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_221),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_220),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_273),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_239),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_229),
.B(n_195),
.Y(n_275)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_232),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_217),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_181),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_240),
.C(n_244),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_195),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_272),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_258),
.A2(n_238),
.B1(n_242),
.B2(n_244),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_281),
.A2(n_305),
.B1(n_307),
.B2(n_179),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_263),
.B(n_243),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_304),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_294),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_299),
.C(n_301),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_256),
.B(n_242),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_228),
.Y(n_296)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_233),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_260),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_251),
.C(n_252),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_300),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_192),
.C(n_164),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_261),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_258),
.A2(n_248),
.B1(n_231),
.B2(n_217),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_277),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_308),
.B(n_273),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_262),
.B(n_192),
.C(n_161),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_280),
.C(n_268),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_330),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_283),
.B1(n_296),
.B2(n_295),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_313),
.A2(n_317),
.B1(n_322),
.B2(n_327),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_265),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_315),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_329),
.C(n_333),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_287),
.A2(n_267),
.B1(n_291),
.B2(n_284),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_293),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_323),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_268),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_321),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_268),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_284),
.A2(n_273),
.B1(n_254),
.B2(n_269),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_290),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_326),
.Y(n_346)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_306),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_297),
.A2(n_254),
.B1(n_276),
.B2(n_264),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_269),
.C(n_179),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_269),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_331),
.A2(n_299),
.B1(n_285),
.B2(n_302),
.Y(n_341)
);

AOI21xp33_ASAP7_75t_L g332 ( 
.A1(n_297),
.A2(n_223),
.B(n_218),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_332),
.A2(n_300),
.B(n_303),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_168),
.C(n_167),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_336),
.A2(n_10),
.B(n_15),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_328),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_340),
.B(n_343),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_341),
.A2(n_324),
.B1(n_331),
.B2(n_175),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_333),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_310),
.B(n_289),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_348),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_315),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_347),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_288),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_281),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_311),
.B(n_285),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_223),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_303),
.Y(n_351)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_351),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_311),
.B(n_316),
.C(n_329),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_353),
.C(n_356),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_301),
.C(n_305),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_322),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_355),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_319),
.A2(n_175),
.B1(n_130),
.B2(n_104),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_223),
.C(n_145),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_359),
.B(n_360),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_337),
.B(n_12),
.Y(n_361)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_339),
.A2(n_132),
.B1(n_153),
.B2(n_126),
.Y(n_363)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_363),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_346),
.B(n_27),
.Y(n_364)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_338),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_371),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_339),
.A2(n_126),
.B1(n_136),
.B2(n_86),
.Y(n_366)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_366),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_124),
.C(n_163),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_349),
.C(n_344),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_356),
.A2(n_139),
.B(n_212),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_370),
.A2(n_373),
.B(n_14),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_334),
.B(n_212),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_350),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_372),
.B(n_376),
.Y(n_379)
);

OAI321xp33_ASAP7_75t_L g375 ( 
.A1(n_353),
.A2(n_335),
.A3(n_348),
.B1(n_342),
.B2(n_349),
.C(n_352),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_375),
.A2(n_128),
.B1(n_106),
.B2(n_11),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_335),
.B(n_124),
.Y(n_376)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_377),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_384),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_121),
.C(n_73),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_386),
.B(n_387),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_367),
.B(n_139),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_360),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_389),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_17),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_136),
.C(n_54),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_106),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_379),
.A2(n_359),
.B(n_369),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_396),
.Y(n_409)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_380),
.Y(n_395)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_395),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_378),
.A2(n_373),
.B(n_374),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_385),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_397),
.B(n_399),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_376),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_85),
.C(n_75),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_383),
.A2(n_361),
.B1(n_363),
.B2(n_366),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_390),
.A2(n_362),
.B(n_368),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_402),
.B(n_12),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_403),
.B(n_11),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_392),
.A2(n_386),
.B1(n_381),
.B2(n_382),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_405),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_393),
.A2(n_382),
.B1(n_370),
.B2(n_391),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_408),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_394),
.A2(n_128),
.B1(n_115),
.B2(n_112),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_115),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_411),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_412),
.B(n_414),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_413),
.A2(n_415),
.B(n_12),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_396),
.A2(n_402),
.B1(n_400),
.B2(n_398),
.Y(n_414)
);

BUFx24_ASAP7_75t_SL g415 ( 
.A(n_397),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_416),
.Y(n_426)
);

AOI21x1_ASAP7_75t_SL g417 ( 
.A1(n_409),
.A2(n_7),
.B(n_15),
.Y(n_417)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_417),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_407),
.A2(n_410),
.B1(n_409),
.B2(n_406),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_420),
.B(n_424),
.Y(n_429)
);

AOI322xp5_ASAP7_75t_L g422 ( 
.A1(n_414),
.A2(n_87),
.A3(n_67),
.B1(n_7),
.B2(n_13),
.C1(n_4),
.C2(n_6),
.Y(n_422)
);

AND2x2_ASAP7_75t_SL g425 ( 
.A(n_422),
.B(n_6),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_407),
.A2(n_112),
.B1(n_70),
.B2(n_4),
.Y(n_424)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_425),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_421),
.A2(n_6),
.B(n_13),
.Y(n_427)
);

AOI31xp67_ASAP7_75t_SL g433 ( 
.A1(n_427),
.A2(n_419),
.A3(n_2),
.B(n_3),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_417),
.A2(n_0),
.B(n_1),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_428),
.A2(n_423),
.B1(n_418),
.B2(n_422),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_432),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_430),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_433),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_434),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_435),
.C(n_429),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_438),
.B(n_426),
.Y(n_439)
);

O2A1O1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_439),
.A2(n_3),
.B(n_0),
.C(n_2),
.Y(n_440)
);


endmodule