module real_jpeg_23896_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_4),
.A2(n_7),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_4),
.A2(n_21),
.B1(n_22),
.B2(n_32),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_4),
.A2(n_32),
.B1(n_47),
.B2(n_48),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_4),
.A2(n_32),
.B1(n_66),
.B2(n_67),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_4),
.B(n_20),
.C(n_22),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_4),
.B(n_19),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_4),
.B(n_44),
.C(n_47),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_4),
.B(n_63),
.C(n_66),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_4),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_4),
.B(n_109),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_4),
.B(n_56),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_6),
.A2(n_21),
.B1(n_22),
.B2(n_53),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_6),
.A2(n_53),
.B1(n_66),
.B2(n_67),
.Y(n_184)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_8),
.A2(n_21),
.B1(n_22),
.B2(n_39),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_8),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_8),
.A2(n_39),
.B1(n_66),
.B2(n_67),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_9),
.A2(n_21),
.B1(n_22),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_9),
.A2(n_29),
.B1(n_47),
.B2(n_48),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_9),
.A2(n_29),
.B1(n_66),
.B2(n_67),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_11),
.Y(n_128)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_11),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_85),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_84),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_69),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_16),
.B(n_69),
.Y(n_84)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_16),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_37),
.CI(n_49),
.CON(n_16),
.SN(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_25),
.B(n_30),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_18),
.A2(n_30),
.B(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_19),
.A2(n_31),
.B1(n_35),
.B2(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_19),
.B(n_35),
.Y(n_102)
);

AO22x1_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_19)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_20),
.A2(n_24),
.B1(n_28),
.B2(n_34),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_21),
.A2(n_22),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

INVx5_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_22),
.B(n_214),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_34),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_42),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_46),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_41),
.A2(n_46),
.B(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_42),
.B(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_42),
.A2(n_56),
.B1(n_83),
.B2(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

OA22x2_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_81),
.B(n_82),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_46),
.A2(n_82),
.B(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_47),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_48),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_47),
.B(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.C(n_57),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_SL g124 ( 
.A(n_50),
.B(n_125),
.C(n_132),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_50),
.A2(n_75),
.B1(n_132),
.B2(n_133),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_50),
.A2(n_75),
.B1(n_111),
.B2(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_50),
.B(n_111),
.C(n_177),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_79),
.C(n_80),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_57),
.A2(n_73),
.B1(n_80),
.B2(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_68),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_59),
.B(n_99),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_61),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_61),
.A2(n_99),
.B1(n_109),
.B2(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_65),
.A2(n_98),
.B(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_66),
.B(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.C(n_77),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_70),
.A2(n_76),
.B1(n_79),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_79),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_76),
.B(n_151),
.C(n_159),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_76),
.A2(n_79),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_76),
.A2(n_79),
.B1(n_159),
.B2(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_77),
.A2(n_78),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_79),
.B(n_132),
.C(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_80),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

OAI211xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_134),
.B(n_141),
.C(n_282),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_119),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_87),
.B(n_119),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_104),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_88),
.B(n_106),
.C(n_114),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_95),
.B(n_100),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_100),
.B1(n_101),
.B2(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_89),
.A2(n_96),
.B1(n_122),
.B2(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_91),
.B(n_186),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_94),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_92),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_93),
.A2(n_127),
.B(n_154),
.Y(n_153)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_93),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_96),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_114),
.B2(n_115),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_107),
.B(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_111),
.B(n_198),
.C(n_200),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_111),
.A2(n_188),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_124),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_123),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_126),
.A2(n_129),
.B1(n_130),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_126),
.Y(n_273)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_129),
.A2(n_130),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_129),
.A2(n_130),
.B1(n_211),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_130),
.B(n_205),
.C(n_211),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_130),
.B(n_182),
.C(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_132),
.A2(n_133),
.B1(n_173),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_132),
.A2(n_133),
.B1(n_157),
.B2(n_170),
.Y(n_250)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_133),
.B(n_157),
.C(n_251),
.Y(n_254)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_SL g141 ( 
.A(n_135),
.B(n_142),
.C(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_136),
.B(n_137),
.Y(n_282)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_163),
.B(n_281),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_161),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_145),
.B(n_161),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_150),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_146),
.B(n_148),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_150),
.B(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_151),
.A2(n_152),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_157),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_155),
.A2(n_184),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_157),
.A2(n_170),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_157),
.B(n_228),
.Y(n_240)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_159),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_276),
.B(n_280),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_201),
.B(n_262),
.C(n_275),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_190),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_166),
.B(n_190),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_176),
.B2(n_189),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_168)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_169),
.B(n_175),
.C(n_189),
.Y(n_263)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_187),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_181),
.A2(n_182),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_182),
.B(n_236),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.C(n_197),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_191),
.A2(n_192),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_197),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_200),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_198),
.B(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_200),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_261),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_220),
.B(n_260),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_217),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_204),
.B(n_217),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_205),
.A2(n_206),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_210),
.B(n_225),
.Y(n_238)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_253),
.B(n_259),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_247),
.B(n_252),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_239),
.B(n_246),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_229),
.B(n_238),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_226),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_235),
.B(n_237),
.Y(n_229)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_240),
.B(n_241),
.Y(n_246)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_244),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_254),
.B(n_255),
.Y(n_259)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_256),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_264),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_274),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_271),
.B2(n_272),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_272),
.C(n_274),
.Y(n_277)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_278),
.Y(n_280)
);


endmodule