module real_aes_8742_n_271 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_271);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_271;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_755;
wire n_656;
wire n_284;
wire n_316;
wire n_532;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_753;
wire n_283;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_475;
wire n_554;
wire n_798;
wire n_668;
wire n_797;
AOI22xp33_ASAP7_75t_SL g556 ( .A1(n_0), .A2(n_234), .B1(n_557), .B2(n_558), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_1), .A2(n_259), .B1(n_329), .B2(n_334), .Y(n_328) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_2), .A2(n_106), .B1(n_560), .B2(n_562), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_3), .A2(n_248), .B1(n_600), .B2(n_650), .Y(n_817) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_4), .A2(n_36), .B1(n_461), .B2(n_600), .C(n_602), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_5), .B(n_327), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_6), .B(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_7), .A2(n_95), .B1(n_339), .B2(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_8), .A2(n_21), .B1(n_303), .B2(n_314), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_9), .A2(n_159), .B1(n_383), .B2(n_499), .Y(n_657) );
XOR2x2_ASAP7_75t_L g451 ( .A(n_10), .B(n_452), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_11), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_12), .A2(n_176), .B1(n_339), .B2(n_455), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_13), .Y(n_666) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_14), .A2(n_116), .B1(n_383), .B2(n_384), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_15), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_16), .A2(n_212), .B1(n_347), .B2(n_500), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_17), .A2(n_213), .B1(n_326), .B2(n_518), .C(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_18), .A2(n_136), .B1(n_378), .B2(n_387), .Y(n_682) );
AOI222xp33_ASAP7_75t_L g350 ( .A1(n_19), .A2(n_108), .B1(n_131), .B2(n_351), .C1(n_354), .C2(n_359), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g377 ( .A1(n_20), .A2(n_184), .B1(n_378), .B2(n_379), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_22), .Y(n_777) );
INVx1_ASAP7_75t_L g747 ( .A(n_23), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_24), .A2(n_264), .B1(n_521), .B2(n_549), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_25), .A2(n_32), .B1(n_314), .B2(n_465), .Y(n_678) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_26), .A2(n_81), .B1(n_293), .B2(n_298), .Y(n_302) );
INVx1_ASAP7_75t_L g799 ( .A(n_26), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_27), .A2(n_44), .B1(n_586), .B2(n_587), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_28), .A2(n_34), .B1(n_356), .B2(n_359), .Y(n_368) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_29), .A2(n_46), .B1(n_443), .B2(n_457), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_30), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_31), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_33), .A2(n_152), .B1(n_345), .B2(n_347), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_35), .A2(n_189), .B1(n_437), .B2(n_439), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_37), .A2(n_163), .B1(n_418), .B2(n_574), .Y(n_573) );
AO22x1_ASAP7_75t_L g397 ( .A1(n_38), .A2(n_398), .B1(n_449), .B2(n_450), .Y(n_397) );
INVx1_ASAP7_75t_L g449 ( .A(n_38), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_39), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_40), .A2(n_215), .B1(n_442), .B2(n_443), .Y(n_441) );
AOI222xp33_ASAP7_75t_L g527 ( .A1(n_41), .A2(n_126), .B1(n_192), .B2(n_351), .C1(n_354), .C2(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_42), .A2(n_263), .B1(n_335), .B2(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_43), .A2(n_231), .B1(n_466), .B2(n_513), .Y(n_675) );
AO22x2_ASAP7_75t_L g300 ( .A1(n_45), .A2(n_84), .B1(n_293), .B2(n_294), .Y(n_300) );
INVx1_ASAP7_75t_L g800 ( .A(n_45), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_47), .A2(n_56), .B1(n_354), .B2(n_528), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_48), .A2(n_186), .B1(n_566), .B2(n_656), .Y(n_655) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_49), .A2(n_96), .B1(n_437), .B2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_50), .A2(n_157), .B1(n_309), .B2(n_314), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_51), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_52), .A2(n_270), .B1(n_309), .B2(n_466), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_53), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_54), .Y(n_767) );
XOR2xp5_ASAP7_75t_L g285 ( .A(n_55), .B(n_286), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_57), .A2(n_235), .B1(n_524), .B2(n_525), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_58), .A2(n_251), .B1(n_433), .B2(n_434), .Y(n_432) );
XNOR2x1_ASAP7_75t_L g659 ( .A(n_59), .B(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_60), .A2(n_135), .B1(n_335), .B2(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_61), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_62), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_63), .A2(n_236), .B1(n_461), .B2(n_462), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_64), .A2(n_187), .B1(n_345), .B2(n_379), .Y(n_718) );
AOI222xp33_ASAP7_75t_L g621 ( .A1(n_65), .A2(n_86), .B1(n_146), .B2(n_417), .C1(n_622), .C2(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_66), .B(n_519), .Y(n_713) );
INVx1_ASAP7_75t_L g473 ( .A(n_67), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_68), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_69), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_70), .A2(n_122), .B1(n_466), .B2(n_502), .C(n_610), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_71), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_72), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_73), .A2(n_153), .B1(n_386), .B2(n_387), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_74), .A2(n_252), .B1(n_357), .B2(n_374), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_75), .A2(n_82), .B1(n_321), .B2(n_326), .Y(n_320) );
AOI22xp33_ASAP7_75t_SL g818 ( .A1(n_76), .A2(n_233), .B1(n_819), .B2(n_821), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_77), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_78), .A2(n_203), .B1(n_334), .B2(n_360), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_79), .A2(n_124), .B1(n_465), .B2(n_466), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_80), .A2(n_142), .B1(n_303), .B2(n_524), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_83), .Y(n_697) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_85), .A2(n_175), .B1(n_584), .B2(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g278 ( .A(n_87), .B(n_279), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_88), .A2(n_109), .B1(n_339), .B2(n_341), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_89), .A2(n_193), .B1(n_329), .B2(n_356), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_90), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_91), .A2(n_183), .B1(n_386), .B2(n_387), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_92), .A2(n_111), .B1(n_341), .B2(n_442), .Y(n_511) );
INVx1_ASAP7_75t_L g275 ( .A(n_93), .Y(n_275) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_94), .A2(n_219), .B1(n_374), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_97), .A2(n_226), .B1(n_303), .B2(n_458), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_98), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_99), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_100), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_101), .A2(n_223), .B1(n_339), .B2(n_587), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_102), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_103), .A2(n_206), .B1(n_455), .B2(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_104), .A2(n_121), .B1(n_341), .B2(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_105), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_107), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_110), .A2(n_132), .B1(n_335), .B2(n_374), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_112), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_113), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_114), .A2(n_208), .B1(n_442), .B2(n_586), .Y(n_771) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_115), .A2(n_225), .B1(n_386), .B2(n_461), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_117), .A2(n_158), .B1(n_378), .B2(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_118), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_119), .B(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_120), .A2(n_211), .B1(n_289), .B2(n_438), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_123), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_125), .A2(n_256), .B1(n_357), .B2(n_359), .Y(n_667) );
AOI22xp33_ASAP7_75t_SL g498 ( .A1(n_127), .A2(n_155), .B1(n_499), .B2(n_500), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_128), .A2(n_199), .B1(n_529), .B2(n_548), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_129), .Y(n_619) );
XOR2x2_ASAP7_75t_L g631 ( .A(n_130), .B(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_133), .A2(n_210), .B1(n_446), .B2(n_566), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_134), .Y(n_552) );
INVx2_ASAP7_75t_L g279 ( .A(n_137), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_138), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_139), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_140), .A2(n_145), .B1(n_458), .B2(n_525), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_141), .A2(n_209), .B1(n_465), .B2(n_584), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_143), .A2(n_224), .B1(n_462), .B2(n_558), .Y(n_825) );
INVx1_ASAP7_75t_L g389 ( .A(n_144), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_147), .B(n_327), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_148), .B(n_321), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_149), .A2(n_265), .B1(n_314), .B2(n_437), .Y(n_772) );
AND2x6_ASAP7_75t_L g274 ( .A(n_150), .B(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_150), .Y(n_793) );
AO22x2_ASAP7_75t_L g292 ( .A1(n_151), .A2(n_218), .B1(n_293), .B2(n_294), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_154), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_156), .A2(n_249), .B1(n_521), .B2(n_549), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_160), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_161), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_162), .A2(n_246), .B1(n_744), .B2(n_746), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_164), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_165), .A2(n_207), .B1(n_330), .B2(n_335), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_166), .B(n_740), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_167), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_168), .A2(n_243), .B1(n_315), .B2(n_560), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_169), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_170), .B(n_371), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_171), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_172), .A2(n_269), .B1(n_321), .B2(n_326), .Y(n_468) );
XNOR2x1_ASAP7_75t_L g567 ( .A(n_173), .B(n_568), .Y(n_567) );
AO22x2_ASAP7_75t_L g297 ( .A1(n_174), .A2(n_237), .B1(n_293), .B2(n_298), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_177), .A2(n_267), .B1(n_303), .B2(n_345), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_178), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_179), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_180), .A2(n_216), .B1(n_345), .B2(n_347), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_181), .A2(n_250), .B1(n_457), .B2(n_458), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_182), .Y(n_663) );
AOI22xp5_ASAP7_75t_SL g479 ( .A1(n_185), .A2(n_480), .B1(n_506), .B2(n_507), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g507 ( .A(n_185), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_188), .Y(n_516) );
INVxp67_ASAP7_75t_L g837 ( .A(n_190), .Y(n_837) );
XNOR2x1_ASAP7_75t_L g839 ( .A(n_190), .B(n_803), .Y(n_839) );
AO22x1_ASAP7_75t_L g597 ( .A1(n_191), .A2(n_598), .B1(n_625), .B2(n_626), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_191), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_194), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_195), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_196), .Y(n_646) );
AOI22xp33_ASAP7_75t_SL g736 ( .A1(n_197), .A2(n_201), .B1(n_529), .B2(n_737), .Y(n_736) );
AOI22xp33_ASAP7_75t_SL g694 ( .A1(n_198), .A2(n_266), .B1(n_383), .B2(n_695), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_200), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_202), .B(n_371), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_204), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_205), .B(n_327), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_214), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_217), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_218), .B(n_798), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_220), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_221), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_222), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_227), .Y(n_686) );
AOI22xp33_ASAP7_75t_SL g823 ( .A1(n_228), .A2(n_232), .B1(n_378), .B2(n_824), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_229), .Y(n_419) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_230), .A2(n_268), .B1(n_349), .B2(n_448), .Y(n_717) );
INVx1_ASAP7_75t_L g796 ( .A(n_237), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_238), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_239), .A2(n_803), .B1(n_826), .B2(n_827), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_239), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_240), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_241), .B(n_529), .Y(n_642) );
OA22x2_ASAP7_75t_L g752 ( .A1(n_242), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_752) );
CKINVDCx16_ASAP7_75t_R g753 ( .A(n_242), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_244), .B(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_245), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_247), .Y(n_539) );
INVx1_ASAP7_75t_L g293 ( .A(n_253), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_253), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_254), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_255), .Y(n_550) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_257), .A2(n_272), .B(n_280), .C(n_801), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_258), .A2(n_261), .B1(n_288), .B2(n_303), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_260), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_262), .Y(n_421) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_275), .Y(n_792) );
OAI21xp5_ASAP7_75t_L g835 ( .A1(n_276), .A2(n_791), .B(n_836), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_277), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_595), .B1(n_786), .B2(n_787), .C(n_788), .Y(n_280) );
INVx1_ASAP7_75t_L g786 ( .A(n_281), .Y(n_786) );
XOR2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_477), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_392), .B2(n_476), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AO22x2_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_362), .B1(n_390), .B2(n_391), .Y(n_284) );
INVx1_ASAP7_75t_L g390 ( .A(n_285), .Y(n_390) );
NAND5xp2_ASAP7_75t_SL g286 ( .A(n_287), .B(n_308), .C(n_319), .D(n_337), .E(n_350), .Y(n_286) );
BUFx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx3_ASAP7_75t_L g383 ( .A(n_289), .Y(n_383) );
INVx6_ASAP7_75t_L g444 ( .A(n_289), .Y(n_444) );
BUFx3_ASAP7_75t_L g558 ( .A(n_289), .Y(n_558) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_299), .Y(n_289) );
AND2x2_ASAP7_75t_L g346 ( .A(n_290), .B(n_311), .Y(n_346) );
AND2x6_ASAP7_75t_L g349 ( .A(n_290), .B(n_324), .Y(n_349) );
AND2x6_ASAP7_75t_L g352 ( .A(n_290), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_296), .Y(n_290) );
AND2x2_ASAP7_75t_L g313 ( .A(n_291), .B(n_297), .Y(n_313) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g306 ( .A(n_292), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_292), .B(n_297), .Y(n_318) );
AND2x2_ASAP7_75t_L g333 ( .A(n_292), .B(n_302), .Y(n_333) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g298 ( .A(n_295), .Y(n_298) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g307 ( .A(n_297), .Y(n_307) );
INVx1_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
AND2x2_ASAP7_75t_L g305 ( .A(n_299), .B(n_306), .Y(n_305) );
AND2x6_ASAP7_75t_L g327 ( .A(n_299), .B(n_313), .Y(n_327) );
NAND2x1p5_ASAP7_75t_L g409 ( .A(n_299), .B(n_313), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_299), .B(n_306), .Y(n_613) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g312 ( .A(n_300), .Y(n_312) );
INVx1_ASAP7_75t_L g317 ( .A(n_300), .Y(n_317) );
OR2x2_ASAP7_75t_L g325 ( .A(n_300), .B(n_301), .Y(n_325) );
AND2x2_ASAP7_75t_L g353 ( .A(n_300), .B(n_302), .Y(n_353) );
AND2x2_ASAP7_75t_L g311 ( .A(n_301), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx5_ASAP7_75t_L g384 ( .A(n_304), .Y(n_384) );
INVx4_ASAP7_75t_L g438 ( .A(n_304), .Y(n_438) );
INVx2_ASAP7_75t_L g457 ( .A(n_304), .Y(n_457) );
BUFx3_ASAP7_75t_L g820 ( .A(n_304), .Y(n_820) );
INVx8_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g340 ( .A(n_306), .B(n_311), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_306), .B(n_311), .Y(n_608) );
INVx1_ASAP7_75t_L g361 ( .A(n_307), .Y(n_361) );
BUFx2_ASAP7_75t_L g566 ( .A(n_309), .Y(n_566) );
BUFx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_310), .Y(n_386) );
INVx2_ASAP7_75t_L g435 ( .A(n_310), .Y(n_435) );
BUFx3_ASAP7_75t_L g465 ( .A(n_310), .Y(n_465) );
BUFx3_ASAP7_75t_L g525 ( .A(n_310), .Y(n_525) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
AND2x4_ASAP7_75t_L g342 ( .A(n_311), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g331 ( .A(n_312), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g388 ( .A(n_312), .Y(n_388) );
AND2x4_ASAP7_75t_L g323 ( .A(n_313), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g405 ( .A(n_313), .Y(n_405) );
BUFx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx4f_ASAP7_75t_SL g439 ( .A(n_315), .Y(n_439) );
BUFx2_ASAP7_75t_L g458 ( .A(n_315), .Y(n_458) );
INVx6_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g562 ( .A(n_316), .Y(n_562) );
INVx1_ASAP7_75t_L g653 ( .A(n_316), .Y(n_653) );
INVx1_ASAP7_75t_SL g821 ( .A(n_316), .Y(n_821) );
OR2x6_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g336 ( .A(n_317), .Y(n_336) );
INVx1_ASAP7_75t_L g343 ( .A(n_318), .Y(n_343) );
AND2x2_ASAP7_75t_SL g319 ( .A(n_320), .B(n_328), .Y(n_319) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g371 ( .A(n_322), .Y(n_371) );
INVx5_ASAP7_75t_L g519 ( .A(n_322), .Y(n_519) );
INVx2_ASAP7_75t_L g742 ( .A(n_322), .Y(n_742) );
INVx4_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g404 ( .A(n_325), .B(n_405), .Y(n_404) );
BUFx4f_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g578 ( .A(n_327), .Y(n_578) );
BUFx2_ASAP7_75t_L g740 ( .A(n_327), .Y(n_740) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_330), .Y(n_374) );
BUFx2_ASAP7_75t_L g412 ( .A(n_330), .Y(n_412) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_330), .Y(n_529) );
BUFx4f_ASAP7_75t_SL g692 ( .A(n_330), .Y(n_692) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g358 ( .A(n_332), .Y(n_358) );
AND2x4_ASAP7_75t_L g335 ( .A(n_333), .B(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g357 ( .A(n_333), .B(n_358), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_333), .B(n_388), .Y(n_423) );
BUFx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g580 ( .A(n_335), .Y(n_580) );
INVx1_ASAP7_75t_L g745 ( .A(n_335), .Y(n_745) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_344), .Y(n_337) );
BUFx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx3_ASAP7_75t_L g378 ( .A(n_340), .Y(n_378) );
BUFx3_ASAP7_75t_L g448 ( .A(n_340), .Y(n_448) );
BUFx3_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx3_ASAP7_75t_L g379 ( .A(n_342), .Y(n_379) );
BUFx3_ASAP7_75t_L g466 ( .A(n_342), .Y(n_466) );
BUFx2_ASAP7_75t_SL g500 ( .A(n_342), .Y(n_500) );
BUFx2_ASAP7_75t_SL g584 ( .A(n_342), .Y(n_584) );
INVx1_ASAP7_75t_L g780 ( .A(n_342), .Y(n_780) );
AND2x2_ASAP7_75t_L g387 ( .A(n_343), .B(n_388), .Y(n_387) );
BUFx3_ASAP7_75t_L g433 ( .A(n_345), .Y(n_433) );
BUFx3_ASAP7_75t_L g557 ( .A(n_345), .Y(n_557) );
INVx3_ASAP7_75t_L g651 ( .A(n_345), .Y(n_651) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx2_ASAP7_75t_SL g461 ( .A(n_346), .Y(n_461) );
INVx2_ASAP7_75t_L g514 ( .A(n_346), .Y(n_514) );
INVx5_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g442 ( .A(n_348), .Y(n_442) );
INVx4_ASAP7_75t_L g587 ( .A(n_348), .Y(n_587) );
INVx2_ASAP7_75t_SL g695 ( .A(n_348), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_348), .A2(n_444), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx11_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx11_ASAP7_75t_L g463 ( .A(n_349), .Y(n_463) );
INVx2_ASAP7_75t_SL g414 ( .A(n_351), .Y(n_414) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g367 ( .A(n_352), .Y(n_367) );
BUFx3_ASAP7_75t_L g472 ( .A(n_352), .Y(n_472) );
INVx2_ASAP7_75t_SL g488 ( .A(n_352), .Y(n_488) );
INVx4_ASAP7_75t_L g571 ( .A(n_352), .Y(n_571) );
AND2x4_ASAP7_75t_L g360 ( .A(n_353), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g428 ( .A(n_353), .Y(n_428) );
INVx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx4f_ASAP7_75t_SL g737 ( .A(n_356), .Y(n_737) );
BUFx12f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_357), .Y(n_418) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_357), .Y(n_549) );
BUFx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_360), .Y(n_521) );
BUFx2_ASAP7_75t_SL g574 ( .A(n_360), .Y(n_574) );
BUFx2_ASAP7_75t_SL g746 ( .A(n_360), .Y(n_746) );
INVx1_ASAP7_75t_L g429 ( .A(n_361), .Y(n_429) );
INVx2_ASAP7_75t_L g391 ( .A(n_362), .Y(n_391) );
XOR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_389), .Y(n_362) );
NAND2x1p5_ASAP7_75t_L g363 ( .A(n_364), .B(n_375), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_369), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_367), .B(n_368), .Y(n_365) );
OAI221xp5_ASAP7_75t_L g639 ( .A1(n_367), .A2(n_416), .B1(n_640), .B2(n_641), .C(n_642), .Y(n_639) );
OAI21xp33_ASAP7_75t_SL g809 ( .A1(n_367), .A2(n_810), .B(n_811), .Y(n_809) );
NAND3xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .C(n_373), .Y(n_369) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_374), .Y(n_544) );
NOR2x1_ASAP7_75t_L g375 ( .A(n_376), .B(n_381), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_380), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_385), .Y(n_381) );
INVx4_ASAP7_75t_L g601 ( .A(n_386), .Y(n_601) );
INVx3_ASAP7_75t_L g394 ( .A(n_391), .Y(n_394) );
INVx1_ASAP7_75t_L g476 ( .A(n_392), .Y(n_476) );
XOR2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_451), .B2(n_475), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g450 ( .A(n_398), .Y(n_450) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_430), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_410), .C(n_420), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_406), .B2(n_407), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_402), .A2(n_635), .B1(n_636), .B2(n_637), .Y(n_634) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_404), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_404), .A2(n_407), .B1(n_663), .B2(n_664), .Y(n_662) );
BUFx3_ASAP7_75t_L g807 ( .A(n_404), .Y(n_807) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g486 ( .A(n_408), .Y(n_486) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx3_ASAP7_75t_L g540 ( .A(n_409), .Y(n_540) );
OAI222xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B1(n_414), .B2(n_415), .C1(n_416), .C2(n_419), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_411), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_668) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B1(n_424), .B2(n_425), .Y(n_420) );
OAI22xp5_ASAP7_75t_SL g551 ( .A1(n_422), .A2(n_425), .B1(n_552), .B2(n_553), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_422), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_617) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx4_ASAP7_75t_L g494 ( .A(n_423), .Y(n_494) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_423), .Y(n_645) );
OAI22xp33_ASAP7_75t_SL g766 ( .A1(n_423), .A2(n_425), .B1(n_767), .B2(n_768), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_425), .A2(n_644), .B1(n_645), .B2(n_646), .Y(n_643) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g620 ( .A(n_426), .Y(n_620) );
CKINVDCx16_ASAP7_75t_R g426 ( .A(n_427), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_427), .A2(n_492), .B1(n_493), .B2(n_495), .Y(n_491) );
OR2x6_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_440), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_436), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g561 ( .A(n_438), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g615 ( .A(n_439), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_441), .B(n_445), .Y(n_440) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g455 ( .A(n_444), .Y(n_455) );
INVx3_ASAP7_75t_L g524 ( .A(n_444), .Y(n_524) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx4f_ASAP7_75t_SL g499 ( .A(n_448), .Y(n_499) );
INVx1_ASAP7_75t_SL g475 ( .A(n_451), .Y(n_475) );
NOR4xp75_ASAP7_75t_L g452 ( .A(n_453), .B(n_459), .C(n_467), .D(n_470), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_454), .B(n_456), .Y(n_453) );
INVx2_ASAP7_75t_L g604 ( .A(n_455), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_460), .B(n_464), .Y(n_459) );
INVx4_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g502 ( .A(n_463), .Y(n_502) );
INVx2_ASAP7_75t_SL g656 ( .A(n_463), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_468), .B(n_469), .Y(n_467) );
OAI21xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_473), .B(n_474), .Y(n_470) );
OAI21xp33_ASAP7_75t_L g665 ( .A1(n_471), .A2(n_666), .B(n_667), .Y(n_665) );
OAI21xp33_ASAP7_75t_SL g763 ( .A1(n_471), .A2(n_764), .B(n_765), .Y(n_763) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_533), .B1(n_593), .B2(n_594), .Y(n_477) );
INVx1_ASAP7_75t_L g594 ( .A(n_478), .Y(n_594) );
AO22x1_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_508), .B1(n_531), .B2(n_532), .Y(n_478) );
INVx1_ASAP7_75t_L g531 ( .A(n_479), .Y(n_531) );
INVx2_ASAP7_75t_L g506 ( .A(n_480), .Y(n_506) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_496), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_487), .C(n_491), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_485), .B2(n_486), .Y(n_482) );
OAI22xp5_ASAP7_75t_SL g538 ( .A1(n_484), .A2(n_539), .B1(n_540), .B2(n_541), .Y(n_538) );
INVx1_ASAP7_75t_L g759 ( .A(n_484), .Y(n_759) );
OA211x2_ASAP7_75t_L g515 ( .A1(n_486), .A2(n_516), .B(n_517), .C(n_520), .Y(n_515) );
OAI21xp5_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_489), .B(n_490), .Y(n_487) );
OAI222xp33_ASAP7_75t_L g542 ( .A1(n_488), .A2(n_543), .B1(n_545), .B2(n_546), .C1(n_547), .C2(n_550), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_493), .A2(n_620), .B1(n_813), .B2(n_814), .Y(n_812) );
INVx3_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g671 ( .A(n_494), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_503), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_501), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g532 ( .A(n_508), .Y(n_532) );
XOR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_530), .Y(n_508) );
NAND4xp75_ASAP7_75t_L g509 ( .A(n_510), .B(n_515), .C(n_522), .D(n_527), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g586 ( .A(n_514), .Y(n_586) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_526), .Y(n_522) );
INVx1_ASAP7_75t_L g778 ( .A(n_525), .Y(n_778) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g624 ( .A(n_529), .Y(n_624) );
INVx1_ASAP7_75t_L g593 ( .A(n_533), .Y(n_593) );
OAI22xp5_ASAP7_75t_SL g533 ( .A1(n_534), .A2(n_567), .B1(n_591), .B2(n_592), .Y(n_533) );
INVx2_ASAP7_75t_L g591 ( .A(n_534), .Y(n_591) );
XNOR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_554), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .C(n_551), .Y(n_537) );
INVx2_ASAP7_75t_L g638 ( .A(n_540), .Y(n_638) );
BUFx3_ASAP7_75t_L g761 ( .A(n_540), .Y(n_761) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx4f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_563), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .Y(n_555) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g592 ( .A(n_567), .Y(n_592) );
AND2x4_ASAP7_75t_L g568 ( .A(n_569), .B(n_581), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_575), .Y(n_569) );
OAI21xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_572), .B(n_573), .Y(n_570) );
INVx4_ASAP7_75t_L g622 ( .A(n_571), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_571), .A2(n_686), .B(n_687), .Y(n_685) );
OAI21xp5_ASAP7_75t_L g709 ( .A1(n_571), .A2(n_710), .B(n_711), .Y(n_709) );
OAI21xp5_ASAP7_75t_SL g734 ( .A1(n_571), .A2(n_735), .B(n_736), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .C(n_579), .Y(n_575) );
NOR2x1_ASAP7_75t_L g581 ( .A(n_582), .B(n_588), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g787 ( .A(n_595), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B1(n_627), .B2(n_785), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g626 ( .A(n_598), .Y(n_626) );
AND4x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_609), .C(n_616), .D(n_621), .Y(n_598) );
INVx4_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B1(n_605), .B2(n_606), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_604), .A2(n_732), .B1(n_774), .B2(n_775), .Y(n_773) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g732 ( .A(n_607), .Y(n_732) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_614), .B2(n_615), .Y(n_610) );
BUFx2_ASAP7_75t_R g612 ( .A(n_613), .Y(n_612) );
INVx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g785 ( .A(n_627), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_700), .B1(n_782), .B2(n_784), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g783 ( .A(n_630), .Y(n_783) );
OA22x2_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_658), .B1(n_698), .B2(n_699), .Y(n_630) );
INVx2_ASAP7_75t_L g698 ( .A(n_631), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_647), .Y(n_632) );
NOR3xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_639), .C(n_643), .Y(n_633) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_654), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_652), .Y(n_648) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_651), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx2_ASAP7_75t_L g699 ( .A(n_658), .Y(n_699) );
XOR2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_679), .Y(n_658) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_672), .Y(n_660) );
NOR3xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_665), .C(n_668), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_676), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
XOR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_697), .Y(n_679) );
NAND3x1_ASAP7_75t_L g680 ( .A(n_681), .B(n_684), .C(n_693), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NOR2x1_ASAP7_75t_L g684 ( .A(n_685), .B(n_688), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .C(n_691), .Y(n_688) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g784 ( .A(n_700), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_749), .B1(n_750), .B2(n_781), .Y(n_700) );
INVx1_ASAP7_75t_L g781 ( .A(n_701), .Y(n_781) );
OA22x2_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_720), .B2(n_748), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_702), .A2(n_703), .B1(n_751), .B2(n_752), .Y(n_750) );
INVx3_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
XOR2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_719), .Y(n_703) );
NAND3x1_ASAP7_75t_SL g704 ( .A(n_705), .B(n_708), .C(n_716), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
NOR2x1_ASAP7_75t_L g708 ( .A(n_709), .B(n_712), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .C(n_715), .Y(n_712) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g748 ( .A(n_720), .Y(n_748) );
XOR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_747), .Y(n_720) );
AND2x2_ASAP7_75t_SL g721 ( .A(n_722), .B(n_733), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_726), .C(n_729), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_738), .Y(n_733) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_741), .C(n_743), .Y(n_738) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_769), .Y(n_755) );
NOR3xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_763), .C(n_766), .Y(n_756) );
OAI22xp5_ASAP7_75t_SL g757 ( .A1(n_758), .A2(n_760), .B1(n_761), .B2(n_762), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_761), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_805) );
NOR3xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_773), .C(n_776), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .B1(n_779), .B2(n_780), .Y(n_776) );
INVx1_ASAP7_75t_L g824 ( .A(n_780), .Y(n_824) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
NOR2x1_ASAP7_75t_L g789 ( .A(n_790), .B(n_794), .Y(n_789) );
OR2x2_ASAP7_75t_SL g842 ( .A(n_790), .B(n_795), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_791), .Y(n_829) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_792), .B(n_833), .Y(n_836) );
CKINVDCx16_ASAP7_75t_R g833 ( .A(n_793), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
OAI322xp33_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_828), .A3(n_830), .B1(n_834), .B2(n_837), .C1(n_838), .C2(n_840), .Y(n_801) );
INVx1_ASAP7_75t_L g827 ( .A(n_803), .Y(n_827) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_815), .Y(n_803) );
NOR3xp33_ASAP7_75t_L g804 ( .A(n_805), .B(n_809), .C(n_812), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_816), .B(n_822), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
INVx3_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_825), .Y(n_822) );
BUFx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
CKINVDCx16_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_841), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_842), .Y(n_841) );
endmodule