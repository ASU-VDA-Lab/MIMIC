module real_aes_9192_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_691;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_753;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_224;
wire n_639;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_241;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_0), .A2(n_133), .B1(n_307), .B2(n_374), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_1), .A2(n_40), .B1(n_450), .B2(n_585), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_2), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_3), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g727 ( .A1(n_4), .A2(n_216), .B1(n_378), .B2(n_483), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_5), .A2(n_109), .B1(n_417), .B2(n_450), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_6), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_7), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_8), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_9), .A2(n_38), .B1(n_389), .B2(n_485), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_10), .A2(n_169), .B1(n_307), .B2(n_313), .Y(n_306) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_11), .A2(n_110), .B1(n_347), .B2(n_407), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_12), .A2(n_220), .B1(n_325), .B2(n_371), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_13), .A2(n_31), .B1(n_584), .B2(n_585), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_14), .A2(n_179), .B1(n_649), .B2(n_650), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_15), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_16), .A2(n_123), .B1(n_402), .B2(n_625), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_17), .A2(n_114), .B1(n_363), .B2(n_573), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_18), .Y(n_545) );
AOI22x1_ASAP7_75t_L g656 ( .A1(n_19), .A2(n_657), .B1(n_686), .B2(n_687), .Y(n_656) );
INVx1_ASAP7_75t_L g686 ( .A(n_19), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_20), .A2(n_214), .B1(n_577), .B2(n_645), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_21), .Y(n_532) );
AO22x2_ASAP7_75t_L g246 ( .A1(n_22), .A2(n_87), .B1(n_247), .B2(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g702 ( .A(n_22), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_23), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_24), .A2(n_58), .B1(n_495), .B2(n_496), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_25), .A2(n_193), .B1(n_450), .B2(n_585), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_26), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_27), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_28), .A2(n_136), .B1(n_327), .B2(n_329), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_29), .A2(n_207), .B1(n_327), .B2(n_425), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_30), .A2(n_126), .B1(n_302), .B2(n_441), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_32), .A2(n_116), .B1(n_446), .B2(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_33), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_34), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_35), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_36), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_37), .A2(n_95), .B1(n_374), .B2(n_419), .Y(n_418) );
AO22x2_ASAP7_75t_L g250 ( .A1(n_39), .A2(n_89), .B1(n_247), .B2(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g703 ( .A(n_39), .Y(n_703) );
INVx1_ASAP7_75t_L g508 ( .A(n_41), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_42), .A2(n_200), .B1(n_556), .B2(n_557), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_43), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_44), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_45), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_46), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_47), .B(n_469), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_48), .A2(n_166), .B1(n_445), .B2(n_446), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_49), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_50), .A2(n_85), .B1(n_320), .B2(n_329), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_51), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_52), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_53), .A2(n_101), .B1(n_369), .B2(n_480), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_54), .A2(n_183), .B1(n_279), .B2(n_407), .Y(n_466) );
AOI22xp33_ASAP7_75t_SL g482 ( .A1(n_55), .A2(n_186), .B1(n_378), .B2(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_56), .A2(n_112), .B1(n_477), .B2(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_57), .A2(n_73), .B1(n_367), .B2(n_370), .Y(n_366) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_59), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_60), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_61), .A2(n_83), .B1(n_272), .B2(n_279), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_62), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_63), .A2(n_115), .B1(n_358), .B2(n_363), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_64), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_65), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_66), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_67), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_68), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_69), .A2(n_177), .B1(n_500), .B2(n_501), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_70), .A2(n_176), .B1(n_409), .B2(n_411), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_71), .A2(n_217), .B1(n_556), .B2(n_649), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_72), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_74), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_75), .A2(n_96), .B1(n_503), .B2(n_504), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_76), .Y(n_589) );
AOI222xp33_ASAP7_75t_L g651 ( .A1(n_77), .A2(n_134), .B1(n_140), .B2(n_407), .C1(n_652), .C2(n_653), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_78), .Y(n_738) );
AO22x2_ASAP7_75t_L g740 ( .A1(n_78), .A2(n_738), .B1(n_741), .B2(n_761), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_79), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_80), .A2(n_181), .B1(n_585), .B2(n_757), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_81), .A2(n_82), .B1(n_318), .B2(n_329), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_84), .A2(n_125), .B1(n_348), .B2(n_352), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_86), .A2(n_158), .B1(n_417), .B2(n_649), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_88), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_90), .B(n_342), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_91), .Y(n_534) );
INVx1_ASAP7_75t_L g230 ( .A(n_92), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_93), .A2(n_203), .B1(n_553), .B2(n_554), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_94), .A2(n_161), .B1(n_503), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_97), .A2(n_160), .B1(n_504), .B2(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g226 ( .A(n_98), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_99), .A2(n_142), .B1(n_329), .B2(n_593), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_100), .A2(n_124), .B1(n_328), .B2(n_424), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_102), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_103), .A2(n_159), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_104), .A2(n_188), .B1(n_441), .B2(n_443), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_105), .A2(n_196), .B1(n_632), .B2(n_633), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_106), .A2(n_215), .B1(n_280), .B2(n_573), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_107), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_108), .B(n_471), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_111), .A2(n_113), .B1(n_419), .B2(n_639), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_117), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_118), .Y(n_679) );
XNOR2x2_ASAP7_75t_L g604 ( .A(n_119), .B(n_605), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_120), .A2(n_187), .B1(n_367), .B2(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g229 ( .A(n_121), .B(n_230), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_122), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_127), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_128), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_129), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_130), .Y(n_355) );
AND2x6_ASAP7_75t_L g225 ( .A(n_131), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_131), .Y(n_696) );
AO22x2_ASAP7_75t_L g256 ( .A1(n_132), .A2(n_178), .B1(n_247), .B2(n_251), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_135), .A2(n_155), .B1(n_318), .B2(n_322), .Y(n_317) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_137), .A2(n_191), .B1(n_350), .B2(n_629), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_138), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_139), .Y(n_464) );
INVx1_ASAP7_75t_L g331 ( .A(n_141), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_143), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_144), .A2(n_154), .B1(n_348), .B2(n_473), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_145), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_146), .B(n_350), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_147), .A2(n_163), .B1(n_328), .B2(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_148), .A2(n_204), .B1(n_650), .B2(n_760), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_149), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_150), .A2(n_171), .B1(n_347), .B2(n_350), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_151), .A2(n_221), .B1(n_477), .B2(n_478), .Y(n_476) );
AO22x2_ASAP7_75t_L g254 ( .A1(n_152), .A2(n_197), .B1(n_247), .B2(n_248), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_153), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_156), .A2(n_201), .B1(n_361), .B2(n_750), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_157), .A2(n_491), .B1(n_525), .B2(n_526), .Y(n_490) );
INVx1_ASAP7_75t_L g525 ( .A(n_157), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_162), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_164), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_165), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_167), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_168), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_170), .A2(n_706), .B1(n_707), .B2(n_729), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_170), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_172), .A2(n_202), .B1(n_299), .B2(n_302), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_173), .B(n_469), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_174), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g594 ( .A(n_175), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_178), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_180), .B(n_518), .Y(n_517) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_182), .A2(n_223), .B(n_231), .C(n_704), .Y(n_222) );
INVx1_ASAP7_75t_L g437 ( .A(n_184), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_185), .Y(n_682) );
OA22x2_ASAP7_75t_L g391 ( .A1(n_189), .A2(n_392), .B1(n_393), .B2(n_426), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_189), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_190), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_192), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_194), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_195), .Y(n_745) );
INVx1_ASAP7_75t_L g699 ( .A(n_197), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_198), .A2(n_208), .B1(n_327), .B2(n_329), .Y(n_326) );
AOI211xp5_ASAP7_75t_L g336 ( .A1(n_199), .A2(n_337), .B(n_338), .C(n_354), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_205), .Y(n_587) );
INVx1_ASAP7_75t_L g247 ( .A(n_206), .Y(n_247) );
INVx1_ASAP7_75t_L g249 ( .A(n_206), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_209), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_210), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_211), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_212), .Y(n_359) );
OA22x2_ASAP7_75t_L g561 ( .A1(n_213), .A2(n_562), .B1(n_563), .B2(n_564), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_213), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_218), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_219), .Y(n_719) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_226), .Y(n_695) );
OAI21xp5_ASAP7_75t_L g736 ( .A1(n_227), .A2(n_694), .B(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_600), .B1(n_689), .B2(n_690), .C(n_691), .Y(n_231) );
INVxp67_ASAP7_75t_L g689 ( .A(n_232), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B1(n_431), .B2(n_599), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_332), .B1(n_429), .B2(n_430), .Y(n_235) );
INVx1_ASAP7_75t_L g429 ( .A(n_236), .Y(n_429) );
XOR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_331), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_296), .Y(n_237) );
NOR3xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_263), .C(n_282), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B1(n_257), .B2(n_258), .Y(n_239) );
INVx1_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g509 ( .A(n_242), .Y(n_509) );
INVx2_ASAP7_75t_L g567 ( .A(n_242), .Y(n_567) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OAI221xp5_ASAP7_75t_L g451 ( .A1(n_243), .A2(n_260), .B1(n_452), .B2(n_453), .C(n_454), .Y(n_451) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_243), .Y(n_540) );
BUFx3_ASAP7_75t_L g712 ( .A(n_243), .Y(n_712) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_252), .Y(n_243) );
INVx2_ASAP7_75t_L g321 ( .A(n_244), .Y(n_321) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_250), .Y(n_244) );
AND2x2_ASAP7_75t_L g262 ( .A(n_245), .B(n_250), .Y(n_262) );
AND2x2_ASAP7_75t_L g301 ( .A(n_245), .B(n_277), .Y(n_301) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g268 ( .A(n_246), .B(n_250), .Y(n_268) );
AND2x2_ASAP7_75t_L g278 ( .A(n_246), .B(n_256), .Y(n_278) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g251 ( .A(n_249), .Y(n_251) );
INVx2_ASAP7_75t_L g277 ( .A(n_250), .Y(n_277) );
INVx1_ASAP7_75t_L g315 ( .A(n_250), .Y(n_315) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2x1p5_ASAP7_75t_L g261 ( .A(n_253), .B(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g325 ( .A(n_253), .B(n_301), .Y(n_325) );
AND2x4_ASAP7_75t_L g345 ( .A(n_253), .B(n_321), .Y(n_345) );
AND2x6_ASAP7_75t_L g413 ( .A(n_253), .B(n_262), .Y(n_413) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g270 ( .A(n_254), .Y(n_270) );
INVx1_ASAP7_75t_L g276 ( .A(n_254), .Y(n_276) );
INVx1_ASAP7_75t_L g295 ( .A(n_254), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_254), .B(n_256), .Y(n_305) );
AND2x2_ASAP7_75t_L g269 ( .A(n_255), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g312 ( .A(n_256), .B(n_295), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_258), .A2(n_537), .B1(n_538), .B2(n_541), .Y(n_536) );
OAI22xp5_ASAP7_75t_SL g566 ( .A1(n_258), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_258), .A2(n_538), .B1(n_675), .B2(n_676), .Y(n_674) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx3_ASAP7_75t_L g340 ( .A(n_260), .Y(n_340) );
BUFx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g512 ( .A(n_261), .Y(n_512) );
AND2x2_ASAP7_75t_L g311 ( .A(n_262), .B(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g328 ( .A(n_262), .B(n_269), .Y(n_328) );
OAI21xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B(n_271), .Y(n_263) );
BUFx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx4_ASAP7_75t_L g652 ( .A(n_266), .Y(n_652) );
OAI21xp5_ASAP7_75t_SL g715 ( .A1(n_266), .A2(n_716), .B(n_717), .Y(n_715) );
INVx4_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
BUFx3_ASAP7_75t_L g337 ( .A(n_267), .Y(n_337) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_267), .Y(n_399) );
INVx2_ASAP7_75t_SL g514 ( .A(n_267), .Y(n_514) );
INVx2_ASAP7_75t_L g622 ( .A(n_267), .Y(n_622) );
AND2x6_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx1_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
AND2x4_ASAP7_75t_L g353 ( .A(n_268), .B(n_294), .Y(n_353) );
AND2x2_ASAP7_75t_L g300 ( .A(n_269), .B(n_301), .Y(n_300) );
AND2x6_ASAP7_75t_L g320 ( .A(n_269), .B(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g396 ( .A(n_273), .Y(n_396) );
INVx4_ASAP7_75t_L g626 ( .A(n_273), .Y(n_626) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_274), .Y(n_358) );
BUFx4f_ASAP7_75t_SL g473 ( .A(n_274), .Y(n_473) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_274), .Y(n_577) );
BUFx2_ASAP7_75t_L g750 ( .A(n_274), .Y(n_750) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_278), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g281 ( .A(n_276), .Y(n_281) );
INVx1_ASAP7_75t_L g287 ( .A(n_277), .Y(n_287) );
AND2x4_ASAP7_75t_L g280 ( .A(n_278), .B(n_281), .Y(n_280) );
NAND2x1p5_ASAP7_75t_L g286 ( .A(n_278), .B(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g348 ( .A(n_278), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g519 ( .A(n_279), .Y(n_519) );
BUFx3_ASAP7_75t_L g681 ( .A(n_279), .Y(n_681) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx12f_ASAP7_75t_L g363 ( .A(n_280), .Y(n_363) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_280), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_288), .B2(n_289), .Y(n_282) );
INVx3_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g522 ( .A(n_285), .Y(n_522) );
INVx4_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx3_ASAP7_75t_L g546 ( .A(n_286), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_286), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_718) );
AND2x2_ASAP7_75t_L g446 ( .A(n_287), .B(n_304), .Y(n_446) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g524 ( .A(n_290), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g290 ( .A(n_291), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_291), .A2(n_522), .B1(n_752), .B2(n_753), .Y(n_751) );
OR2x6_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_316), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_306), .Y(n_297) );
INVx1_ASAP7_75t_L g588 ( .A(n_299), .Y(n_588) );
BUFx2_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_300), .Y(n_369) );
INVx2_ASAP7_75t_L g442 ( .A(n_300), .Y(n_442) );
AND2x4_ASAP7_75t_L g303 ( .A(n_301), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g330 ( .A(n_301), .B(n_312), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_301), .B(n_312), .Y(n_383) );
INVx1_ASAP7_75t_SL g590 ( .A(n_302), .Y(n_590) );
BUFx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
BUFx3_ASAP7_75t_L g390 ( .A(n_303), .Y(n_390) );
BUFx2_ASAP7_75t_L g417 ( .A(n_303), .Y(n_417) );
BUFx3_ASAP7_75t_L g480 ( .A(n_303), .Y(n_480) );
BUFx2_ASAP7_75t_SL g610 ( .A(n_303), .Y(n_610) );
BUFx3_ASAP7_75t_L g650 ( .A(n_303), .Y(n_650) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x6_ASAP7_75t_L g314 ( .A(n_305), .B(n_315), .Y(n_314) );
INVx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_309), .Y(n_503) );
INVx4_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx3_ASAP7_75t_L g420 ( .A(n_310), .Y(n_420) );
INVx5_ASAP7_75t_L g445 ( .A(n_310), .Y(n_445) );
INVx3_ASAP7_75t_L g483 ( .A(n_310), .Y(n_483) );
INVx1_ASAP7_75t_L g582 ( .A(n_310), .Y(n_582) );
INVx2_ASAP7_75t_L g757 ( .A(n_310), .Y(n_757) );
INVx8_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_SL g374 ( .A(n_314), .Y(n_374) );
INVx6_ASAP7_75t_SL g505 ( .A(n_314), .Y(n_505) );
INVx1_ASAP7_75t_L g349 ( .A(n_315), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_326), .Y(n_316) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx4_ASAP7_75t_L g443 ( .A(n_319), .Y(n_443) );
INVx3_ASAP7_75t_L g501 ( .A(n_319), .Y(n_501) );
INVx11_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx11_ASAP7_75t_L g372 ( .A(n_320), .Y(n_372) );
INVx4_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_323), .A2(n_614), .B1(n_615), .B2(n_616), .Y(n_613) );
INVx4_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g386 ( .A(n_325), .Y(n_386) );
BUFx3_ASAP7_75t_L g450 ( .A(n_325), .Y(n_450) );
BUFx3_ASAP7_75t_L g556 ( .A(n_325), .Y(n_556) );
BUFx3_ASAP7_75t_L g584 ( .A(n_325), .Y(n_584) );
BUFx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx6_ASAP7_75t_L g379 ( .A(n_328), .Y(n_379) );
BUFx3_ASAP7_75t_L g495 ( .A(n_328), .Y(n_495) );
BUFx3_ASAP7_75t_L g668 ( .A(n_328), .Y(n_668) );
BUFx2_ASAP7_75t_L g496 ( .A(n_329), .Y(n_496) );
BUFx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx3_ASAP7_75t_L g425 ( .A(n_330), .Y(n_425) );
BUFx3_ASAP7_75t_L g478 ( .A(n_330), .Y(n_478) );
INVx1_ASAP7_75t_L g430 ( .A(n_332), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_391), .B1(n_427), .B2(n_428), .Y(n_332) );
INVx2_ASAP7_75t_L g428 ( .A(n_333), .Y(n_428) );
XNOR2x1_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_364), .Y(n_335) );
INVx3_ASAP7_75t_L g456 ( .A(n_337), .Y(n_456) );
OAI211xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B(n_341), .C(n_346), .Y(n_338) );
BUFx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx5_ASAP7_75t_L g410 ( .A(n_344), .Y(n_410) );
INVx2_ASAP7_75t_L g469 ( .A(n_344), .Y(n_469) );
INVx2_ASAP7_75t_L g632 ( .A(n_344), .Y(n_632) );
INVx4_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g630 ( .A(n_348), .Y(n_630) );
BUFx3_ASAP7_75t_L g645 ( .A(n_348), .Y(n_645) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_SL g407 ( .A(n_353), .Y(n_407) );
BUFx2_ASAP7_75t_SL g573 ( .A(n_353), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_359), .B2(n_360), .Y(n_354) );
OAI221xp5_ASAP7_75t_L g513 ( .A1(n_356), .A2(n_514), .B1(n_515), .B2(n_516), .C(n_517), .Y(n_513) );
OAI222xp33_ASAP7_75t_L g677 ( .A1(n_356), .A2(n_398), .B1(n_678), .B2(n_679), .C1(n_680), .C2(n_682), .Y(n_677) );
INVx2_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_SL g720 ( .A(n_357), .Y(n_720) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g544 ( .A(n_358), .Y(n_544) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx4f_ASAP7_75t_SL g653 ( .A(n_363), .Y(n_653) );
NOR3xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_375), .C(n_384), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_373), .Y(n_365) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI221xp5_ASAP7_75t_SL g659 ( .A1(n_368), .A2(n_660), .B1(n_661), .B2(n_663), .C(n_664), .Y(n_659) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx3_ASAP7_75t_L g500 ( .A(n_369), .Y(n_500) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_369), .Y(n_609) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g615 ( .A(n_371), .Y(n_615) );
INVx5_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx4_ASAP7_75t_L g477 ( .A(n_372), .Y(n_477) );
INVx1_ASAP7_75t_L g593 ( .A(n_372), .Y(n_593) );
INVx2_ASAP7_75t_SL g760 ( .A(n_372), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B1(n_380), .B2(n_381), .Y(n_375) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g553 ( .A(n_379), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_379), .A2(n_596), .B1(n_618), .B2(n_619), .Y(n_617) );
INVx2_ASAP7_75t_L g639 ( .A(n_379), .Y(n_639) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g596 ( .A(n_382), .Y(n_596) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_387), .B2(n_388), .Y(n_384) );
INVx2_ASAP7_75t_L g485 ( .A(n_386), .Y(n_485) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g427 ( .A(n_391), .Y(n_427) );
INVx1_ASAP7_75t_SL g426 ( .A(n_393), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_414), .Y(n_393) );
NOR2x1_ASAP7_75t_L g394 ( .A(n_395), .B(n_405), .Y(n_394) );
OAI222xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_398), .B2(n_400), .C1(n_401), .C2(n_404), .Y(n_395) );
INVx2_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g465 ( .A(n_399), .Y(n_465) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx4f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g533 ( .A(n_403), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_408), .Y(n_405) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
BUFx4f_ASAP7_75t_L g471 ( .A(n_413), .Y(n_471) );
BUFx2_ASAP7_75t_L g633 ( .A(n_413), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_421), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
BUFx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g599 ( .A(n_431), .Y(n_599) );
AOI22xp5_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_560), .B1(n_597), .B2(n_598), .Y(n_431) );
INVx1_ASAP7_75t_L g597 ( .A(n_432), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_488), .B2(n_559), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI22xp5_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_436), .B1(n_459), .B2(n_487), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
XNOR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
NOR4xp75_ASAP7_75t_L g438 ( .A(n_439), .B(n_447), .C(n_451), .D(n_455), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_440), .B(n_444), .Y(n_439) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx3_ASAP7_75t_L g649 ( .A(n_442), .Y(n_649) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_445), .Y(n_554) );
BUFx2_ASAP7_75t_L g672 ( .A(n_445), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_448), .B(n_449), .Y(n_447) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_450), .Y(n_662) );
OAI21xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_457), .B(n_458), .Y(n_455) );
OAI21xp33_ASAP7_75t_L g570 ( .A1(n_456), .A2(n_571), .B(n_572), .Y(n_570) );
OAI21xp33_ASAP7_75t_L g747 ( .A1(n_456), .A2(n_748), .B(n_749), .Y(n_747) );
INVx2_ASAP7_75t_SL g487 ( .A(n_459), .Y(n_487) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
XOR2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_486), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_462), .B(n_474), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_467), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B(n_466), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g531 ( .A1(n_465), .A2(n_532), .B1(n_533), .B2(n_534), .C(n_535), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .C(n_472), .Y(n_467) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_481), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_479), .Y(n_475) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_480), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
INVx1_ASAP7_75t_L g559 ( .A(n_488), .Y(n_559) );
OAI22xp5_ASAP7_75t_SL g488 ( .A1(n_489), .A2(n_490), .B1(n_527), .B2(n_528), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g526 ( .A(n_491), .Y(n_526) );
AND2x2_ASAP7_75t_SL g491 ( .A(n_492), .B(n_506), .Y(n_491) );
NOR2xp33_ASAP7_75t_SL g492 ( .A(n_493), .B(n_498), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_497), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_502), .Y(n_498) );
BUFx4f_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_L g557 ( .A(n_505), .Y(n_557) );
BUFx2_ASAP7_75t_L g585 ( .A(n_505), .Y(n_585) );
BUFx2_ASAP7_75t_L g612 ( .A(n_505), .Y(n_612) );
NOR3xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_513), .C(n_520), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B1(n_510), .B2(n_511), .Y(n_507) );
OA211x2_ASAP7_75t_L g641 ( .A1(n_511), .A2(n_642), .B(n_643), .C(n_644), .Y(n_641) );
INVx1_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g714 ( .A(n_512), .Y(n_714) );
INVx2_ASAP7_75t_L g746 ( .A(n_512), .Y(n_746) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B1(n_523), .B2(n_524), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_522), .A2(n_524), .B1(n_684), .B2(n_685), .Y(n_683) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
XOR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_558), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_547), .Y(n_529) );
NOR3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .C(n_542), .Y(n_530) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_545), .B2(n_546), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_546), .A2(n_575), .B1(n_576), .B2(n_578), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx1_ASAP7_75t_SL g598 ( .A(n_560), .Y(n_598) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_579), .Y(n_564) );
NOR3xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_570), .C(n_574), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_567), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_577), .Y(n_576) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_586), .C(n_591), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B1(n_589), .B2(n_590), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI221xp5_ASAP7_75t_SL g666 ( .A1(n_596), .A2(n_667), .B1(n_669), .B2(n_670), .C(n_671), .Y(n_666) );
INVx1_ASAP7_75t_L g690 ( .A(n_600), .Y(n_690) );
AOI22xp5_ASAP7_75t_SL g600 ( .A1(n_601), .A2(n_602), .B1(n_656), .B2(n_688), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B1(n_634), .B2(n_655), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_606), .B(n_620), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_613), .C(n_617), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_627), .Y(n_620) );
OAI21xp5_ASAP7_75t_SL g621 ( .A1(n_622), .A2(n_623), .B(n_624), .Y(n_621) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g655 ( .A(n_634), .Y(n_655) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
XOR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_654), .Y(n_635) );
NAND4xp75_ASAP7_75t_L g636 ( .A(n_637), .B(n_641), .C(n_646), .D(n_651), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx2_ASAP7_75t_L g688 ( .A(n_656), .Y(n_688) );
INVx1_ASAP7_75t_SL g687 ( .A(n_657), .Y(n_687) );
AND2x2_ASAP7_75t_SL g657 ( .A(n_658), .B(n_673), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_666), .Y(n_658) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx3_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_677), .C(n_683), .Y(n_673) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
NOR2x1_ASAP7_75t_L g692 ( .A(n_693), .B(n_697), .Y(n_692) );
OR2x2_ASAP7_75t_SL g764 ( .A(n_693), .B(n_698), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_695), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_695), .B(n_734), .Y(n_737) );
CKINVDCx16_ASAP7_75t_R g734 ( .A(n_696), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
OAI322xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_730), .A3(n_731), .B1(n_735), .B2(n_738), .C1(n_739), .C2(n_762), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_707), .Y(n_706) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_722), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_715), .C(n_718), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_726), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g761 ( .A(n_741), .Y(n_761) );
AND2x2_ASAP7_75t_SL g741 ( .A(n_742), .B(n_754), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .C(n_751), .Y(n_742) );
AND4x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .C(n_758), .D(n_759), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
endmodule