module fake_jpeg_21529_n_94 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_94);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_94;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_24),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_0),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_15),
.B(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_14),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_0),
.B(n_1),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_25),
.B(n_16),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_21),
.C(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_45),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_57),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_58),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_40),
.B1(n_41),
.B2(n_35),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_52),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_16),
.B(n_29),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_21),
.B1(n_28),
.B2(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_60),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_28),
.B(n_19),
.C(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_22),
.B1(n_23),
.B2(n_20),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_2),
.B(n_3),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_20),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_45),
.C(n_53),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_73),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_53),
.C(n_55),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_70),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_74),
.B(n_66),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_44),
.B(n_43),
.Y(n_77)
);

AOI322xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_60),
.A3(n_66),
.B1(n_67),
.B2(n_52),
.C1(n_56),
.C2(n_23),
.Y(n_78)
);

OAI221xp5_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_76),
.B1(n_56),
.B2(n_18),
.C(n_13),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_73),
.C(n_74),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_81),
.C(n_69),
.Y(n_88)
);

INVxp33_ASAP7_75t_SL g83 ( 
.A(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_80),
.B(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_84),
.B(n_85),
.Y(n_86)
);

AOI32xp33_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_79),
.A3(n_81),
.B1(n_75),
.B2(n_18),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_87),
.B(n_88),
.Y(n_90)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_11),
.B(n_6),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_88),
.B(n_6),
.Y(n_91)
);

OAI321xp33_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_92),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C(n_19),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_2),
.Y(n_94)
);


endmodule