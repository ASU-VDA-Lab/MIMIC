module fake_jpeg_25369_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_39),
.Y(n_66)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_44),
.Y(n_63)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_46),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_19),
.B(n_1),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_27),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_27),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_54),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_51),
.B(n_58),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_28),
.B1(n_22),
.B2(n_30),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_53),
.A2(n_19),
.B1(n_29),
.B2(n_35),
.Y(n_116)
);

HAxp5_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_24),
.CON(n_54),
.SN(n_54)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_28),
.B1(n_23),
.B2(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_56),
.A2(n_57),
.B1(n_61),
.B2(n_29),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_28),
.B1(n_23),
.B2(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_65),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_28),
.B1(n_23),
.B2(n_22),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_22),
.B1(n_27),
.B2(n_16),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_62),
.A2(n_69),
.B1(n_74),
.B2(n_70),
.Y(n_89)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_39),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_17),
.B1(n_33),
.B2(n_16),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_20),
.B1(n_31),
.B2(n_46),
.Y(n_95)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_16),
.B1(n_31),
.B2(n_20),
.Y(n_74)
);

INVx5_ASAP7_75t_SL g75 ( 
.A(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_21),
.Y(n_97)
);

NAND2x1_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_29),
.Y(n_77)
);

NAND2x1_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_29),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_79),
.B(n_95),
.Y(n_143)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_97),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_77),
.B(n_46),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_103),
.C(n_107),
.Y(n_119)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_77),
.A2(n_33),
.B1(n_43),
.B2(n_42),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_84),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_89),
.A2(n_112),
.B1(n_63),
.B2(n_55),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_67),
.A2(n_45),
.B(n_41),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_100),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_43),
.B1(n_42),
.B2(n_32),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_94),
.A2(n_102),
.B1(n_29),
.B2(n_35),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_26),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_99),
.B(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_46),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_31),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_104),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_43),
.B1(n_32),
.B2(n_20),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_68),
.B(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_48),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_62),
.A2(n_48),
.B(n_40),
.C(n_36),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_55),
.B1(n_60),
.B2(n_65),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_48),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_40),
.Y(n_144)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_59),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_117),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_51),
.B1(n_75),
.B2(n_60),
.Y(n_121)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_121),
.A2(n_127),
.B1(n_136),
.B2(n_141),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_63),
.A3(n_50),
.B1(n_60),
.B2(n_55),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_95),
.Y(n_163)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_133),
.Y(n_149)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_134),
.A2(n_146),
.B1(n_78),
.B2(n_88),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_137),
.B(n_80),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_105),
.B(n_107),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_40),
.B1(n_36),
.B2(n_19),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_106),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_89),
.A2(n_40),
.B1(n_26),
.B2(n_21),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_153),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_100),
.C(n_82),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_158),
.C(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_151),
.B(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_107),
.B(n_82),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_155),
.A2(n_159),
.B(n_165),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_133),
.B(n_96),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_118),
.C(n_144),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_104),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_163),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_92),
.B(n_93),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_167),
.B(n_114),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_103),
.C(n_79),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_166),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_101),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_103),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_92),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_91),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_143),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_129),
.Y(n_184)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_125),
.B(n_14),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g206 ( 
.A(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_134),
.B(n_78),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_174),
.Y(n_182)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_88),
.B1(n_111),
.B2(n_110),
.Y(n_202)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_35),
.B(n_25),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_126),
.B(n_132),
.Y(n_183)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_129),
.B(n_13),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_181),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_183),
.A2(n_190),
.B1(n_202),
.B2(n_213),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_188),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_130),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_149),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_189),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_164),
.A2(n_126),
.B1(n_130),
.B2(n_117),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_139),
.C(n_124),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_197),
.C(n_198),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_139),
.C(n_124),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_86),
.C(n_109),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_171),
.C(n_153),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_86),
.C(n_25),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_159),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_166),
.B(n_128),
.CI(n_25),
.CON(n_204),
.SN(n_204)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_167),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_152),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_209),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_177),
.A2(n_145),
.B1(n_128),
.B2(n_86),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_185),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_218),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_215),
.B(n_223),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_201),
.A2(n_161),
.B(n_163),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_165),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_239),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_205),
.A2(n_177),
.B1(n_176),
.B2(n_179),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_226),
.B1(n_194),
.B2(n_204),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_153),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_228),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_189),
.B(n_148),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_167),
.B1(n_165),
.B2(n_172),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_152),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_191),
.B1(n_209),
.B2(n_210),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_128),
.C(n_9),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_233),
.C(n_187),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_9),
.C(n_13),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_192),
.B(n_14),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_185),
.B(n_1),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_193),
.B(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_238),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_187),
.B(n_12),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_240),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_240),
.A2(n_183),
.B1(n_200),
.B2(n_199),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_241),
.A2(n_249),
.B1(n_251),
.B2(n_257),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_248),
.B(n_216),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_217),
.A2(n_201),
.B1(n_182),
.B2(n_197),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_214),
.A2(n_196),
.B1(n_198),
.B2(n_194),
.Y(n_251)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_254),
.A2(n_256),
.B1(n_259),
.B2(n_237),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_221),
.A2(n_204),
.B1(n_208),
.B2(n_210),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_219),
.A2(n_235),
.B1(n_224),
.B2(n_220),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_224),
.A2(n_208),
.B1(n_191),
.B2(n_184),
.Y(n_258)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_195),
.B1(n_206),
.B2(n_5),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_12),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_233),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_262),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_229),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_268),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_271),
.B1(n_249),
.B2(n_251),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_245),
.Y(n_268)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_239),
.C(n_232),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_269),
.B(n_270),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_216),
.C(n_228),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_254),
.A2(n_236),
.B1(n_230),
.B2(n_231),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_272),
.B(n_277),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_230),
.C(n_9),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_275),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_3),
.B(n_4),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_3),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_278),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_241),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_3),
.Y(n_280)
);

XOR2x2_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_257),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_289),
.Y(n_298)
);

NOR4xp25_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_255),
.C(n_248),
.D(n_243),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_288),
.B(n_266),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_242),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_267),
.B1(n_263),
.B2(n_274),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_243),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_294),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_247),
.B1(n_262),
.B2(n_259),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_292),
.B(n_293),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_261),
.B1(n_10),
.B2(n_11),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_10),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_296),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_276),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_267),
.C(n_268),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_286),
.C(n_282),
.Y(n_307)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_304),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_280),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_303),
.B(n_279),
.Y(n_310)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_275),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_287),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_308),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_281),
.C(n_286),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_312),
.Y(n_318)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_310),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_263),
.C(n_279),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_299),
.C(n_295),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_302),
.B(n_301),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_315),
.A2(n_319),
.B(n_306),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_305),
.B(n_299),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

AOI21x1_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_10),
.B(n_11),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_322),
.Y(n_323)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

AOI322xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_316),
.A3(n_320),
.B1(n_317),
.B2(n_314),
.C1(n_12),
.C2(n_7),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_7),
.B(n_5),
.Y(n_326)
);

MAJx2_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_6),
.C(n_7),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_6),
.Y(n_328)
);


endmodule