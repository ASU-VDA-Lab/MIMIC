module fake_jpeg_17218_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_1),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_52),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_59),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_74),
.Y(n_79)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_51),
.B1(n_48),
.B2(n_43),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_50),
.B1(n_47),
.B2(n_45),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_58),
.A2(n_40),
.B1(n_43),
.B2(n_37),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_65),
.A2(n_67),
.B1(n_71),
.B2(n_46),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_37),
.B1(n_47),
.B2(n_44),
.Y(n_67)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_39),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_2),
.Y(n_85)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_85),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_63),
.C(n_50),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_90),
.C(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_36),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_42),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_84),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_86),
.B1(n_88),
.B2(n_4),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_89),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_88)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_3),
.Y(n_91)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_96),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_102),
.Y(n_105)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_79),
.C(n_86),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_103),
.B(n_101),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_88),
.B1(n_29),
.B2(n_30),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_109),
.B(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

AOI221xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.C(n_115),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_106),
.A2(n_92),
.B1(n_97),
.B2(n_96),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_108),
.A2(n_102),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_118),
.A2(n_119),
.B(n_12),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_114),
.A2(n_103),
.B1(n_107),
.B2(n_105),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_10),
.B(n_11),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_121),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_119),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_13),
.B1(n_15),
.B2(n_20),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_21),
.A3(n_25),
.B1(n_26),
.B2(n_27),
.C1(n_28),
.C2(n_31),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

XOR2x2_ASAP7_75t_R g130 ( 
.A(n_129),
.B(n_33),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_34),
.Y(n_131)
);


endmodule