module fake_netlist_1_5013_n_458 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_458);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_458;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_141;
wire n_119;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g68 ( .A(n_59), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_36), .Y(n_69) );
CKINVDCx16_ASAP7_75t_R g70 ( .A(n_55), .Y(n_70) );
CKINVDCx5p33_ASAP7_75t_R g71 ( .A(n_54), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_6), .Y(n_72) );
BUFx5_ASAP7_75t_L g73 ( .A(n_41), .Y(n_73) );
INVx2_ASAP7_75t_L g74 ( .A(n_23), .Y(n_74) );
INVx1_ASAP7_75t_SL g75 ( .A(n_42), .Y(n_75) );
INVx1_ASAP7_75t_SL g76 ( .A(n_63), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_31), .Y(n_77) );
BUFx6f_ASAP7_75t_L g78 ( .A(n_13), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_7), .Y(n_79) );
BUFx3_ASAP7_75t_L g80 ( .A(n_12), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_47), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_29), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_11), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_35), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_67), .Y(n_85) );
INVx3_ASAP7_75t_L g86 ( .A(n_51), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_65), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_49), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_53), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_34), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_12), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_62), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_56), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_64), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_43), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_7), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_60), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_27), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_61), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_2), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_66), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_58), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_9), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_26), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_19), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_68), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_70), .Y(n_107) );
INVx3_ASAP7_75t_L g108 ( .A(n_86), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_80), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_68), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_70), .B(n_0), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_89), .B(n_0), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_86), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_71), .Y(n_114) );
NOR2xp67_ASAP7_75t_L g115 ( .A(n_86), .B(n_1), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_69), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_72), .B(n_79), .Y(n_117) );
AND2x2_ASAP7_75t_SL g118 ( .A(n_69), .B(n_28), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_80), .B(n_1), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_77), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_86), .Y(n_121) );
CKINVDCx14_ASAP7_75t_R g122 ( .A(n_84), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_80), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_73), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_74), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_95), .B(n_2), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_93), .B(n_3), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_113), .B(n_93), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_113), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_109), .B(n_96), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_109), .B(n_96), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_113), .Y(n_132) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_107), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_113), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_111), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_123), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_108), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_108), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_122), .B(n_94), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_108), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_126), .Y(n_141) );
BUFx2_ASAP7_75t_L g142 ( .A(n_123), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_108), .Y(n_143) );
BUFx6f_ASAP7_75t_SL g144 ( .A(n_118), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_108), .B(n_72), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_121), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_124), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_126), .B(n_79), .Y(n_148) );
OR2x2_ASAP7_75t_SL g149 ( .A(n_117), .B(n_83), .Y(n_149) );
OAI221xp5_ASAP7_75t_L g150 ( .A1(n_117), .A2(n_105), .B1(n_91), .B2(n_103), .C(n_100), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_108), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_129), .Y(n_152) );
NOR2xp33_ASAP7_75t_R g153 ( .A(n_136), .B(n_107), .Y(n_153) );
NAND3xp33_ASAP7_75t_SL g154 ( .A(n_135), .B(n_114), .C(n_111), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_131), .B(n_111), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_131), .B(n_122), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g157 ( .A1(n_142), .A2(n_118), .B1(n_100), .B2(n_105), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_137), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_145), .B(n_112), .Y(n_159) );
OR2x6_ASAP7_75t_L g160 ( .A(n_141), .B(n_148), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_145), .B(n_112), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_137), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
INVx2_ASAP7_75t_SL g164 ( .A(n_148), .Y(n_164) );
INVx5_ASAP7_75t_L g165 ( .A(n_141), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
NOR2xp33_ASAP7_75t_R g167 ( .A(n_144), .B(n_118), .Y(n_167) );
INVx1_ASAP7_75t_SL g168 ( .A(n_142), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_148), .B(n_112), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_146), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
NOR3xp33_ASAP7_75t_SL g174 ( .A(n_150), .B(n_127), .C(n_91), .Y(n_174) );
BUFx8_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
BUFx4f_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
OR2x2_ASAP7_75t_L g177 ( .A(n_149), .B(n_119), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_146), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_139), .Y(n_180) );
NOR3xp33_ASAP7_75t_SL g181 ( .A(n_149), .B(n_127), .C(n_83), .Y(n_181) );
NOR2xp33_ASAP7_75t_R g182 ( .A(n_144), .B(n_118), .Y(n_182) );
OAI22xp33_ASAP7_75t_L g183 ( .A1(n_163), .A2(n_141), .B1(n_144), .B2(n_128), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_159), .B(n_130), .Y(n_184) );
INVx5_ASAP7_75t_L g185 ( .A(n_160), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_158), .Y(n_186) );
OR2x6_ASAP7_75t_SL g187 ( .A(n_175), .B(n_97), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_158), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_159), .B(n_130), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_162), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_162), .Y(n_192) );
INVx3_ASAP7_75t_SL g193 ( .A(n_168), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_165), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_157), .A2(n_141), .B1(n_130), .B2(n_126), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_170), .B(n_126), .Y(n_197) );
OR2x2_ASAP7_75t_L g198 ( .A(n_163), .B(n_128), .Y(n_198) );
O2A1O1Ixp5_ASAP7_75t_SL g199 ( .A1(n_166), .A2(n_125), .B(n_77), .C(n_81), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_166), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_170), .A2(n_151), .B1(n_143), .B2(n_119), .Y(n_201) );
OAI22xp5_ASAP7_75t_SL g202 ( .A1(n_180), .A2(n_103), .B1(n_104), .B2(n_85), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_167), .A2(n_126), .B1(n_119), .B2(n_151), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_165), .Y(n_205) );
NAND3xp33_ASAP7_75t_L g206 ( .A(n_174), .B(n_134), .C(n_147), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_169), .A2(n_132), .B(n_129), .Y(n_207) );
CKINVDCx11_ASAP7_75t_R g208 ( .A(n_160), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_170), .B(n_126), .Y(n_209) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_160), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_170), .B(n_115), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_204), .A2(n_176), .B1(n_120), .B2(n_106), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_198), .B(n_155), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_197), .A2(n_182), .B1(n_176), .B2(n_154), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_186), .Y(n_215) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_183), .A2(n_115), .B(n_120), .Y(n_216) );
OAI221xp5_ASAP7_75t_L g217 ( .A1(n_195), .A2(n_156), .B1(n_181), .B2(n_155), .C(n_177), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_186), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_198), .A2(n_164), .B1(n_177), .B2(n_160), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_188), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_188), .A2(n_120), .B1(n_106), .B2(n_110), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_190), .Y(n_222) );
NAND3xp33_ASAP7_75t_L g223 ( .A(n_199), .B(n_110), .C(n_116), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_190), .Y(n_224) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_207), .A2(n_116), .B(n_74), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_189), .B(n_161), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_193), .B(n_165), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_192), .A2(n_169), .B(n_178), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_200), .Y(n_229) );
AOI22xp33_ASAP7_75t_SL g230 ( .A1(n_185), .A2(n_153), .B1(n_175), .B2(n_116), .Y(n_230) );
NAND2x1_ASAP7_75t_L g231 ( .A(n_203), .B(n_172), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_197), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_197), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_209), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_209), .A2(n_175), .B1(n_165), .B2(n_178), .Y(n_235) );
OAI221xp5_ASAP7_75t_L g236 ( .A1(n_202), .A2(n_173), .B1(n_152), .B2(n_82), .C(n_90), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_212), .A2(n_208), .B1(n_211), .B2(n_209), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_217), .A2(n_208), .B1(n_211), .B2(n_189), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_215), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_215), .Y(n_240) );
AOI22xp33_ASAP7_75t_SL g241 ( .A1(n_219), .A2(n_185), .B1(n_175), .B2(n_187), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_215), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_220), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_213), .B(n_184), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_226), .B(n_185), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_220), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_212), .A2(n_187), .B1(n_185), .B2(n_201), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_236), .A2(n_211), .B1(n_210), .B2(n_206), .Y(n_248) );
AOI21x1_ASAP7_75t_L g249 ( .A1(n_225), .A2(n_121), .B(n_171), .Y(n_249) );
OR2x2_ASAP7_75t_L g250 ( .A(n_222), .B(n_191), .Y(n_250) );
OAI221xp5_ASAP7_75t_L g251 ( .A1(n_214), .A2(n_203), .B1(n_205), .B2(n_196), .C(n_121), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_222), .Y(n_252) );
OAI221xp5_ASAP7_75t_L g253 ( .A1(n_230), .A2(n_205), .B1(n_196), .B2(n_121), .C(n_125), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_222), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_226), .B(n_194), .Y(n_255) );
AOI21x1_ASAP7_75t_L g256 ( .A1(n_225), .A2(n_223), .B(n_231), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_238), .A2(n_234), .B1(n_233), .B2(n_232), .Y(n_257) );
INVx4_ASAP7_75t_R g258 ( .A(n_239), .Y(n_258) );
NOR4xp25_ASAP7_75t_SL g259 ( .A(n_253), .B(n_102), .C(n_90), .D(n_98), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_240), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_247), .A2(n_221), .B1(n_224), .B2(n_229), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_240), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_240), .Y(n_263) );
OAI221xp5_ASAP7_75t_L g264 ( .A1(n_241), .A2(n_235), .B1(n_234), .B2(n_233), .C(n_232), .Y(n_264) );
NAND2xp33_ASAP7_75t_R g265 ( .A(n_239), .B(n_227), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_246), .B(n_224), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_242), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_242), .B(n_224), .Y(n_268) );
NAND2xp33_ASAP7_75t_R g269 ( .A(n_243), .B(n_225), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_244), .B(n_218), .Y(n_270) );
INVx4_ASAP7_75t_L g271 ( .A(n_246), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_243), .Y(n_272) );
AOI322xp5_ASAP7_75t_L g273 ( .A1(n_237), .A2(n_125), .A3(n_92), .B1(n_102), .B2(n_101), .C1(n_98), .C2(n_81), .Y(n_273) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_256), .A2(n_223), .B(n_228), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_245), .A2(n_216), .B1(n_229), .B2(n_225), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_246), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_267), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_267), .Y(n_278) );
NOR3xp33_ASAP7_75t_L g279 ( .A(n_264), .B(n_251), .C(n_101), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_266), .B(n_252), .Y(n_280) );
OAI221xp5_ASAP7_75t_L g281 ( .A1(n_257), .A2(n_248), .B1(n_254), .B2(n_252), .C(n_255), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_271), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_260), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_260), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_272), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_262), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_272), .B(n_254), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g288 ( .A1(n_270), .A2(n_78), .B1(n_255), .B2(n_125), .C(n_87), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_263), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_269), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_266), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_258), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_268), .B(n_252), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_263), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_266), .B(n_250), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_268), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_266), .A2(n_216), .B(n_250), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_271), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_271), .Y(n_299) );
NOR3xp33_ASAP7_75t_L g300 ( .A(n_261), .B(n_87), .C(n_88), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_276), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_276), .B(n_256), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_275), .B(n_216), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_299), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_280), .B(n_274), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_283), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_283), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_277), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_282), .B(n_261), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_286), .B(n_274), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_277), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_280), .B(n_274), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_304), .B(n_274), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_299), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_278), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_283), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_304), .B(n_73), .Y(n_318) );
CKINVDCx8_ASAP7_75t_R g319 ( .A(n_292), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_296), .B(n_4), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_284), .Y(n_321) );
AOI31xp33_ASAP7_75t_L g322 ( .A1(n_292), .A2(n_265), .A3(n_258), .B(n_88), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_285), .B(n_273), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_284), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_292), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_285), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_284), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_295), .B(n_73), .Y(n_328) );
AO22x1_ASAP7_75t_L g329 ( .A1(n_290), .A2(n_92), .B1(n_78), .B2(n_95), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_286), .B(n_78), .Y(n_330) );
NOR4xp25_ASAP7_75t_SL g331 ( .A(n_281), .B(n_99), .C(n_259), .D(n_8), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_287), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_293), .B(n_78), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_293), .B(n_78), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_282), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_302), .B(n_291), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_282), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_287), .B(n_125), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_289), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_289), .Y(n_340) );
NOR4xp25_ASAP7_75t_SL g341 ( .A(n_294), .B(n_5), .C(n_6), .D(n_8), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_294), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_309), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_315), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_310), .A2(n_300), .B1(n_279), .B2(n_288), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_318), .B(n_297), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_318), .B(n_297), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_305), .B(n_302), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_328), .B(n_298), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_315), .B(n_298), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_332), .B(n_303), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_335), .B(n_301), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_312), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_325), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g355 ( .A1(n_320), .A2(n_95), .B1(n_76), .B2(n_75), .C(n_124), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_332), .B(n_73), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_335), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_336), .B(n_73), .Y(n_358) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_330), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_316), .B(n_73), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_326), .B(n_73), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_322), .A2(n_249), .B1(n_205), .B2(n_191), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_308), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_339), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_333), .B(n_5), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_310), .A2(n_73), .B1(n_194), .B2(n_146), .Y(n_366) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_329), .A2(n_337), .B(n_333), .C(n_310), .Y(n_367) );
AOI21xp33_ASAP7_75t_SL g368 ( .A1(n_329), .A2(n_10), .B(n_11), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_319), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_340), .B(n_249), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_310), .A2(n_194), .B1(n_146), .B2(n_171), .Y(n_371) );
AOI31xp33_ASAP7_75t_L g372 ( .A1(n_319), .A2(n_13), .A3(n_14), .B(n_15), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_308), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_308), .Y(n_374) );
A2O1A1Ixp33_ASAP7_75t_L g375 ( .A1(n_323), .A2(n_15), .B(n_16), .C(n_17), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_342), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_334), .Y(n_377) );
AOI21xp33_ASAP7_75t_L g378 ( .A1(n_372), .A2(n_338), .B(n_311), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_351), .B(n_311), .Y(n_379) );
NOR2xp33_ASAP7_75t_R g380 ( .A(n_369), .B(n_345), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_351), .B(n_314), .Y(n_381) );
NAND2xp33_ASAP7_75t_L g382 ( .A(n_369), .B(n_317), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_358), .B(n_314), .Y(n_383) );
INVx1_ASAP7_75t_SL g384 ( .A(n_354), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_364), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_343), .Y(n_386) );
NOR4xp25_ASAP7_75t_SL g387 ( .A(n_368), .B(n_341), .C(n_331), .D(n_19), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_376), .B(n_306), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_359), .B(n_306), .Y(n_389) );
OAI21xp5_ASAP7_75t_SL g390 ( .A1(n_362), .A2(n_313), .B(n_317), .Y(n_390) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_367), .B(n_341), .C(n_331), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_350), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_346), .B(n_313), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_346), .B(n_327), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_347), .B(n_324), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_347), .B(n_324), .Y(n_397) );
INVxp67_ASAP7_75t_L g398 ( .A(n_344), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g399 ( .A(n_356), .B(n_321), .C(n_307), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_363), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_373), .Y(n_401) );
NOR3xp33_ASAP7_75t_SL g402 ( .A(n_375), .B(n_18), .C(n_20), .Y(n_402) );
AOI21xp33_ASAP7_75t_L g403 ( .A1(n_356), .A2(n_307), .B(n_22), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_352), .B(n_21), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_360), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_352), .B(n_374), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_360), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_361), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_379), .Y(n_409) );
OAI31xp33_ASAP7_75t_L g410 ( .A1(n_390), .A2(n_357), .A3(n_365), .B(n_361), .Y(n_410) );
NAND4xp25_ASAP7_75t_L g411 ( .A(n_378), .B(n_355), .C(n_366), .D(n_349), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_379), .Y(n_412) );
NOR2xp33_ASAP7_75t_SL g413 ( .A(n_384), .B(n_348), .Y(n_413) );
INVx2_ASAP7_75t_SL g414 ( .A(n_392), .Y(n_414) );
O2A1O1Ixp5_ASAP7_75t_L g415 ( .A1(n_389), .A2(n_377), .B(n_370), .C(n_371), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_386), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_393), .B(n_370), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_386), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_385), .Y(n_419) );
NAND4xp25_ASAP7_75t_L g420 ( .A(n_391), .B(n_179), .C(n_147), .D(n_132), .Y(n_420) );
XNOR2xp5_ASAP7_75t_L g421 ( .A(n_381), .B(n_24), .Y(n_421) );
XOR2xp5_ASAP7_75t_L g422 ( .A(n_383), .B(n_25), .Y(n_422) );
OAI21xp33_ASAP7_75t_SL g423 ( .A1(n_381), .A2(n_30), .B(n_32), .Y(n_423) );
A2O1A1Ixp33_ASAP7_75t_SL g424 ( .A1(n_387), .A2(n_147), .B(n_37), .C(n_38), .Y(n_424) );
O2A1O1Ixp33_ASAP7_75t_L g425 ( .A1(n_402), .A2(n_33), .B(n_39), .C(n_40), .Y(n_425) );
OAI21xp33_ASAP7_75t_SL g426 ( .A1(n_398), .A2(n_44), .B(n_45), .Y(n_426) );
OAI32xp33_ASAP7_75t_L g427 ( .A1(n_399), .A2(n_46), .A3(n_48), .B1(n_50), .B2(n_52), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_394), .A2(n_146), .B1(n_129), .B2(n_57), .Y(n_428) );
INVx3_ASAP7_75t_SL g429 ( .A(n_414), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_409), .B(n_397), .Y(n_430) );
OAI211xp5_ASAP7_75t_L g431 ( .A1(n_423), .A2(n_380), .B(n_408), .C(n_407), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g432 ( .A1(n_410), .A2(n_405), .B1(n_394), .B2(n_395), .C(n_388), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_417), .B(n_395), .Y(n_433) );
OAI21xp33_ASAP7_75t_L g434 ( .A1(n_413), .A2(n_406), .B(n_382), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_416), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_417), .B(n_396), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_418), .Y(n_437) );
NOR2xp67_ASAP7_75t_L g438 ( .A(n_426), .B(n_400), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_411), .A2(n_404), .B1(n_401), .B2(n_403), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_419), .Y(n_440) );
OAI311xp33_ASAP7_75t_L g441 ( .A1(n_420), .A2(n_425), .A3(n_428), .B1(n_415), .C1(n_422), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_427), .A2(n_423), .B(n_410), .Y(n_442) );
XNOR2x2_ASAP7_75t_L g443 ( .A(n_424), .B(n_421), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_413), .A2(n_411), .B1(n_412), .B2(n_409), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_409), .B(n_412), .Y(n_445) );
OR3x2_ASAP7_75t_L g446 ( .A(n_443), .B(n_441), .C(n_442), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_444), .B(n_432), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_438), .A2(n_429), .B1(n_431), .B2(n_434), .Y(n_448) );
OAI322xp33_ASAP7_75t_L g449 ( .A1(n_439), .A2(n_445), .A3(n_440), .B1(n_436), .B2(n_433), .C1(n_435), .C2(n_437), .Y(n_449) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_430), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_450), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_446), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_447), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_452), .B(n_448), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_451), .Y(n_455) );
OR3x2_ASAP7_75t_L g456 ( .A(n_454), .B(n_453), .C(n_449), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_456), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_457), .A2(n_453), .B(n_455), .Y(n_458) );
endmodule