module fake_jpeg_5771_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_43),
.Y(n_51)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_18),
.Y(n_54)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_19),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_22),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_16),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_46),
.B(n_49),
.C(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_71),
.B(n_72),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_19),
.B1(n_33),
.B2(n_23),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_73),
.A2(n_77),
.B1(n_78),
.B2(n_90),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_75),
.B(n_95),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_76),
.Y(n_124)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_19),
.B1(n_33),
.B2(n_23),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_33),
.B(n_22),
.C(n_30),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_84),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_24),
.B1(n_18),
.B2(n_25),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_92),
.B1(n_30),
.B2(n_32),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_38),
.B(n_37),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_94),
.B(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_34),
.Y(n_89)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_33),
.B1(n_23),
.B2(n_29),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_53),
.A2(n_47),
.B(n_56),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_34),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_32),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_23),
.B1(n_30),
.B2(n_52),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_109),
.B1(n_110),
.B2(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_101),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_21),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_112),
.B1(n_96),
.B2(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_21),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_108),
.Y(n_135)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_64),
.B(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_32),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_29),
.B1(n_37),
.B2(n_38),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_24),
.B1(n_25),
.B2(n_18),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_21),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_52),
.Y(n_115)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_58),
.B1(n_27),
.B2(n_28),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_63),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_58),
.Y(n_120)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_80),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_126),
.B1(n_91),
.B2(n_24),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_82),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_93),
.Y(n_152)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_132),
.Y(n_168)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_79),
.B(n_98),
.C(n_85),
.D(n_96),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_130),
.B(n_107),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_97),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_74),
.C(n_72),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_155),
.C(n_115),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_112),
.A2(n_74),
.B1(n_68),
.B2(n_77),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_90),
.B1(n_73),
.B2(n_78),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_157),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_68),
.B1(n_77),
.B2(n_80),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_144),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_141),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_103),
.A2(n_119),
.B1(n_109),
.B2(n_110),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_106),
.B(n_113),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_143),
.A2(n_147),
.B(n_107),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g146 ( 
.A(n_127),
.Y(n_146)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_96),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_156),
.Y(n_161)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_154),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_86),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_70),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_76),
.C(n_70),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_31),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_102),
.A2(n_91),
.B1(n_25),
.B2(n_28),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_120),
.B(n_105),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_128),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_163),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_155),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_14),
.Y(n_209)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_177),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_176),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_124),
.C(n_105),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_187),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_113),
.B1(n_126),
.B2(n_102),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_189),
.B1(n_131),
.B2(n_17),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_171),
.A2(n_129),
.B1(n_132),
.B2(n_137),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_107),
.Y(n_178)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_179),
.B(n_183),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_153),
.A2(n_127),
.B1(n_116),
.B2(n_123),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_180),
.A2(n_191),
.B1(n_7),
.B2(n_13),
.Y(n_205)
);

AO22x2_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_104),
.B1(n_111),
.B2(n_27),
.Y(n_181)
);

AO22x2_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_31),
.Y(n_182)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_31),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_130),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_192),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_93),
.Y(n_186)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_93),
.C(n_31),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_26),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_147),
.A2(n_26),
.B1(n_31),
.B2(n_17),
.Y(n_189)
);

BUFx24_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_17),
.B(n_1),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_0),
.Y(n_192)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_150),
.A3(n_135),
.B1(n_142),
.B2(n_139),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_171),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_213),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_200),
.A2(n_209),
.B(n_191),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_193),
.A2(n_17),
.B1(n_9),
.B2(n_10),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_216),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_7),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_217),
.C(n_221),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_205),
.A2(n_222),
.B1(n_181),
.B2(n_184),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_219),
.Y(n_229)
);

OAI21x1_ASAP7_75t_R g211 ( 
.A1(n_160),
.A2(n_0),
.B(n_1),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_212),
.B1(n_181),
.B2(n_164),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_176),
.Y(n_213)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_161),
.B(n_13),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_168),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_170),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_161),
.B(n_13),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_166),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_222)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_165),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_223),
.B(n_224),
.Y(n_249)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_225),
.B(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_220),
.A2(n_166),
.B1(n_178),
.B2(n_172),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_230),
.A2(n_239),
.B1(n_215),
.B2(n_190),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_233),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_159),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_167),
.C(n_169),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_210),
.C(n_202),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_237),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_216),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_187),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_244),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_200),
.A2(n_181),
.B1(n_183),
.B2(n_179),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_207),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_242),
.A2(n_245),
.B(n_223),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_212),
.A2(n_181),
.B1(n_189),
.B2(n_162),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_243),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_182),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_160),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_204),
.B(n_190),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_212),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_252),
.C(n_258),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_221),
.C(n_195),
.Y(n_252)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_239),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_218),
.C(n_214),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_224),
.A2(n_212),
.B1(n_208),
.B2(n_162),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_268),
.B1(n_230),
.B2(n_231),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_264),
.C(n_265),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_263),
.A2(n_245),
.B1(n_234),
.B2(n_228),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_175),
.C(n_2),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_1),
.Y(n_266)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_11),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_228),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_256),
.A2(n_246),
.B1(n_236),
.B2(n_240),
.Y(n_270)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_273),
.B(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_276),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_243),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_278),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_279),
.A2(n_282),
.B(n_285),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_248),
.B(n_245),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_284),
.Y(n_293)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_255),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_258),
.C(n_254),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_292),
.C(n_295),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_288),
.A2(n_298),
.B(n_279),
.Y(n_302)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_250),
.B(n_251),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_249),
.B(n_4),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_254),
.C(n_252),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_267),
.C(n_265),
.Y(n_295)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

INVx11_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_268),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_281),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_289),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_302),
.A2(n_303),
.B(n_304),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_287),
.B(n_264),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_297),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_293),
.Y(n_306)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_272),
.Y(n_307)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

OAI21x1_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_249),
.B(n_276),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_12),
.C1(n_301),
.C2(n_310),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_247),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_309),
.A2(n_294),
.B(n_295),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_SL g312 ( 
.A1(n_310),
.A2(n_291),
.B(n_288),
.C(n_6),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_314),
.C(n_317),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_11),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_315),
.Y(n_325)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_3),
.A3(n_12),
.B1(n_302),
.B2(n_309),
.C1(n_300),
.C2(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_316),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_305),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_323),
.B(n_324),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_3),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_312),
.Y(n_327)
);

OAI21xp33_ASAP7_75t_SL g330 ( 
.A1(n_327),
.A2(n_329),
.B(n_321),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_312),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_330),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_328),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_325),
.Y(n_333)
);


endmodule