module fake_ariane_452_n_2038 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2038);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2038;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_355;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1856;
wire n_2016;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx10_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_120),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_52),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_182),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_63),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_29),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_160),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_49),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_194),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_3),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_112),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_18),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_150),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_93),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_118),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_177),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_121),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_61),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_174),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_11),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_168),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_133),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_105),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_33),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_95),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_142),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_113),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_12),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_80),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_18),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_137),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_83),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_109),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_159),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_127),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_61),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_101),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_9),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_77),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_13),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_166),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_12),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_25),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_22),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_161),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_1),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_91),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_16),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_2),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_132),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_149),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_128),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_131),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_115),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_169),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_76),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_81),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_92),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_22),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_147),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_98),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_136),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_73),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_8),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_191),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_70),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_55),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_178),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_193),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_78),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_123),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_42),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_157),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_171),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_107),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_49),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_96),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_5),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_28),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_79),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_154),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_26),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_190),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_53),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_87),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_148),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_184),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_68),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_82),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_13),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_11),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_165),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_85),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_117),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_100),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_15),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_179),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_3),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_43),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_2),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_36),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_126),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_90),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_46),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_8),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_33),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_124),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_72),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_158),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_102),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_134),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_145),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_152),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_24),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_172),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_114),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_67),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_141),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_40),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_0),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_163),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_64),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_94),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_106),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_14),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_60),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_59),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_24),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_7),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_200),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_84),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_48),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_104),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_43),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_58),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_41),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_36),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_162),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_10),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_99),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_26),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_188),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_138),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_16),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_139),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_156),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_46),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_103),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_1),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_7),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_129),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_71),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_9),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_0),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_48),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_189),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_44),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_122),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_40),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_42),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_23),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_196),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_35),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_69),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_35),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_86),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_140),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_50),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_119),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_45),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_6),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_180),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_5),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_67),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_45),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_181),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_41),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_14),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_27),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_47),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_108),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_30),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_58),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_10),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_28),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_75),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_97),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_183),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_130),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_6),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_203),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_224),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_335),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_258),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_335),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_278),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_387),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_283),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_318),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_368),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_372),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_387),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_231),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_274),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_387),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_220),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_382),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_277),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_268),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_244),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_247),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_337),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_249),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_359),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_220),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_252),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_294),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_349),
.B(n_4),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_294),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_330),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_386),
.B(n_4),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_330),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_363),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_360),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_285),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_201),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_259),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_286),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_360),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_289),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_201),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_292),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_298),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_371),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_201),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_218),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_390),
.Y(n_453)
);

INVxp33_ASAP7_75t_SL g454 ( 
.A(n_209),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_400),
.B(n_15),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_306),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_218),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_271),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_271),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_399),
.B(n_17),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_268),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_205),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_221),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_308),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_209),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_310),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_314),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_210),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_238),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_296),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_327),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_254),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_216),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_256),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_221),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_221),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_296),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_269),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_282),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_329),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_288),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_243),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_215),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_332),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_336),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_354),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_215),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_300),
.Y(n_488)
);

NOR2xp67_ASAP7_75t_L g489 ( 
.A(n_311),
.B(n_17),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_315),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_316),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_339),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_364),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_202),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_346),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_357),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_216),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_365),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_367),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_370),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_243),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_424),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_497),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_483),
.B(n_206),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_403),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_482),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_405),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_482),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_404),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_404),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_470),
.B(n_375),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_483),
.B(n_207),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_482),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_406),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_406),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_421),
.B(n_383),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_470),
.B(n_384),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_482),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_482),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_407),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_453),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_407),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_455),
.A2(n_324),
.B1(n_214),
.B2(n_309),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_420),
.B(n_212),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_410),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_410),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_415),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_409),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_415),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_409),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_416),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_416),
.Y(n_533)
);

INVxp33_ASAP7_75t_SL g534 ( 
.A(n_426),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_419),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_424),
.B(n_461),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_425),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_419),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_432),
.B(n_388),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_452),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_452),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_457),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_457),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_423),
.A2(n_226),
.B1(n_228),
.B2(n_232),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_458),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_465),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_458),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_501),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_459),
.A2(n_246),
.B(n_234),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_459),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_494),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_494),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_487),
.B(n_501),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_461),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_487),
.B(n_260),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_430),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_430),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_434),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_434),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_435),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_435),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_439),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_439),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_454),
.B(n_436),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_444),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_444),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_449),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_449),
.Y(n_568)
);

BUFx8_ASAP7_75t_L g569 ( 
.A(n_455),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_450),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_450),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_462),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_462),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_500),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_500),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_473),
.Y(n_576)
);

OA21x2_ASAP7_75t_L g577 ( 
.A1(n_468),
.A2(n_272),
.B(n_264),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_468),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_437),
.B(n_273),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_469),
.Y(n_580)
);

OA21x2_ASAP7_75t_L g581 ( 
.A1(n_469),
.A2(n_290),
.B(n_287),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_502),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_553),
.B(n_417),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_502),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_531),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_531),
.Y(n_586)
);

INVx4_ASAP7_75t_SL g587 ( 
.A(n_551),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_506),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_548),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_531),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_548),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_506),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_505),
.B(n_417),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_510),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_524),
.A2(n_478),
.B1(n_342),
.B2(n_253),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_504),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_508),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_553),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_531),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_505),
.B(n_428),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_548),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_536),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_551),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_532),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_536),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_532),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_513),
.B(n_431),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_510),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_572),
.B(n_481),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_551),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_513),
.B(n_442),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_532),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_572),
.B(n_472),
.Y(n_613)
);

NOR2x1p5_ASAP7_75t_L g614 ( 
.A(n_555),
.B(n_443),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_534),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_551),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_569),
.A2(n_460),
.B1(n_489),
.B2(n_433),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_578),
.B(n_243),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_578),
.B(n_472),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_511),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_541),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_580),
.B(n_474),
.Y(n_622)
);

AND2x6_ASAP7_75t_L g623 ( 
.A(n_580),
.B(n_243),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_569),
.A2(n_489),
.B1(n_433),
.B2(n_477),
.Y(n_624)
);

BUFx8_ASAP7_75t_SL g625 ( 
.A(n_504),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_548),
.B(n_445),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_532),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_L g628 ( 
.A(n_555),
.B(n_250),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_541),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_564),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_541),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_511),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_515),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_503),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_551),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_551),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_569),
.A2(n_394),
.B1(n_395),
.B2(n_389),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_517),
.B(n_474),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_541),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_564),
.A2(n_548),
.B1(n_546),
.B2(n_569),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_503),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_504),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_541),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_541),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_503),
.B(n_447),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_577),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_509),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_569),
.A2(n_446),
.B1(n_475),
.B2(n_441),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_503),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_577),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_524),
.A2(n_476),
.B1(n_463),
.B2(n_451),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_515),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_516),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_573),
.Y(n_654)
);

OR2x6_ASAP7_75t_L g655 ( 
.A(n_544),
.B(n_479),
.Y(n_655)
);

BUFx4f_ASAP7_75t_L g656 ( 
.A(n_577),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_573),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_508),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_573),
.Y(n_659)
);

BUFx4f_ASAP7_75t_L g660 ( 
.A(n_577),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_573),
.B(n_250),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_517),
.B(n_479),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_554),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_541),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_522),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_551),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_551),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_546),
.B(n_456),
.C(n_448),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_534),
.A2(n_464),
.B1(n_498),
.B2(n_466),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_522),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_574),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_525),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_577),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_541),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_577),
.A2(n_492),
.B1(n_467),
.B2(n_480),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_517),
.A2(n_471),
.B1(n_484),
.B2(n_485),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_539),
.A2(n_486),
.B1(n_493),
.B2(n_373),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_537),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_539),
.B(n_440),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_574),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_537),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_574),
.B(n_488),
.Y(n_682)
);

CKINVDCx6p67_ASAP7_75t_R g683 ( 
.A(n_576),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_543),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_574),
.B(n_488),
.Y(n_685)
);

INVx6_ASAP7_75t_L g686 ( 
.A(n_512),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_543),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_581),
.A2(n_499),
.B1(n_496),
.B2(n_495),
.Y(n_688)
);

OR2x6_ASAP7_75t_L g689 ( 
.A(n_544),
.B(n_499),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_554),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_543),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_576),
.B(n_418),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_516),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_525),
.B(n_579),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_512),
.B(n_518),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_543),
.Y(n_696)
);

INVx4_ASAP7_75t_L g697 ( 
.A(n_581),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_543),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_543),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_543),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_539),
.B(n_401),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_521),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_543),
.Y(n_703)
);

INVx8_ASAP7_75t_L g704 ( 
.A(n_512),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_509),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_554),
.B(n_490),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_554),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_554),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_547),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_575),
.B(n_490),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_581),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_547),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_581),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_547),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_579),
.Y(n_715)
);

INVxp67_ASAP7_75t_SL g716 ( 
.A(n_552),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_540),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_512),
.B(n_408),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_552),
.B(n_491),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_521),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_523),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_523),
.Y(n_722)
);

OR2x6_ASAP7_75t_L g723 ( 
.A(n_512),
.B(n_491),
.Y(n_723)
);

NAND3xp33_ASAP7_75t_L g724 ( 
.A(n_581),
.B(n_228),
.C(n_226),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_581),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_547),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_549),
.Y(n_727)
);

NAND2xp33_ASAP7_75t_L g728 ( 
.A(n_575),
.B(n_250),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_518),
.B(n_575),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_575),
.B(n_495),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_518),
.A2(n_236),
.B1(n_232),
.B2(n_301),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_518),
.B(n_411),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_549),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_SL g734 ( 
.A(n_518),
.B(n_413),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_694),
.B(n_557),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_676),
.B(n_630),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_585),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_630),
.B(n_414),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_630),
.B(n_600),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_672),
.B(n_557),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_582),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_602),
.B(n_557),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_605),
.B(n_557),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_585),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_583),
.A2(n_422),
.B1(n_540),
.B2(n_542),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_607),
.B(n_557),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_611),
.B(n_717),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_591),
.B(n_204),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_593),
.B(n_402),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_591),
.B(n_204),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_L g751 ( 
.A(n_589),
.B(n_250),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_717),
.B(n_638),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_638),
.B(n_552),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_638),
.B(n_552),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_586),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_591),
.B(n_208),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_662),
.B(n_542),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_586),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_662),
.B(n_545),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_662),
.B(n_545),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_609),
.B(n_550),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_609),
.B(n_550),
.Y(n_762)
);

NAND2xp33_ASAP7_75t_L g763 ( 
.A(n_589),
.B(n_250),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_613),
.B(n_556),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_704),
.B(n_556),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_678),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_582),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_626),
.B(n_208),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_669),
.B(n_211),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_613),
.B(n_559),
.Y(n_770)
);

O2A1O1Ixp5_ASAP7_75t_L g771 ( 
.A1(n_603),
.A2(n_559),
.B(n_570),
.C(n_561),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_692),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_619),
.B(n_561),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_590),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_622),
.B(n_566),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_SL g776 ( 
.A1(n_715),
.A2(n_427),
.B1(n_429),
.B2(n_438),
.Y(n_776)
);

AO221x1_ASAP7_75t_L g777 ( 
.A1(n_595),
.A2(n_362),
.B1(n_356),
.B2(n_243),
.C(n_352),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_640),
.A2(n_338),
.B1(n_393),
.B2(n_301),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_692),
.B(n_567),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_723),
.B(n_570),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_590),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_665),
.B(n_412),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_665),
.B(n_236),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_725),
.A2(n_549),
.B1(n_547),
.B2(n_565),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_601),
.B(n_558),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_601),
.B(n_211),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_725),
.A2(n_549),
.B1(n_350),
.B2(n_213),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_645),
.B(n_558),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_677),
.B(n_213),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_584),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_682),
.B(n_558),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_682),
.B(n_558),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_584),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_R g794 ( 
.A(n_615),
.B(n_217),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_598),
.B(n_217),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_685),
.B(n_562),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_599),
.Y(n_797)
);

NAND3xp33_ASAP7_75t_L g798 ( 
.A(n_675),
.B(n_668),
.C(n_658),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_598),
.B(n_219),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_617),
.A2(n_549),
.B1(n_353),
.B2(n_219),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_685),
.B(n_562),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_588),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_598),
.B(n_222),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_599),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_710),
.B(n_562),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_615),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_588),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_673),
.B(n_250),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_681),
.B(n_222),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_715),
.A2(n_549),
.B1(n_547),
.B2(n_565),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_597),
.B(n_223),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_723),
.B(n_496),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_604),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_724),
.A2(n_547),
.B1(n_565),
.B2(n_563),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_701),
.B(n_338),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_597),
.B(n_223),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_658),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_604),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_670),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_710),
.B(n_730),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_670),
.B(n_562),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_637),
.B(n_225),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_606),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_730),
.B(n_568),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_606),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_729),
.B(n_568),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_704),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_612),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_718),
.B(n_679),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_656),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_729),
.B(n_568),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_704),
.Y(n_832)
);

NOR2x1_ASAP7_75t_L g833 ( 
.A(n_614),
.B(n_241),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_704),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_729),
.B(n_568),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_592),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_592),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_628),
.A2(n_519),
.B(n_514),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_688),
.B(n_571),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_594),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_612),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_716),
.B(n_571),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_663),
.B(n_571),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_673),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_718),
.B(n_225),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_734),
.B(n_227),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_627),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_594),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_663),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_732),
.B(n_344),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_656),
.A2(n_351),
.B1(n_344),
.B2(n_345),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_596),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_723),
.B(n_571),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_690),
.B(n_707),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_624),
.B(n_227),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_690),
.B(n_707),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_642),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_608),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_723),
.B(n_560),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_627),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_654),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_708),
.B(n_560),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_608),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_708),
.B(n_560),
.Y(n_864)
);

NAND2xp33_ASAP7_75t_SL g865 ( 
.A(n_646),
.B(n_345),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_656),
.B(n_229),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_660),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_634),
.B(n_560),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_620),
.A2(n_538),
.B(n_529),
.C(n_533),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_620),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_657),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_632),
.B(n_560),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_632),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_633),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_633),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_652),
.B(n_560),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_683),
.B(n_347),
.Y(n_877)
);

NAND2xp33_ASAP7_75t_L g878 ( 
.A(n_713),
.B(n_250),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_660),
.B(n_229),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_625),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_652),
.B(n_560),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_653),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_653),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_693),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_659),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_693),
.B(n_560),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_702),
.B(n_563),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_702),
.B(n_563),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_628),
.A2(n_340),
.B1(n_341),
.B2(n_398),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_720),
.B(n_721),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_660),
.A2(n_547),
.B1(n_565),
.B2(n_563),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_671),
.Y(n_892)
);

NAND2xp33_ASAP7_75t_L g893 ( 
.A(n_713),
.B(n_250),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_720),
.B(n_563),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_721),
.B(n_563),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_686),
.B(n_347),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_686),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_722),
.A2(n_538),
.B(n_535),
.C(n_533),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_722),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_680),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_641),
.Y(n_901)
);

AOI221xp5_ASAP7_75t_L g902 ( 
.A1(n_731),
.A2(n_351),
.B1(n_392),
.B2(n_393),
.C(n_380),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_686),
.Y(n_903)
);

OR2x2_ASAP7_75t_SL g904 ( 
.A(n_655),
.B(n_689),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_751),
.A2(n_733),
.B(n_610),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_737),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_747),
.B(n_686),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_751),
.A2(n_733),
.B(n_610),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_759),
.B(n_683),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_759),
.B(n_695),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_766),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_760),
.B(n_695),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_763),
.A2(n_610),
.B(n_603),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_812),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_777),
.A2(n_655),
.B1(n_689),
.B2(n_727),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_763),
.A2(n_616),
.B(n_603),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_830),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_735),
.A2(n_635),
.B(n_616),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_771),
.A2(n_650),
.B(n_646),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_741),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_746),
.A2(n_635),
.B(n_616),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_829),
.B(n_655),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_760),
.B(n_695),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_827),
.B(n_695),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_821),
.B(n_706),
.Y(n_925)
);

AOI21x1_ASAP7_75t_L g926 ( 
.A1(n_839),
.A2(n_649),
.B(n_643),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_827),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_890),
.A2(n_636),
.B(n_635),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_834),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_834),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_741),
.Y(n_931)
);

NOR3xp33_ASAP7_75t_L g932 ( 
.A(n_736),
.B(n_378),
.C(n_369),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_812),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_820),
.A2(n_719),
.B(n_655),
.C(n_689),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_844),
.A2(n_788),
.B(n_785),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_737),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_780),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_821),
.B(n_689),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_767),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_767),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_830),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_744),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_740),
.A2(n_864),
.B(n_862),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_749),
.B(n_727),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_739),
.B(n_727),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_812),
.B(n_646),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_790),
.Y(n_947)
);

OAI21xp33_ASAP7_75t_L g948 ( 
.A1(n_783),
.A2(n_392),
.B(n_385),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_742),
.A2(n_666),
.B(n_636),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_832),
.B(n_650),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_L g951 ( 
.A(n_832),
.B(n_621),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_806),
.Y(n_952)
);

OAI21xp33_ASAP7_75t_L g953 ( 
.A1(n_902),
.A2(n_381),
.B(n_651),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_772),
.B(n_648),
.Y(n_954)
);

OAI321xp33_ASAP7_75t_L g955 ( 
.A1(n_778),
.A2(n_529),
.A3(n_535),
.B1(n_297),
.B2(n_376),
.C(n_303),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_817),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_790),
.A2(n_728),
.B(n_661),
.C(n_674),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_743),
.A2(n_697),
.B(n_650),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_838),
.A2(n_643),
.B(n_639),
.Y(n_959)
);

INVx11_ASAP7_75t_L g960 ( 
.A(n_852),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_765),
.B(n_697),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_752),
.B(n_697),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_843),
.A2(n_868),
.B(n_856),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_744),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_891),
.A2(n_711),
.B(n_664),
.Y(n_965)
);

NOR3xp33_ASAP7_75t_L g966 ( 
.A(n_738),
.B(n_674),
.C(n_661),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_761),
.B(n_762),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_764),
.A2(n_728),
.B(n_674),
.C(n_712),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_782),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_872),
.A2(n_711),
.B(n_664),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_836),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_757),
.B(n_711),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_854),
.A2(n_666),
.B(n_636),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_819),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_830),
.B(n_621),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_808),
.A2(n_667),
.B(n_666),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_770),
.B(n_773),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_808),
.A2(n_667),
.B(n_639),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_SL g979 ( 
.A1(n_748),
.A2(n_684),
.B(n_714),
.C(n_712),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_878),
.A2(n_667),
.B(n_684),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_876),
.A2(n_691),
.B(n_687),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_780),
.B(n_621),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_836),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_755),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_837),
.A2(n_691),
.B(n_714),
.C(n_696),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_878),
.A2(n_698),
.B(n_696),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_775),
.A2(n_703),
.B(n_700),
.C(n_698),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_837),
.A2(n_699),
.B1(n_700),
.B2(n_703),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_893),
.A2(n_629),
.B(n_621),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_840),
.A2(n_726),
.B(n_709),
.C(n_621),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_893),
.A2(n_631),
.B(n_629),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_857),
.B(n_625),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_791),
.A2(n_527),
.B(n_528),
.C(n_304),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_780),
.B(n_824),
.Y(n_994)
);

BUFx12f_ASAP7_75t_L g995 ( 
.A(n_806),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_881),
.A2(n_631),
.B(n_629),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_758),
.Y(n_997)
);

NAND2xp33_ASAP7_75t_L g998 ( 
.A(n_840),
.B(n_629),
.Y(n_998)
);

OAI21xp33_ASAP7_75t_L g999 ( 
.A1(n_794),
.A2(n_233),
.B(n_230),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_848),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_758),
.Y(n_1001)
);

INVx4_ASAP7_75t_L g1002 ( 
.A(n_765),
.Y(n_1002)
);

OAI321xp33_ASAP7_75t_L g1003 ( 
.A1(n_800),
.A2(n_305),
.A3(n_307),
.B1(n_313),
.B2(n_320),
.C(n_325),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_848),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_779),
.Y(n_1005)
);

O2A1O1Ixp5_ASAP7_75t_L g1006 ( 
.A1(n_866),
.A2(n_507),
.B(n_519),
.C(n_514),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_886),
.A2(n_631),
.B(n_629),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_858),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_858),
.Y(n_1009)
);

NOR2xp67_ASAP7_75t_SL g1010 ( 
.A(n_795),
.B(n_631),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_887),
.A2(n_644),
.B(n_631),
.Y(n_1011)
);

BUFx4f_ASAP7_75t_L g1012 ( 
.A(n_765),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_888),
.A2(n_709),
.B(n_644),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_776),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_779),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_894),
.A2(n_709),
.B(n_644),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_863),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_897),
.B(n_903),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_824),
.B(n_644),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_895),
.A2(n_705),
.B(n_647),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_896),
.B(n_644),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_877),
.B(n_563),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_753),
.B(n_709),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_754),
.B(n_709),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_792),
.A2(n_705),
.B(n_647),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_879),
.A2(n_726),
.B(n_705),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_796),
.A2(n_726),
.B(n_705),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_801),
.A2(n_726),
.B(n_705),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_805),
.A2(n_647),
.B(n_507),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_870),
.A2(n_874),
.B(n_875),
.C(n_873),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_853),
.B(n_726),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_853),
.B(n_793),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_877),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_880),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_765),
.B(n_563),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_833),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_842),
.A2(n_647),
.B(n_519),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_904),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_861),
.A2(n_647),
.B(n_507),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_802),
.B(n_565),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_786),
.A2(n_514),
.B(n_519),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_870),
.A2(n_528),
.B(n_527),
.C(n_377),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_897),
.B(n_230),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_798),
.B(n_565),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_774),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_903),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_830),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_807),
.B(n_565),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_873),
.B(n_565),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_874),
.B(n_875),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_882),
.B(n_587),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_882),
.A2(n_884),
.B(n_883),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_883),
.B(n_587),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_904),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_859),
.B(n_587),
.Y(n_1055)
);

NOR2xp67_ASAP7_75t_L g1056 ( 
.A(n_745),
.B(n_527),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_884),
.A2(n_514),
.B(n_507),
.Y(n_1057)
);

NAND2x1p5_ASAP7_75t_L g1058 ( 
.A(n_859),
.B(n_527),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_899),
.A2(n_379),
.B(n_527),
.C(n_528),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_899),
.A2(n_507),
.B(n_239),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_826),
.B(n_587),
.Y(n_1061)
);

O2A1O1Ixp5_ASAP7_75t_L g1062 ( 
.A1(n_865),
.A2(n_528),
.B(n_530),
.C(n_618),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_781),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_768),
.A2(n_240),
.B(n_239),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_831),
.B(n_233),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_861),
.A2(n_240),
.B(n_237),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_835),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_871),
.A2(n_237),
.B(n_235),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_871),
.A2(n_340),
.B(n_341),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_815),
.B(n_528),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_867),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_781),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_849),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_851),
.B(n_343),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_885),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_885),
.A2(n_343),
.B(n_348),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_892),
.A2(n_348),
.B(n_350),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_867),
.B(n_353),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_810),
.B(n_355),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_892),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_900),
.A2(n_355),
.B(n_358),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_845),
.B(n_618),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_850),
.B(n_358),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_849),
.Y(n_1084)
);

AND2x2_ASAP7_75t_SL g1085 ( 
.A(n_787),
.B(n_352),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_849),
.B(n_901),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_869),
.A2(n_530),
.B(n_242),
.C(n_251),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_811),
.B(n_816),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_797),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_750),
.A2(n_391),
.B(n_396),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_922),
.A2(n_865),
.B(n_846),
.C(n_898),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_977),
.A2(n_756),
.B(n_799),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_1002),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_935),
.A2(n_803),
.B(n_860),
.Y(n_1094)
);

AO21x1_ASAP7_75t_L g1095 ( 
.A1(n_944),
.A2(n_855),
.B(n_789),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_998),
.A2(n_818),
.B(n_860),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_967),
.A2(n_970),
.B(n_1052),
.Y(n_1097)
);

NOR2xp67_ASAP7_75t_L g1098 ( 
.A(n_952),
.B(n_809),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1015),
.B(n_769),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_969),
.A2(n_822),
.B(n_847),
.C(n_841),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_929),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_956),
.Y(n_1102)
);

BUFx4_ASAP7_75t_SL g1103 ( 
.A(n_1034),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_994),
.B(n_797),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_905),
.A2(n_818),
.B(n_847),
.Y(n_1105)
);

BUFx5_ASAP7_75t_L g1106 ( 
.A(n_961),
.Y(n_1106)
);

BUFx12f_ASAP7_75t_L g1107 ( 
.A(n_995),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_922),
.B(n_804),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_908),
.A2(n_823),
.B(n_841),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_963),
.A2(n_828),
.B(n_825),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1075),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_1005),
.B(n_804),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_943),
.A2(n_828),
.B(n_825),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_976),
.A2(n_823),
.B(n_813),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_906),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1005),
.B(n_969),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_909),
.B(n_889),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_1002),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_913),
.A2(n_813),
.B(n_784),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1085),
.A2(n_814),
.B1(n_398),
.B2(n_397),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_914),
.B(n_777),
.Y(n_1121)
);

CKINVDCx16_ASAP7_75t_R g1122 ( 
.A(n_992),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_914),
.B(n_933),
.Y(n_1123)
);

INVx8_ASAP7_75t_L g1124 ( 
.A(n_1035),
.Y(n_1124)
);

CKINVDCx8_ASAP7_75t_R g1125 ( 
.A(n_1038),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_960),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_933),
.B(n_391),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_916),
.A2(n_317),
.B(n_248),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_SL g1129 ( 
.A(n_934),
.B(n_932),
.C(n_1083),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_911),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_938),
.B(n_396),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1067),
.B(n_1032),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1067),
.B(n_397),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_937),
.B(n_245),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_948),
.A2(n_530),
.B(n_20),
.C(n_21),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1085),
.A2(n_530),
.B1(n_321),
.B2(n_366),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_956),
.B(n_526),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1080),
.Y(n_1138)
);

NAND2x1p5_ASAP7_75t_L g1139 ( 
.A(n_937),
.B(n_1012),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1012),
.B(n_255),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_924),
.B(n_257),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1050),
.B(n_526),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_929),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_924),
.B(n_261),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_920),
.A2(n_302),
.B1(n_299),
.B2(n_295),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_929),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_931),
.B(n_526),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1054),
.B(n_1055),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_939),
.A2(n_293),
.B1(n_291),
.B2(n_284),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_936),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_940),
.B(n_947),
.Y(n_1151)
);

NAND2x1_ASAP7_75t_L g1152 ( 
.A(n_1047),
.B(n_618),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_1033),
.A2(n_267),
.B1(n_266),
.B2(n_265),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_942),
.Y(n_1154)
);

NAND2x1p5_ASAP7_75t_L g1155 ( 
.A(n_917),
.B(n_526),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1025),
.A2(n_328),
.B(n_263),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_971),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_983),
.B(n_526),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_929),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_964),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1000),
.B(n_526),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_944),
.B(n_19),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1004),
.A2(n_1008),
.B1(n_1017),
.B2(n_1009),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1021),
.A2(n_331),
.B(n_270),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_930),
.B(n_262),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_910),
.B(n_19),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_953),
.A2(n_623),
.B1(n_618),
.B2(n_333),
.Y(n_1167)
);

AOI21x1_ASAP7_75t_L g1168 ( 
.A1(n_959),
.A2(n_526),
.B(n_623),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1089),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1030),
.A2(n_276),
.B1(n_275),
.B2(n_279),
.Y(n_1170)
);

AOI22x1_ASAP7_75t_L g1171 ( 
.A1(n_918),
.A2(n_526),
.B1(n_281),
.B2(n_280),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_974),
.B(n_312),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_958),
.A2(n_319),
.B(n_322),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1089),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_984),
.Y(n_1175)
);

BUFx12f_ASAP7_75t_L g1176 ( 
.A(n_1036),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_974),
.B(n_374),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_934),
.A2(n_1074),
.B(n_932),
.C(n_1088),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_954),
.B(n_1088),
.Y(n_1179)
);

CKINVDCx16_ASAP7_75t_R g1180 ( 
.A(n_1014),
.Y(n_1180)
);

AND2x2_ASAP7_75t_SL g1181 ( 
.A(n_915),
.B(n_362),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_925),
.B(n_623),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_997),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_912),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_930),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_923),
.B(n_25),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1087),
.A2(n_361),
.B(n_326),
.C(n_334),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_930),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_930),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1001),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_917),
.B(n_323),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_919),
.A2(n_623),
.B(n_618),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_961),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1022),
.B(n_27),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_915),
.A2(n_362),
.B1(n_356),
.B2(n_352),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_999),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_951),
.A2(n_991),
.B(n_989),
.Y(n_1197)
);

AOI21x1_ASAP7_75t_L g1198 ( 
.A1(n_926),
.A2(n_975),
.B(n_1010),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1078),
.A2(n_31),
.B(n_32),
.C(n_34),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1046),
.B(n_945),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1058),
.B(n_32),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1045),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_921),
.A2(n_362),
.B(n_356),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1063),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_917),
.B(n_520),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1046),
.B(n_34),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_945),
.B(n_37),
.Y(n_1207)
);

CKINVDCx14_ASAP7_75t_R g1208 ( 
.A(n_1035),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1072),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_SL g1210 ( 
.A1(n_1035),
.A2(n_1082),
.B1(n_1058),
.B2(n_1065),
.Y(n_1210)
);

AND2x4_ASAP7_75t_SL g1211 ( 
.A(n_927),
.B(n_356),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_978),
.A2(n_352),
.B(n_520),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1040),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_1031),
.Y(n_1214)
);

AO32x2_ASAP7_75t_L g1215 ( 
.A1(n_988),
.A2(n_37),
.A3(n_38),
.B1(n_39),
.B2(n_44),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1018),
.B(n_39),
.Y(n_1216)
);

NOR3xp33_ASAP7_75t_SL g1217 ( 
.A(n_1064),
.B(n_47),
.C(n_50),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1087),
.A2(n_352),
.B(n_520),
.C(n_509),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1048),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1049),
.Y(n_1220)
);

OR2x6_ASAP7_75t_SL g1221 ( 
.A(n_907),
.B(n_1079),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1019),
.A2(n_972),
.B1(n_957),
.B2(n_1086),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_917),
.B(n_520),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1073),
.B(n_51),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_R g1225 ( 
.A(n_927),
.B(n_941),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_962),
.A2(n_990),
.B1(n_982),
.B2(n_1024),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1071),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1071),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_SL g1229 ( 
.A1(n_966),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1071),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_980),
.A2(n_520),
.B(n_509),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1055),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1071),
.B(n_520),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1020),
.A2(n_520),
.B(n_509),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_R g1235 ( 
.A(n_941),
.B(n_110),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1070),
.B(n_54),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_955),
.A2(n_520),
.B(n_509),
.C(n_56),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1073),
.B(n_54),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1056),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1084),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_941),
.B(n_509),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_SL g1242 ( 
.A1(n_950),
.A2(n_55),
.B(n_56),
.C(n_57),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1003),
.A2(n_509),
.B(n_59),
.C(n_60),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1044),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_949),
.A2(n_125),
.B(n_198),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_941),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_996),
.A2(n_111),
.B(n_195),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1162),
.A2(n_1043),
.B1(n_1084),
.B2(n_1023),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1179),
.B(n_1090),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1130),
.Y(n_1250)
);

BUFx5_ASAP7_75t_L g1251 ( 
.A(n_1220),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1116),
.B(n_1044),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1115),
.Y(n_1253)
);

OA21x2_ASAP7_75t_L g1254 ( 
.A1(n_1097),
.A2(n_1212),
.B(n_1203),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1197),
.A2(n_968),
.B(n_965),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1117),
.B(n_1082),
.Y(n_1256)
);

BUFx8_ASAP7_75t_SL g1257 ( 
.A(n_1107),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1103),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1207),
.A2(n_968),
.B(n_928),
.Y(n_1259)
);

OR2x6_ASAP7_75t_L g1260 ( 
.A(n_1124),
.B(n_946),
.Y(n_1260)
);

AOI21xp33_ASAP7_75t_L g1261 ( 
.A1(n_1178),
.A2(n_993),
.B(n_987),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1222),
.A2(n_1027),
.B(n_1028),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1181),
.A2(n_1081),
.B1(n_1077),
.B2(n_1076),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1222),
.A2(n_987),
.B(n_1053),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1150),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1131),
.A2(n_966),
.B1(n_1047),
.B2(n_975),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1101),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1168),
.A2(n_986),
.B(n_1011),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_SL g1269 ( 
.A1(n_1091),
.A2(n_1059),
.B(n_1051),
.C(n_985),
.Y(n_1269)
);

BUFx10_ASAP7_75t_L g1270 ( 
.A(n_1126),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_1195),
.A2(n_1061),
.A3(n_1007),
.B(n_1013),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1094),
.A2(n_1016),
.B(n_1029),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1226),
.A2(n_979),
.B(n_973),
.Y(n_1273)
);

AOI21x1_ASAP7_75t_SL g1274 ( 
.A1(n_1238),
.A2(n_1060),
.B(n_1006),
.Y(n_1274)
);

NOR4xp25_ASAP7_75t_L g1275 ( 
.A(n_1129),
.B(n_1042),
.C(n_993),
.D(n_981),
.Y(n_1275)
);

INVx8_ASAP7_75t_L g1276 ( 
.A(n_1176),
.Y(n_1276)
);

AOI221xp5_ASAP7_75t_SL g1277 ( 
.A1(n_1199),
.A2(n_1069),
.B1(n_1068),
.B2(n_1066),
.C(n_1042),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1226),
.A2(n_1039),
.B(n_1026),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_SL g1279 ( 
.A1(n_1238),
.A2(n_1057),
.B(n_1041),
.C(n_1037),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1180),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1111),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1154),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1102),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1142),
.A2(n_1006),
.B(n_1062),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1172),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1092),
.A2(n_1062),
.B(n_62),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1160),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1138),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1110),
.A2(n_89),
.B(n_187),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1132),
.B(n_57),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1173),
.A2(n_62),
.B(n_63),
.Y(n_1291)
);

OR2x6_ASAP7_75t_L g1292 ( 
.A(n_1124),
.B(n_64),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1113),
.A2(n_143),
.B(n_175),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1195),
.A2(n_135),
.A3(n_167),
.B(n_155),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1157),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1169),
.B(n_1174),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1119),
.A2(n_88),
.A3(n_146),
.B(n_144),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1139),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1136),
.A2(n_1237),
.B(n_1135),
.C(n_1187),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1125),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1122),
.B(n_65),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1142),
.A2(n_74),
.B(n_199),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1099),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1114),
.A2(n_65),
.B(n_66),
.Y(n_1304)
);

AO21x1_ASAP7_75t_L g1305 ( 
.A1(n_1136),
.A2(n_66),
.B(n_68),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1200),
.A2(n_1120),
.B(n_1156),
.Y(n_1306)
);

AOI31xp67_ASAP7_75t_L g1307 ( 
.A1(n_1241),
.A2(n_1233),
.A3(n_1230),
.B(n_1228),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1163),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1112),
.B(n_1151),
.Y(n_1309)
);

OAI22x1_ASAP7_75t_L g1310 ( 
.A1(n_1239),
.A2(n_1144),
.B1(n_1141),
.B2(n_1193),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1177),
.A2(n_1210),
.B1(n_1120),
.B2(n_1098),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1243),
.A2(n_1196),
.B(n_1218),
.C(n_1100),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1216),
.A2(n_1108),
.B(n_1244),
.C(n_1184),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1101),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1231),
.A2(n_1105),
.B(n_1109),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1236),
.A2(n_1186),
.B(n_1166),
.C(n_1217),
.Y(n_1316)
);

AO21x1_ASAP7_75t_L g1317 ( 
.A1(n_1170),
.A2(n_1163),
.B(n_1121),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1096),
.A2(n_1192),
.B(n_1234),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1151),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1192),
.A2(n_1213),
.B(n_1219),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1148),
.Y(n_1321)
);

INVxp67_ASAP7_75t_SL g1322 ( 
.A(n_1123),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1214),
.B(n_1148),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_1227),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_SL g1325 ( 
.A1(n_1229),
.A2(n_1191),
.B(n_1224),
.C(n_1134),
.Y(n_1325)
);

NOR2x1_ASAP7_75t_SL g1326 ( 
.A(n_1101),
.B(n_1185),
.Y(n_1326)
);

AOI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1198),
.A2(n_1182),
.B(n_1223),
.Y(n_1327)
);

A2O1A1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1206),
.A2(n_1194),
.B(n_1164),
.C(n_1128),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1202),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1245),
.A2(n_1161),
.B(n_1158),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1104),
.A2(n_1133),
.B(n_1140),
.C(n_1167),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1214),
.B(n_1232),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1188),
.Y(n_1333)
);

AO21x1_ASAP7_75t_L g1334 ( 
.A1(n_1147),
.A2(n_1158),
.B(n_1161),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1204),
.A2(n_1175),
.A3(n_1209),
.B(n_1190),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1147),
.A2(n_1247),
.B(n_1205),
.Y(n_1336)
);

INVxp67_ASAP7_75t_SL g1337 ( 
.A(n_1232),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1171),
.A2(n_1152),
.B(n_1155),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1124),
.A2(n_1211),
.B(n_1240),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1155),
.A2(n_1093),
.B(n_1118),
.Y(n_1340)
);

AO21x2_ASAP7_75t_L g1341 ( 
.A1(n_1183),
.A2(n_1165),
.B(n_1235),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1137),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1153),
.A2(n_1149),
.A3(n_1145),
.B(n_1159),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1225),
.Y(n_1344)
);

AO21x2_ASAP7_75t_L g1345 ( 
.A1(n_1242),
.A2(n_1127),
.B(n_1149),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_SL g1346 ( 
.A1(n_1139),
.A2(n_1246),
.B(n_1185),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1143),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1221),
.B(n_1106),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1215),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1106),
.B(n_1201),
.Y(n_1350)
);

AOI221x1_ASAP7_75t_L g1351 ( 
.A1(n_1145),
.A2(n_1093),
.B1(n_1118),
.B2(n_1246),
.C(n_1159),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1208),
.A2(n_1246),
.B(n_1143),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1143),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1106),
.A2(n_1146),
.B(n_1185),
.Y(n_1354)
);

OAI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1146),
.A2(n_1189),
.B1(n_1215),
.B2(n_1106),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1189),
.A2(n_922),
.B1(n_969),
.B2(n_1162),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1215),
.B(n_1106),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1189),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1195),
.A2(n_1119),
.A3(n_1095),
.B(n_1218),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1195),
.A2(n_1119),
.A3(n_1095),
.B(n_1218),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1157),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1115),
.Y(n_1362)
);

A2O1A1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1178),
.A2(n_934),
.B(n_922),
.C(n_1207),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1207),
.A2(n_944),
.B(n_607),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1195),
.A2(n_1119),
.A3(n_1095),
.B(n_1218),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1097),
.A2(n_998),
.B(n_763),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1097),
.A2(n_998),
.B(n_763),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1157),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1097),
.A2(n_998),
.B(n_763),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1179),
.B(n_1012),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1162),
.A2(n_922),
.B1(n_969),
.B2(n_1207),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1111),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1097),
.A2(n_1212),
.B(n_1203),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1179),
.B(n_1005),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1162),
.A2(n_922),
.B1(n_969),
.B2(n_1207),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1179),
.B(n_1005),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1232),
.B(n_937),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1097),
.A2(n_998),
.B(n_763),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1207),
.A2(n_944),
.B(n_607),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1097),
.A2(n_998),
.B(n_763),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1097),
.A2(n_998),
.B(n_763),
.Y(n_1381)
);

AO22x2_ASAP7_75t_L g1382 ( 
.A1(n_1195),
.A2(n_1136),
.B1(n_1120),
.B2(n_1129),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1115),
.Y(n_1383)
);

O2A1O1Ixp5_ASAP7_75t_L g1384 ( 
.A1(n_1207),
.A2(n_1162),
.B(n_1095),
.C(n_944),
.Y(n_1384)
);

NAND2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1130),
.B(n_937),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1097),
.A2(n_998),
.B(n_763),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1168),
.A2(n_959),
.B(n_1110),
.Y(n_1387)
);

BUFx10_ASAP7_75t_L g1388 ( 
.A(n_1126),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1115),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1179),
.B(n_1116),
.Y(n_1390)
);

BUFx10_ASAP7_75t_L g1391 ( 
.A(n_1126),
.Y(n_1391)
);

AOI221xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1199),
.A2(n_948),
.B1(n_969),
.B2(n_564),
.C(n_1207),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1179),
.B(n_1005),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1130),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1168),
.A2(n_959),
.B(n_1110),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1179),
.B(n_1015),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1123),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1111),
.Y(n_1398)
);

AO31x2_ASAP7_75t_L g1399 ( 
.A1(n_1195),
.A2(n_1119),
.A3(n_1095),
.B(n_1218),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1178),
.A2(n_934),
.B(n_922),
.C(n_1207),
.Y(n_1400)
);

INVx5_ASAP7_75t_L g1401 ( 
.A(n_1124),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_SL g1402 ( 
.A1(n_1162),
.A2(n_1091),
.B(n_739),
.C(n_1030),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1207),
.A2(n_944),
.B(n_607),
.Y(n_1403)
);

AOI221x1_ASAP7_75t_L g1404 ( 
.A1(n_1195),
.A2(n_1136),
.B1(n_1120),
.B2(n_1129),
.C(n_1207),
.Y(n_1404)
);

BUFx4_ASAP7_75t_SL g1405 ( 
.A(n_1126),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1130),
.Y(n_1406)
);

CKINVDCx16_ASAP7_75t_R g1407 ( 
.A(n_1107),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1130),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1097),
.A2(n_998),
.B(n_763),
.Y(n_1409)
);

AND2x6_ASAP7_75t_L g1410 ( 
.A(n_1093),
.B(n_961),
.Y(n_1410)
);

AOI221x1_ASAP7_75t_L g1411 ( 
.A1(n_1195),
.A2(n_1136),
.B1(n_1120),
.B2(n_1129),
.C(n_1207),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1179),
.A2(n_922),
.B1(n_782),
.B2(n_749),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1405),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1283),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1296),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1412),
.A2(n_1375),
.B1(n_1371),
.B2(n_1382),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1382),
.A2(n_1364),
.B1(n_1379),
.B2(n_1403),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1295),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1324),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_SL g1420 ( 
.A1(n_1256),
.A2(n_1249),
.B1(n_1291),
.B2(n_1306),
.Y(n_1420)
);

OAI22x1_ASAP7_75t_L g1421 ( 
.A1(n_1311),
.A2(n_1285),
.B1(n_1301),
.B2(n_1348),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1305),
.A2(n_1317),
.B1(n_1390),
.B2(n_1393),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1276),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1353),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1309),
.Y(n_1425)
);

BUFx8_ASAP7_75t_L g1426 ( 
.A(n_1344),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1374),
.A2(n_1376),
.B1(n_1303),
.B2(n_1252),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1363),
.A2(n_1400),
.B1(n_1316),
.B2(n_1308),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1361),
.Y(n_1429)
);

INVx3_ASAP7_75t_SL g1430 ( 
.A(n_1280),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1368),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1394),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1406),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1319),
.A2(n_1292),
.B1(n_1349),
.B2(n_1396),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1370),
.A2(n_1356),
.B1(n_1292),
.B2(n_1310),
.Y(n_1435)
);

BUFx8_ASAP7_75t_SL g1436 ( 
.A(n_1257),
.Y(n_1436)
);

CKINVDCx6p67_ASAP7_75t_R g1437 ( 
.A(n_1407),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1321),
.B(n_1408),
.Y(n_1438)
);

OAI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1404),
.A2(n_1411),
.B1(n_1290),
.B2(n_1319),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1267),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1281),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1281),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1258),
.Y(n_1443)
);

CKINVDCx11_ASAP7_75t_R g1444 ( 
.A(n_1270),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1385),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1288),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1288),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1366),
.A2(n_1378),
.B(n_1409),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1372),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1372),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1345),
.A2(n_1397),
.B1(n_1322),
.B2(n_1398),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1323),
.B(n_1332),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1270),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1250),
.A2(n_1350),
.B1(n_1266),
.B2(n_1260),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1398),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1357),
.A2(n_1342),
.B1(n_1263),
.B2(n_1355),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1335),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1261),
.A2(n_1341),
.B1(n_1286),
.B2(n_1253),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1341),
.A2(n_1248),
.B1(n_1259),
.B2(n_1410),
.Y(n_1459)
);

CKINVDCx11_ASAP7_75t_R g1460 ( 
.A(n_1388),
.Y(n_1460)
);

AOI21xp33_ASAP7_75t_L g1461 ( 
.A1(n_1392),
.A2(n_1384),
.B(n_1299),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1410),
.A2(n_1377),
.B1(n_1260),
.B2(n_1300),
.Y(n_1462)
);

AOI21xp33_ASAP7_75t_L g1463 ( 
.A1(n_1313),
.A2(n_1331),
.B(n_1277),
.Y(n_1463)
);

CKINVDCx20_ASAP7_75t_R g1464 ( 
.A(n_1276),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_SL g1465 ( 
.A1(n_1410),
.A2(n_1251),
.B1(n_1298),
.B2(n_1304),
.Y(n_1465)
);

BUFx12f_ASAP7_75t_L g1466 ( 
.A(n_1388),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1265),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1282),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1410),
.A2(n_1251),
.B1(n_1298),
.B2(n_1337),
.Y(n_1469)
);

BUFx12f_ASAP7_75t_L g1470 ( 
.A(n_1391),
.Y(n_1470)
);

OAI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1351),
.A2(n_1333),
.B1(n_1320),
.B2(n_1377),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1251),
.A2(n_1402),
.B1(n_1325),
.B2(n_1358),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1391),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1251),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1251),
.Y(n_1475)
);

CKINVDCx6p67_ASAP7_75t_R g1476 ( 
.A(n_1267),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1287),
.A2(n_1362),
.B1(n_1329),
.B2(n_1389),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1383),
.A2(n_1334),
.B1(n_1255),
.B2(n_1264),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1307),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1314),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1339),
.A2(n_1278),
.B1(n_1302),
.B2(n_1294),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1294),
.A2(n_1347),
.B1(n_1380),
.B2(n_1386),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1327),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1343),
.B(n_1347),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1314),
.Y(n_1485)
);

CKINVDCx11_ASAP7_75t_R g1486 ( 
.A(n_1314),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1294),
.A2(n_1381),
.B1(n_1367),
.B2(n_1369),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1284),
.A2(n_1352),
.B1(n_1330),
.B2(n_1318),
.Y(n_1488)
);

INVx4_ASAP7_75t_L g1489 ( 
.A(n_1254),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1343),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1354),
.Y(n_1491)
);

INVxp67_ASAP7_75t_SL g1492 ( 
.A(n_1326),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1273),
.A2(n_1336),
.B1(n_1262),
.B2(n_1343),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1340),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1297),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1346),
.B(n_1275),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1312),
.A2(n_1254),
.B1(n_1373),
.B2(n_1293),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1297),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1297),
.Y(n_1499)
);

OAI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1272),
.A2(n_1399),
.B1(n_1359),
.B2(n_1365),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1328),
.A2(n_1399),
.B1(n_1359),
.B2(n_1365),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1359),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1373),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1289),
.A2(n_1399),
.B1(n_1365),
.B2(n_1360),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1338),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1360),
.Y(n_1506)
);

BUFx4f_ASAP7_75t_SL g1507 ( 
.A(n_1274),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1360),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1269),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1279),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1271),
.A2(n_1268),
.B1(n_1315),
.B2(n_1387),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1395),
.A2(n_1085),
.B1(n_1181),
.B2(n_922),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1271),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_SL g1514 ( 
.A1(n_1301),
.A2(n_922),
.B1(n_1179),
.B2(n_1280),
.Y(n_1514)
);

CKINVDCx11_ASAP7_75t_R g1515 ( 
.A(n_1407),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1412),
.A2(n_1085),
.B1(n_1181),
.B2(n_922),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1412),
.A2(n_1085),
.B1(n_1181),
.B2(n_922),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1412),
.A2(n_1085),
.B1(n_1181),
.B2(n_922),
.Y(n_1518)
);

BUFx12f_ASAP7_75t_L g1519 ( 
.A(n_1270),
.Y(n_1519)
);

OAI21xp33_ASAP7_75t_L g1520 ( 
.A1(n_1364),
.A2(n_1403),
.B(n_1379),
.Y(n_1520)
);

BUFx4f_ASAP7_75t_L g1521 ( 
.A(n_1276),
.Y(n_1521)
);

BUFx12f_ASAP7_75t_L g1522 ( 
.A(n_1270),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1412),
.A2(n_1085),
.B1(n_1181),
.B2(n_922),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1374),
.B(n_1376),
.Y(n_1524)
);

AOI22x1_ASAP7_75t_SL g1525 ( 
.A1(n_1280),
.A2(n_1258),
.B1(n_277),
.B2(n_337),
.Y(n_1525)
);

INVx4_ASAP7_75t_L g1526 ( 
.A(n_1276),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1412),
.A2(n_922),
.B1(n_782),
.B2(n_1371),
.Y(n_1527)
);

BUFx2_ASAP7_75t_SL g1528 ( 
.A(n_1270),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1412),
.A2(n_922),
.B1(n_782),
.B2(n_1371),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1344),
.Y(n_1530)
);

INVx6_ASAP7_75t_L g1531 ( 
.A(n_1401),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1296),
.Y(n_1532)
);

CKINVDCx11_ASAP7_75t_R g1533 ( 
.A(n_1407),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1412),
.A2(n_1085),
.B1(n_1181),
.B2(n_922),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1412),
.A2(n_922),
.B1(n_782),
.B2(n_1371),
.Y(n_1535)
);

BUFx12f_ASAP7_75t_L g1536 ( 
.A(n_1270),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_1257),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1412),
.A2(n_1085),
.B1(n_1181),
.B2(n_922),
.Y(n_1538)
);

BUFx8_ASAP7_75t_L g1539 ( 
.A(n_1344),
.Y(n_1539)
);

INVx6_ASAP7_75t_L g1540 ( 
.A(n_1401),
.Y(n_1540)
);

CKINVDCx6p67_ASAP7_75t_R g1541 ( 
.A(n_1407),
.Y(n_1541)
);

CKINVDCx11_ASAP7_75t_R g1542 ( 
.A(n_1407),
.Y(n_1542)
);

CKINVDCx16_ASAP7_75t_R g1543 ( 
.A(n_1407),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1412),
.A2(n_1085),
.B1(n_1181),
.B2(n_922),
.Y(n_1544)
);

CKINVDCx11_ASAP7_75t_R g1545 ( 
.A(n_1407),
.Y(n_1545)
);

BUFx2_ASAP7_75t_SL g1546 ( 
.A(n_1270),
.Y(n_1546)
);

INVx4_ASAP7_75t_SL g1547 ( 
.A(n_1410),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1296),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1374),
.B(n_1376),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1412),
.A2(n_1085),
.B1(n_1181),
.B2(n_922),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1412),
.A2(n_1371),
.B1(n_1375),
.B2(n_1285),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1412),
.A2(n_1371),
.B1(n_1375),
.B2(n_1285),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1296),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1405),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1412),
.A2(n_1085),
.B1(n_1181),
.B2(n_922),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1412),
.A2(n_1371),
.B1(n_1375),
.B2(n_1285),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1405),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1296),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1296),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1448),
.A2(n_1511),
.B(n_1497),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1441),
.Y(n_1561)
);

OAI21x1_ASAP7_75t_L g1562 ( 
.A1(n_1497),
.A2(n_1487),
.B(n_1488),
.Y(n_1562)
);

INVxp33_ASAP7_75t_L g1563 ( 
.A(n_1438),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1558),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1441),
.B(n_1449),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1491),
.B(n_1484),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1491),
.B(n_1494),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1450),
.B(n_1506),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1494),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1442),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1479),
.A2(n_1482),
.B(n_1478),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1446),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1447),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1455),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1432),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1425),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1457),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1432),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1433),
.Y(n_1579)
);

INVxp67_ASAP7_75t_R g1580 ( 
.A(n_1496),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1433),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1490),
.Y(n_1582)
);

AO21x2_ASAP7_75t_L g1583 ( 
.A1(n_1495),
.A2(n_1499),
.B(n_1498),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1418),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1508),
.B(n_1502),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1451),
.Y(n_1586)
);

OA21x2_ASAP7_75t_L g1587 ( 
.A1(n_1504),
.A2(n_1478),
.B(n_1482),
.Y(n_1587)
);

OA21x2_ASAP7_75t_L g1588 ( 
.A1(n_1504),
.A2(n_1481),
.B(n_1458),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1429),
.Y(n_1589)
);

AND2x6_ASAP7_75t_L g1590 ( 
.A(n_1474),
.B(n_1475),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1431),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1524),
.B(n_1549),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1415),
.Y(n_1593)
);

INVx4_ASAP7_75t_R g1594 ( 
.A(n_1530),
.Y(n_1594)
);

AO21x2_ASAP7_75t_L g1595 ( 
.A1(n_1500),
.A2(n_1493),
.B(n_1439),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1424),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_SL g1597 ( 
.A(n_1426),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1483),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1513),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1503),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1513),
.Y(n_1601)
);

OAI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1527),
.A2(n_1535),
.B1(n_1529),
.B2(n_1552),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1516),
.A2(n_1555),
.B1(n_1550),
.B2(n_1518),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1474),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1458),
.A2(n_1472),
.B(n_1451),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1467),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1475),
.B(n_1547),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1468),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1501),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1516),
.A2(n_1555),
.B1(n_1544),
.B2(n_1523),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1547),
.B(n_1505),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1489),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1489),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1428),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_SL g1615 ( 
.A1(n_1551),
.A2(n_1556),
.B1(n_1514),
.B2(n_1525),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1532),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1548),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1553),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1559),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1456),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1456),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1507),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1452),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1510),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1510),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1471),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1416),
.B(n_1417),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1459),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1509),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1530),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1509),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1440),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1485),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1547),
.B(n_1492),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1416),
.B(n_1417),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1427),
.B(n_1434),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1445),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1420),
.B(n_1422),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1520),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1476),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1422),
.A2(n_1512),
.B(n_1434),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1445),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1421),
.Y(n_1643)
);

AO21x2_ASAP7_75t_L g1644 ( 
.A1(n_1463),
.A2(n_1461),
.B(n_1454),
.Y(n_1644)
);

AOI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1414),
.A2(n_1465),
.B(n_1435),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1427),
.B(n_1419),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1480),
.B(n_1518),
.Y(n_1647)
);

BUFx12f_ASAP7_75t_L g1648 ( 
.A(n_1515),
.Y(n_1648)
);

AO21x2_ASAP7_75t_L g1649 ( 
.A1(n_1462),
.A2(n_1512),
.B(n_1544),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1517),
.A2(n_1538),
.B1(n_1534),
.B2(n_1523),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1477),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1477),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1469),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1543),
.A2(n_1437),
.B1(n_1541),
.B2(n_1550),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1517),
.B(n_1538),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1534),
.B(n_1430),
.Y(n_1656)
);

OA21x2_ASAP7_75t_L g1657 ( 
.A1(n_1473),
.A2(n_1540),
.B(n_1531),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1540),
.A2(n_1486),
.B(n_1426),
.Y(n_1658)
);

AOI222xp33_ASAP7_75t_L g1659 ( 
.A1(n_1515),
.A2(n_1545),
.B1(n_1533),
.B2(n_1542),
.C1(n_1521),
.C2(n_1539),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1426),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1539),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1430),
.B(n_1546),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1539),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1528),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1545),
.B(n_1423),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1466),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1466),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1470),
.Y(n_1668)
);

BUFx3_ASAP7_75t_L g1669 ( 
.A(n_1470),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1519),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1638),
.A2(n_1443),
.B1(n_1537),
.B2(n_1526),
.C(n_1464),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1578),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1579),
.B(n_1557),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1566),
.B(n_1526),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1593),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1584),
.B(n_1460),
.Y(n_1676)
);

OA21x2_ASAP7_75t_L g1677 ( 
.A1(n_1560),
.A2(n_1413),
.B(n_1554),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1615),
.A2(n_1521),
.B1(n_1536),
.B2(n_1519),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_SL g1679 ( 
.A1(n_1638),
.A2(n_1522),
.B1(n_1536),
.B2(n_1460),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1584),
.B(n_1444),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1627),
.A2(n_1522),
.B1(n_1453),
.B2(n_1436),
.Y(n_1681)
);

O2A1O1Ixp33_ASAP7_75t_SL g1682 ( 
.A1(n_1602),
.A2(n_1614),
.B(n_1622),
.C(n_1654),
.Y(n_1682)
);

OA21x2_ASAP7_75t_L g1683 ( 
.A1(n_1560),
.A2(n_1562),
.B(n_1605),
.Y(n_1683)
);

AND2x6_ASAP7_75t_L g1684 ( 
.A(n_1611),
.B(n_1634),
.Y(n_1684)
);

AO21x2_ASAP7_75t_L g1685 ( 
.A1(n_1605),
.A2(n_1586),
.B(n_1626),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1589),
.B(n_1591),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1603),
.A2(n_1650),
.B1(n_1610),
.B2(n_1614),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1594),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1589),
.B(n_1591),
.Y(n_1689)
);

OR2x6_ASAP7_75t_L g1690 ( 
.A(n_1611),
.B(n_1657),
.Y(n_1690)
);

AND2x2_ASAP7_75t_SL g1691 ( 
.A(n_1627),
.B(n_1635),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1576),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1566),
.B(n_1611),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1564),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1561),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1595),
.A2(n_1644),
.B(n_1655),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1570),
.Y(n_1697)
);

NAND4xp25_ASAP7_75t_L g1698 ( 
.A(n_1639),
.B(n_1664),
.C(n_1622),
.D(n_1659),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1566),
.B(n_1611),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1635),
.A2(n_1626),
.B(n_1562),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1657),
.A2(n_1634),
.B(n_1595),
.Y(n_1701)
);

NOR2x1_ASAP7_75t_SL g1702 ( 
.A(n_1629),
.B(n_1631),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1595),
.A2(n_1644),
.B(n_1587),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_SL g1704 ( 
.A1(n_1656),
.A2(n_1629),
.B(n_1631),
.C(n_1664),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1561),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1580),
.B(n_1575),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1641),
.A2(n_1628),
.B(n_1645),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1644),
.B(n_1630),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1620),
.A2(n_1621),
.B1(n_1628),
.B2(n_1653),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1580),
.B(n_1575),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1641),
.A2(n_1620),
.B(n_1621),
.C(n_1636),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1581),
.B(n_1563),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1572),
.B(n_1573),
.Y(n_1713)
);

A2O1A1Ixp33_ASAP7_75t_L g1714 ( 
.A1(n_1636),
.A2(n_1653),
.B(n_1643),
.C(n_1647),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1645),
.A2(n_1609),
.B(n_1571),
.Y(n_1715)
);

OAI211xp5_ASAP7_75t_L g1716 ( 
.A1(n_1609),
.A2(n_1643),
.B(n_1633),
.C(n_1587),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1623),
.B(n_1592),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1565),
.B(n_1616),
.Y(n_1718)
);

OAI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1646),
.A2(n_1588),
.B1(n_1587),
.B2(n_1637),
.C(n_1642),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1574),
.Y(n_1720)
);

OAI21x1_ASAP7_75t_SL g1721 ( 
.A1(n_1668),
.A2(n_1661),
.B(n_1660),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1587),
.B(n_1604),
.Y(n_1722)
);

OAI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1588),
.A2(n_1596),
.B(n_1613),
.C(n_1612),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1617),
.B(n_1619),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1604),
.B(n_1588),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1597),
.A2(n_1663),
.B1(n_1660),
.B2(n_1661),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1663),
.B(n_1665),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1617),
.Y(n_1728)
);

AO21x2_ASAP7_75t_L g1729 ( 
.A1(n_1583),
.A2(n_1598),
.B(n_1599),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1658),
.Y(n_1730)
);

A2O1A1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1658),
.A2(n_1619),
.B(n_1652),
.C(n_1651),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1568),
.B(n_1618),
.Y(n_1732)
);

NOR3xp33_ASAP7_75t_L g1733 ( 
.A(n_1632),
.B(n_1640),
.C(n_1624),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_SL g1734 ( 
.A1(n_1648),
.A2(n_1669),
.B1(n_1670),
.B2(n_1666),
.Y(n_1734)
);

OR2x6_ASAP7_75t_L g1735 ( 
.A(n_1657),
.B(n_1567),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1725),
.Y(n_1736)
);

INVxp67_ASAP7_75t_SL g1737 ( 
.A(n_1708),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1675),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1720),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1695),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1687),
.A2(n_1648),
.B1(n_1625),
.B2(n_1624),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1695),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1691),
.A2(n_1625),
.B1(n_1670),
.B2(n_1666),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1672),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1705),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1691),
.A2(n_1709),
.B1(n_1678),
.B2(n_1714),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1700),
.A2(n_1649),
.B1(n_1642),
.B2(n_1601),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1707),
.A2(n_1649),
.B1(n_1696),
.B2(n_1719),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1722),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1722),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1692),
.B(n_1694),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_SL g1752 ( 
.A1(n_1731),
.A2(n_1657),
.B(n_1607),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1721),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1693),
.B(n_1699),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1685),
.A2(n_1649),
.B1(n_1601),
.B2(n_1599),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_SL g1756 ( 
.A1(n_1716),
.A2(n_1607),
.B1(n_1590),
.B2(n_1569),
.Y(n_1756)
);

NOR2xp67_ASAP7_75t_L g1757 ( 
.A(n_1723),
.B(n_1600),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1718),
.B(n_1585),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1693),
.B(n_1590),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1699),
.B(n_1590),
.Y(n_1760)
);

INVx4_ASAP7_75t_L g1761 ( 
.A(n_1684),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1697),
.Y(n_1762)
);

NOR2x1_ASAP7_75t_L g1763 ( 
.A(n_1701),
.B(n_1730),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1685),
.A2(n_1606),
.B1(n_1608),
.B2(n_1577),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1717),
.B(n_1582),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1713),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1740),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1746),
.A2(n_1714),
.B1(n_1711),
.B2(n_1681),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1739),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1765),
.B(n_1686),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1754),
.B(n_1676),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1758),
.B(n_1724),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1740),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1742),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1761),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1753),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1746),
.A2(n_1703),
.B1(n_1715),
.B2(n_1698),
.Y(n_1777)
);

AND2x2_ASAP7_75t_SL g1778 ( 
.A(n_1761),
.B(n_1677),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1744),
.B(n_1666),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1742),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1754),
.B(n_1676),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1736),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1761),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1752),
.A2(n_1682),
.B(n_1704),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1736),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1736),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1743),
.A2(n_1681),
.B1(n_1679),
.B2(n_1688),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1754),
.B(n_1712),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1761),
.Y(n_1789)
);

OAI31xp33_ASAP7_75t_L g1790 ( 
.A1(n_1741),
.A2(n_1682),
.A3(n_1743),
.B(n_1711),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1753),
.Y(n_1791)
);

INVx1_ASAP7_75t_SL g1792 ( 
.A(n_1753),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1741),
.A2(n_1688),
.B1(n_1731),
.B2(n_1671),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1754),
.B(n_1680),
.Y(n_1794)
);

OAI33xp33_ASAP7_75t_L g1795 ( 
.A1(n_1751),
.A2(n_1726),
.A3(n_1734),
.B1(n_1728),
.B2(n_1732),
.B3(n_1667),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1758),
.B(n_1686),
.Y(n_1796)
);

INVx3_ASAP7_75t_L g1797 ( 
.A(n_1759),
.Y(n_1797)
);

INVxp67_ASAP7_75t_SL g1798 ( 
.A(n_1757),
.Y(n_1798)
);

AO21x2_ASAP7_75t_L g1799 ( 
.A1(n_1757),
.A2(n_1729),
.B(n_1752),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1759),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_L g1801 ( 
.A(n_1748),
.B(n_1683),
.C(n_1677),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1745),
.Y(n_1802)
);

AOI21xp33_ASAP7_75t_L g1803 ( 
.A1(n_1763),
.A2(n_1677),
.B(n_1683),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1749),
.B(n_1750),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1737),
.A2(n_1704),
.B(n_1702),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1747),
.A2(n_1690),
.B1(n_1683),
.B2(n_1735),
.Y(n_1806)
);

NAND4xp25_ASAP7_75t_L g1807 ( 
.A(n_1751),
.B(n_1680),
.C(n_1673),
.D(n_1727),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1750),
.B(n_1689),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1756),
.A2(n_1674),
.B1(n_1706),
.B2(n_1710),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1739),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1767),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1800),
.B(n_1797),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1767),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1796),
.B(n_1750),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1799),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1797),
.B(n_1771),
.Y(n_1816)
);

INVx2_ASAP7_75t_SL g1817 ( 
.A(n_1791),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1773),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_R g1819 ( 
.A(n_1779),
.B(n_1666),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1799),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1807),
.B(n_1670),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1799),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1769),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1773),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1771),
.B(n_1759),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1781),
.B(n_1760),
.Y(n_1826)
);

BUFx2_ASAP7_75t_L g1827 ( 
.A(n_1791),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1810),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1796),
.B(n_1766),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1770),
.B(n_1762),
.Y(n_1830)
);

NAND4xp25_ASAP7_75t_L g1831 ( 
.A(n_1790),
.B(n_1662),
.C(n_1665),
.D(n_1669),
.Y(n_1831)
);

OAI21x1_ASAP7_75t_L g1832 ( 
.A1(n_1805),
.A2(n_1755),
.B(n_1764),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1799),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1795),
.B(n_1738),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1774),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1774),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1772),
.B(n_1808),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1780),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1772),
.B(n_1766),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1780),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1782),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1781),
.B(n_1760),
.Y(n_1842)
);

CKINVDCx16_ASAP7_75t_R g1843 ( 
.A(n_1768),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1808),
.B(n_1765),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1794),
.B(n_1760),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1791),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1837),
.B(n_1804),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1834),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1811),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1811),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1843),
.B(n_1802),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1837),
.B(n_1844),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1825),
.B(n_1794),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1813),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1825),
.B(n_1775),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1813),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1843),
.B(n_1782),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1834),
.B(n_1785),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1818),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1831),
.A2(n_1768),
.B1(n_1777),
.B2(n_1790),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1827),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1828),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_1827),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1815),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1826),
.B(n_1775),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1815),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1815),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1818),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1820),
.Y(n_1869)
);

INVx2_ASAP7_75t_SL g1870 ( 
.A(n_1812),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1826),
.B(n_1783),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1842),
.B(n_1783),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1824),
.Y(n_1873)
);

INVxp67_ASAP7_75t_SL g1874 ( 
.A(n_1828),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1820),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1844),
.B(n_1804),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1839),
.B(n_1785),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1842),
.B(n_1789),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1823),
.B(n_1785),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1824),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1823),
.B(n_1786),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1835),
.Y(n_1882)
);

INVxp67_ASAP7_75t_SL g1883 ( 
.A(n_1846),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1839),
.B(n_1830),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1845),
.B(n_1789),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1835),
.B(n_1786),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1830),
.B(n_1786),
.Y(n_1887)
);

INVxp67_ASAP7_75t_L g1888 ( 
.A(n_1821),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1836),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1845),
.B(n_1788),
.Y(n_1890)
);

INVxp67_ASAP7_75t_SL g1891 ( 
.A(n_1846),
.Y(n_1891)
);

BUFx2_ASAP7_75t_L g1892 ( 
.A(n_1817),
.Y(n_1892)
);

OAI21xp33_ASAP7_75t_L g1893 ( 
.A1(n_1860),
.A2(n_1848),
.B(n_1831),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1874),
.B(n_1836),
.Y(n_1894)
);

OR2x6_ASAP7_75t_L g1895 ( 
.A(n_1857),
.B(n_1784),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1862),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1849),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1870),
.B(n_1819),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1849),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1883),
.B(n_1817),
.Y(n_1900)
);

AOI211xp5_ASAP7_75t_L g1901 ( 
.A1(n_1851),
.A2(n_1787),
.B(n_1793),
.C(n_1801),
.Y(n_1901)
);

INVx1_ASAP7_75t_SL g1902 ( 
.A(n_1851),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1852),
.B(n_1838),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1850),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1850),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1852),
.B(n_1829),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1854),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1858),
.B(n_1829),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1888),
.B(n_1807),
.Y(n_1909)
);

INVxp67_ASAP7_75t_SL g1910 ( 
.A(n_1891),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1858),
.B(n_1838),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1861),
.B(n_1863),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1861),
.B(n_1863),
.Y(n_1913)
);

NOR3xp33_ASAP7_75t_L g1914 ( 
.A(n_1892),
.B(n_1801),
.C(n_1817),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1884),
.B(n_1847),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1854),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1884),
.B(n_1814),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1853),
.B(n_1816),
.Y(n_1918)
);

NAND3xp33_ASAP7_75t_L g1919 ( 
.A(n_1892),
.B(n_1803),
.C(n_1820),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1890),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1847),
.B(n_1814),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1890),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1856),
.B(n_1840),
.Y(n_1923)
);

INVx2_ASAP7_75t_SL g1924 ( 
.A(n_1855),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1856),
.B(n_1840),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1853),
.B(n_1816),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1859),
.Y(n_1927)
);

AOI21xp33_ASAP7_75t_L g1928 ( 
.A1(n_1857),
.A2(n_1833),
.B(n_1822),
.Y(n_1928)
);

INVx2_ASAP7_75t_SL g1929 ( 
.A(n_1855),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1897),
.Y(n_1930)
);

OAI32xp33_ASAP7_75t_L g1931 ( 
.A1(n_1893),
.A2(n_1870),
.A3(n_1792),
.B1(n_1776),
.B2(n_1879),
.Y(n_1931)
);

XNOR2x1_ASAP7_75t_L g1932 ( 
.A(n_1895),
.B(n_1832),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1910),
.B(n_1776),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1899),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1901),
.A2(n_1798),
.B1(n_1832),
.B2(n_1806),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1918),
.Y(n_1936)
);

O2A1O1Ixp33_ASAP7_75t_L g1937 ( 
.A1(n_1912),
.A2(n_1822),
.B(n_1833),
.C(n_1881),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1902),
.B(n_1896),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1924),
.B(n_1792),
.Y(n_1939)
);

AOI322xp5_ASAP7_75t_L g1940 ( 
.A1(n_1909),
.A2(n_1822),
.A3(n_1833),
.B1(n_1879),
.B2(n_1881),
.C1(n_1864),
.C2(n_1875),
.Y(n_1940)
);

CKINVDCx16_ASAP7_75t_R g1941 ( 
.A(n_1895),
.Y(n_1941)
);

AOI21xp33_ASAP7_75t_SL g1942 ( 
.A1(n_1895),
.A2(n_1929),
.B(n_1914),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1900),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1920),
.B(n_1865),
.Y(n_1944)
);

AOI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1911),
.A2(n_1832),
.B1(n_1778),
.B2(n_1809),
.Y(n_1945)
);

OAI211xp5_ASAP7_75t_L g1946 ( 
.A1(n_1913),
.A2(n_1865),
.B(n_1871),
.C(n_1885),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1913),
.B(n_1871),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1904),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1905),
.Y(n_1949)
);

INVxp33_ASAP7_75t_L g1950 ( 
.A(n_1900),
.Y(n_1950)
);

AOI21xp33_ASAP7_75t_L g1951 ( 
.A1(n_1911),
.A2(n_1868),
.B(n_1859),
.Y(n_1951)
);

NAND2xp33_ASAP7_75t_L g1952 ( 
.A(n_1915),
.B(n_1872),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1922),
.Y(n_1953)
);

OAI22xp5_ASAP7_75t_SL g1954 ( 
.A1(n_1894),
.A2(n_1669),
.B1(n_1670),
.B2(n_1919),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1908),
.A2(n_1778),
.B1(n_1756),
.B2(n_1841),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1907),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1943),
.Y(n_1957)
);

OAI221xp5_ASAP7_75t_L g1958 ( 
.A1(n_1932),
.A2(n_1928),
.B1(n_1903),
.B2(n_1921),
.C(n_1894),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1930),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1947),
.B(n_1906),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1934),
.Y(n_1961)
);

OAI21xp33_ASAP7_75t_L g1962 ( 
.A1(n_1945),
.A2(n_1903),
.B(n_1917),
.Y(n_1962)
);

NAND3xp33_ASAP7_75t_L g1963 ( 
.A(n_1940),
.B(n_1928),
.C(n_1927),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1948),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1935),
.A2(n_1916),
.B1(n_1875),
.B2(n_1867),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1949),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1956),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1947),
.B(n_1926),
.Y(n_1968)
);

INVx1_ASAP7_75t_SL g1969 ( 
.A(n_1941),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1943),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1953),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1936),
.B(n_1872),
.Y(n_1972)
);

INVx1_ASAP7_75t_SL g1973 ( 
.A(n_1952),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1953),
.Y(n_1974)
);

NOR3xp33_ASAP7_75t_L g1975 ( 
.A(n_1942),
.B(n_1925),
.C(n_1923),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1938),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1944),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1969),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1957),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1973),
.B(n_1950),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1957),
.Y(n_1981)
);

NOR3x1_ASAP7_75t_L g1982 ( 
.A(n_1958),
.B(n_1960),
.C(n_1968),
.Y(n_1982)
);

INVxp67_ASAP7_75t_L g1983 ( 
.A(n_1970),
.Y(n_1983)
);

OAI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1965),
.A2(n_1950),
.B1(n_1955),
.B2(n_1933),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1977),
.B(n_1933),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1963),
.B(n_1951),
.Y(n_1986)
);

OAI31xp33_ASAP7_75t_L g1987 ( 
.A1(n_1965),
.A2(n_1954),
.A3(n_1937),
.B(n_1946),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1970),
.Y(n_1988)
);

OAI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1975),
.A2(n_1931),
.B(n_1939),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1971),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1987),
.A2(n_1962),
.B(n_1977),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1978),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1978),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1985),
.B(n_1974),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1985),
.Y(n_1995)
);

INVx2_ASAP7_75t_SL g1996 ( 
.A(n_1980),
.Y(n_1996)
);

NOR3xp33_ASAP7_75t_L g1997 ( 
.A(n_1980),
.B(n_1976),
.C(n_1966),
.Y(n_1997)
);

AOI211xp5_ASAP7_75t_L g1998 ( 
.A1(n_1986),
.A2(n_1989),
.B(n_1984),
.C(n_1990),
.Y(n_1998)
);

OAI211xp5_ASAP7_75t_L g1999 ( 
.A1(n_1986),
.A2(n_1961),
.B(n_1959),
.C(n_1964),
.Y(n_1999)
);

INVx2_ASAP7_75t_SL g2000 ( 
.A(n_1990),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1979),
.Y(n_2001)
);

NAND3xp33_ASAP7_75t_L g2002 ( 
.A(n_1983),
.B(n_1967),
.C(n_1961),
.Y(n_2002)
);

AOI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1998),
.A2(n_1988),
.B1(n_1981),
.B2(n_1939),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1992),
.Y(n_2004)
);

AOI211xp5_ASAP7_75t_L g2005 ( 
.A1(n_1998),
.A2(n_1959),
.B(n_1982),
.C(n_1972),
.Y(n_2005)
);

OAI211xp5_ASAP7_75t_SL g2006 ( 
.A1(n_1991),
.A2(n_1898),
.B(n_1667),
.C(n_1668),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1996),
.B(n_1923),
.Y(n_2007)
);

NAND3xp33_ASAP7_75t_L g2008 ( 
.A(n_1999),
.B(n_1925),
.C(n_1873),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1995),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_2004),
.B(n_1993),
.Y(n_2010)
);

NOR2x1_ASAP7_75t_L g2011 ( 
.A(n_2009),
.B(n_2002),
.Y(n_2011)
);

OAI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_2003),
.A2(n_1994),
.B1(n_2001),
.B2(n_2000),
.Y(n_2012)
);

AOI221xp5_ASAP7_75t_L g2013 ( 
.A1(n_2005),
.A2(n_1997),
.B1(n_1869),
.B2(n_1866),
.C(n_1875),
.Y(n_2013)
);

NAND3xp33_ASAP7_75t_L g2014 ( 
.A(n_2007),
.B(n_1873),
.C(n_1868),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_2008),
.Y(n_2015)
);

AOI221xp5_ASAP7_75t_L g2016 ( 
.A1(n_2006),
.A2(n_1869),
.B1(n_1864),
.B2(n_1866),
.C(n_1867),
.Y(n_2016)
);

OAI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_2011),
.A2(n_1889),
.B1(n_1880),
.B2(n_1882),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_2010),
.Y(n_2018)
);

INVx3_ASAP7_75t_L g2019 ( 
.A(n_2015),
.Y(n_2019)
);

NOR2x1_ASAP7_75t_L g2020 ( 
.A(n_2012),
.B(n_1662),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_2013),
.B(n_2014),
.Y(n_2021)
);

INVx1_ASAP7_75t_SL g2022 ( 
.A(n_2016),
.Y(n_2022)
);

BUFx2_ASAP7_75t_L g2023 ( 
.A(n_2020),
.Y(n_2023)
);

OAI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_2018),
.A2(n_1889),
.B1(n_1880),
.B2(n_1882),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_2019),
.B(n_1876),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_2023),
.B(n_2025),
.Y(n_2026)
);

OAI22x1_ASAP7_75t_L g2027 ( 
.A1(n_2026),
.A2(n_2022),
.B1(n_2021),
.B2(n_2017),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2027),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_2027),
.Y(n_2029)
);

CKINVDCx20_ASAP7_75t_R g2030 ( 
.A(n_2028),
.Y(n_2030)
);

OAI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_2029),
.A2(n_2024),
.B1(n_1887),
.B2(n_1866),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_2030),
.A2(n_1867),
.B(n_1869),
.Y(n_2032)
);

OAI21xp5_ASAP7_75t_SL g2033 ( 
.A1(n_2031),
.A2(n_1864),
.B(n_1640),
.Y(n_2033)
);

AOI22xp33_ASAP7_75t_SL g2034 ( 
.A1(n_2032),
.A2(n_1778),
.B1(n_1886),
.B2(n_1887),
.Y(n_2034)
);

AO21x2_ASAP7_75t_L g2035 ( 
.A1(n_2034),
.A2(n_2033),
.B(n_1886),
.Y(n_2035)
);

HB1xp67_ASAP7_75t_L g2036 ( 
.A(n_2035),
.Y(n_2036)
);

OAI221xp5_ASAP7_75t_R g2037 ( 
.A1(n_2036),
.A2(n_1885),
.B1(n_1878),
.B2(n_1812),
.C(n_1733),
.Y(n_2037)
);

OAI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_2037),
.A2(n_1876),
.B1(n_1877),
.B2(n_1878),
.Y(n_2038)
);


endmodule