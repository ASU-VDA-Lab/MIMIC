module real_aes_2319_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_0), .B(n_511), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_1), .A2(n_514), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_2), .B(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_3), .B(n_217), .Y(n_517) );
INVx1_ASAP7_75t_L g149 ( .A(n_4), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_5), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_6), .B(n_217), .Y(n_587) );
INVx1_ASAP7_75t_L g181 ( .A(n_7), .Y(n_181) );
CKINVDCx16_ASAP7_75t_R g832 ( .A(n_8), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_9), .Y(n_196) );
NAND2xp33_ASAP7_75t_L g572 ( .A(n_10), .B(n_214), .Y(n_572) );
INVx2_ASAP7_75t_L g141 ( .A(n_11), .Y(n_141) );
AOI221x1_ASAP7_75t_L g521 ( .A1(n_12), .A2(n_24), .B1(n_511), .B2(n_514), .C(n_522), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_13), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_14), .B(n_511), .Y(n_568) );
INVx1_ASAP7_75t_L g215 ( .A(n_15), .Y(n_215) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_16), .A2(n_178), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_17), .B(n_172), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_18), .B(n_217), .Y(n_561) );
AO21x1_ASAP7_75t_L g510 ( .A1(n_19), .A2(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g116 ( .A(n_20), .Y(n_116) );
INVx1_ASAP7_75t_L g212 ( .A(n_21), .Y(n_212) );
INVx1_ASAP7_75t_SL g266 ( .A(n_22), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_23), .B(n_164), .Y(n_228) );
AOI33xp33_ASAP7_75t_L g252 ( .A1(n_25), .A2(n_54), .A3(n_146), .B1(n_157), .B2(n_253), .B3(n_254), .Y(n_252) );
NAND2x1_ASAP7_75t_L g532 ( .A(n_26), .B(n_217), .Y(n_532) );
NAND2x1_ASAP7_75t_L g586 ( .A(n_27), .B(n_214), .Y(n_586) );
INVx1_ASAP7_75t_L g189 ( .A(n_28), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_29), .Y(n_118) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_30), .A2(n_87), .B(n_141), .Y(n_140) );
OR2x2_ASAP7_75t_L g174 ( .A(n_30), .B(n_87), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g834 ( .A(n_31), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_32), .B(n_144), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_33), .B(n_214), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_34), .B(n_217), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_35), .A2(n_64), .B1(n_819), .B2(n_820), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_35), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_36), .B(n_214), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_37), .A2(n_514), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g151 ( .A(n_38), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g156 ( .A(n_38), .Y(n_156) );
AND2x2_ASAP7_75t_L g170 ( .A(n_38), .B(n_149), .Y(n_170) );
OR2x6_ASAP7_75t_L g114 ( .A(n_39), .B(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_40), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_41), .B(n_511), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_42), .B(n_144), .Y(n_143) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_43), .A2(n_139), .B1(n_206), .B2(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_44), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_45), .B(n_164), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_46), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_47), .A2(n_95), .B1(n_803), .B2(n_804), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_47), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_48), .B(n_214), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_49), .B(n_178), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_50), .B(n_164), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_51), .A2(n_514), .B(n_585), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_52), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_53), .B(n_214), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_55), .B(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g147 ( .A(n_56), .Y(n_147) );
INVx1_ASAP7_75t_L g166 ( .A(n_56), .Y(n_166) );
AND2x2_ASAP7_75t_L g171 ( .A(n_57), .B(n_172), .Y(n_171) );
AOI221xp5_ASAP7_75t_L g179 ( .A1(n_58), .A2(n_76), .B1(n_144), .B2(n_154), .C(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_59), .B(n_144), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_60), .B(n_217), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_61), .B(n_139), .Y(n_198) );
AOI21xp5_ASAP7_75t_SL g236 ( .A1(n_62), .A2(n_154), .B(n_237), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_63), .A2(n_514), .B(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_64), .Y(n_819) );
INVx1_ASAP7_75t_L g209 ( .A(n_65), .Y(n_209) );
AO21x1_ASAP7_75t_L g513 ( .A1(n_66), .A2(n_514), .B(n_515), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_67), .B(n_511), .Y(n_577) );
INVx1_ASAP7_75t_L g161 ( .A(n_68), .Y(n_161) );
AOI22xp33_ASAP7_75t_SL g805 ( .A1(n_69), .A2(n_802), .B1(n_806), .B2(n_810), .Y(n_805) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_70), .B(n_511), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_71), .A2(n_154), .B(n_160), .Y(n_153) );
AND2x2_ASAP7_75t_L g545 ( .A(n_72), .B(n_173), .Y(n_545) );
INVx1_ASAP7_75t_L g152 ( .A(n_73), .Y(n_152) );
INVx1_ASAP7_75t_L g168 ( .A(n_73), .Y(n_168) );
AND2x2_ASAP7_75t_L g589 ( .A(n_74), .B(n_138), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_75), .B(n_144), .Y(n_255) );
AND2x2_ASAP7_75t_L g268 ( .A(n_77), .B(n_138), .Y(n_268) );
INVx1_ASAP7_75t_L g210 ( .A(n_78), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_79), .A2(n_154), .B(n_265), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_80), .A2(n_154), .B(n_227), .C(n_231), .Y(n_226) );
INVx1_ASAP7_75t_L g117 ( .A(n_81), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_82), .B(n_511), .Y(n_563) );
AND2x2_ASAP7_75t_SL g234 ( .A(n_83), .B(n_138), .Y(n_234) );
AND2x2_ASAP7_75t_L g575 ( .A(n_84), .B(n_138), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_85), .A2(n_154), .B1(n_250), .B2(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_L g512 ( .A(n_86), .B(n_206), .Y(n_512) );
AND2x2_ASAP7_75t_L g535 ( .A(n_88), .B(n_138), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_89), .B(n_214), .Y(n_562) );
INVx1_ASAP7_75t_L g238 ( .A(n_90), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_91), .B(n_217), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_92), .B(n_214), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_93), .A2(n_514), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g256 ( .A(n_94), .B(n_138), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_95), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_96), .B(n_217), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_97), .A2(n_187), .B(n_188), .C(n_191), .Y(n_186) );
BUFx2_ASAP7_75t_L g106 ( .A(n_98), .Y(n_106) );
BUFx2_ASAP7_75t_SL g823 ( .A(n_98), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_99), .A2(n_514), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_100), .B(n_164), .Y(n_239) );
AOI21xp33_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_824), .B(n_833), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_119), .B(n_814), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
NAND3xp33_ASAP7_75t_L g814 ( .A(n_107), .B(n_815), .C(n_822), .Y(n_814) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_118), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g815 ( .A(n_108), .B(n_816), .Y(n_815) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g829 ( .A(n_111), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
OR2x6_ASAP7_75t_SL g125 ( .A(n_112), .B(n_113), .Y(n_125) );
AND2x6_ASAP7_75t_SL g501 ( .A(n_112), .B(n_114), .Y(n_501) );
OR2x2_ASAP7_75t_L g813 ( .A(n_112), .B(n_114), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
OAI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_802), .B(n_805), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_126), .B1(n_498), .B2(n_502), .Y(n_121) );
BUFx4f_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_124), .Y(n_809) );
CKINVDCx11_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_127), .A2(n_807), .B1(n_808), .B2(n_809), .Y(n_806) );
NAND4xp75_ASAP7_75t_L g127 ( .A(n_128), .B(n_370), .C(n_415), .D(n_484), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NAND2x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_330), .Y(n_129) );
NOR3xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_286), .C(n_311), .Y(n_130) );
OAI222xp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_200), .B1(n_241), .B2(n_257), .C1(n_273), .C2(n_280), .Y(n_131) );
INVxp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_175), .Y(n_133) );
AND2x2_ASAP7_75t_L g495 ( .A(n_134), .B(n_309), .Y(n_495) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_136), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_136), .B(n_184), .Y(n_285) );
INVx3_ASAP7_75t_L g300 ( .A(n_136), .Y(n_300) );
AND2x2_ASAP7_75t_L g433 ( .A(n_136), .B(n_434), .Y(n_433) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_142), .B(n_171), .Y(n_136) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_137), .A2(n_138), .B1(n_186), .B2(n_192), .Y(n_185) );
AO21x2_ASAP7_75t_L g318 ( .A1(n_137), .A2(n_142), .B(n_171), .Y(n_318) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_137), .A2(n_529), .B(n_535), .Y(n_528) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_137), .A2(n_539), .B(n_545), .Y(n_538) );
AO21x2_ASAP7_75t_L g550 ( .A1(n_137), .A2(n_529), .B(n_535), .Y(n_550) );
AO21x2_ASAP7_75t_L g552 ( .A1(n_137), .A2(n_539), .B(n_545), .Y(n_552) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx4_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_139), .B(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx4f_ASAP7_75t_L g178 ( .A(n_140), .Y(n_178) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_141), .B(n_174), .Y(n_173) );
AND2x4_ASAP7_75t_L g206 ( .A(n_141), .B(n_174), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_153), .Y(n_142) );
INVx1_ASAP7_75t_L g199 ( .A(n_144), .Y(n_199) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_150), .Y(n_144) );
INVx1_ASAP7_75t_L g223 ( .A(n_145), .Y(n_223) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
OR2x6_ASAP7_75t_L g162 ( .A(n_146), .B(n_158), .Y(n_162) );
INVxp33_ASAP7_75t_L g253 ( .A(n_146), .Y(n_253) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g159 ( .A(n_147), .B(n_149), .Y(n_159) );
AND2x4_ASAP7_75t_L g217 ( .A(n_147), .B(n_167), .Y(n_217) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g224 ( .A(n_150), .Y(n_224) );
BUFx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x6_ASAP7_75t_L g514 ( .A(n_151), .B(n_159), .Y(n_514) );
INVx2_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
AND2x6_ASAP7_75t_L g214 ( .A(n_152), .B(n_165), .Y(n_214) );
INVxp67_ASAP7_75t_L g197 ( .A(n_154), .Y(n_197) );
AND2x4_ASAP7_75t_L g154 ( .A(n_155), .B(n_159), .Y(n_154) );
NOR2x1p5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx1_ASAP7_75t_L g254 ( .A(n_157), .Y(n_254) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_163), .C(n_169), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_SL g180 ( .A1(n_162), .A2(n_169), .B(n_181), .C(n_182), .Y(n_180) );
INVxp67_ASAP7_75t_L g187 ( .A(n_162), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_162), .A2(n_190), .B1(n_209), .B2(n_210), .Y(n_208) );
INVx2_ASAP7_75t_L g230 ( .A(n_162), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_162), .A2(n_169), .B(n_238), .C(n_239), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_SL g265 ( .A1(n_162), .A2(n_169), .B(n_266), .C(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g190 ( .A(n_164), .Y(n_190) );
AND2x4_ASAP7_75t_L g511 ( .A(n_164), .B(n_170), .Y(n_511) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_167), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_169), .B(n_206), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_169), .A2(n_228), .B(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g250 ( .A(n_169), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_169), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_169), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_169), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_169), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_169), .A2(n_561), .B(n_562), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_169), .A2(n_571), .B(n_572), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_169), .A2(n_580), .B(n_581), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_169), .A2(n_586), .B(n_587), .Y(n_585) );
INVx5_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_170), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_172), .Y(n_261) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_172), .A2(n_521), .B(n_525), .Y(n_520) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_172), .A2(n_521), .B(n_525), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_172), .A2(n_577), .B(n_578), .Y(n_576) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g363 ( .A(n_175), .B(n_316), .Y(n_363) );
AND2x2_ASAP7_75t_L g365 ( .A(n_175), .B(n_366), .Y(n_365) );
INVx3_ASAP7_75t_L g400 ( .A(n_175), .Y(n_400) );
AND2x4_ASAP7_75t_L g175 ( .A(n_176), .B(n_184), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVxp67_ASAP7_75t_L g283 ( .A(n_177), .Y(n_283) );
INVx1_ASAP7_75t_L g302 ( .A(n_177), .Y(n_302) );
AND2x4_ASAP7_75t_L g309 ( .A(n_177), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_177), .B(n_247), .Y(n_325) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_177), .Y(n_434) );
INVx1_ASAP7_75t_L g444 ( .A(n_177), .Y(n_444) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_183), .Y(n_177) );
INVx2_ASAP7_75t_SL g231 ( .A(n_178), .Y(n_231) );
INVx1_ASAP7_75t_L g244 ( .A(n_184), .Y(n_244) );
INVx2_ASAP7_75t_L g297 ( .A(n_184), .Y(n_297) );
INVx1_ASAP7_75t_L g378 ( .A(n_184), .Y(n_378) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_193), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_197), .B1(n_198), .B2(n_199), .Y(n_193) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_202), .B(n_232), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_202), .B(n_259), .Y(n_353) );
INVx2_ASAP7_75t_L g374 ( .A(n_202), .Y(n_374) );
AND2x2_ASAP7_75t_L g382 ( .A(n_202), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_219), .Y(n_202) );
AND2x4_ASAP7_75t_L g272 ( .A(n_203), .B(n_220), .Y(n_272) );
INVx1_ASAP7_75t_L g279 ( .A(n_203), .Y(n_279) );
AND2x2_ASAP7_75t_L g455 ( .A(n_203), .B(n_260), .Y(n_455) );
INVx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g293 ( .A(n_204), .B(n_220), .Y(n_293) );
INVx2_ASAP7_75t_L g329 ( .A(n_204), .Y(n_329) );
AND2x2_ASAP7_75t_L g408 ( .A(n_204), .B(n_260), .Y(n_408) );
NOR2x1_ASAP7_75t_SL g451 ( .A(n_204), .B(n_233), .Y(n_451) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_207), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_206), .A2(n_236), .B(n_240), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_206), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_SL g557 ( .A(n_206), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_206), .A2(n_568), .B(n_569), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_211), .B(n_218), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B1(n_215), .B2(n_216), .Y(n_211) );
INVxp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVxp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g291 ( .A(n_219), .Y(n_291) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g305 ( .A(n_220), .B(n_233), .Y(n_305) );
INVx1_ASAP7_75t_L g321 ( .A(n_220), .Y(n_321) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_220), .Y(n_429) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_226), .Y(n_220) );
NOR3xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .C(n_225), .Y(n_222) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_231), .A2(n_248), .B(n_256), .Y(n_247) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_231), .A2(n_248), .B(n_256), .Y(n_298) );
AND2x2_ASAP7_75t_L g292 ( .A(n_232), .B(n_293), .Y(n_292) );
OR2x6_ASAP7_75t_L g373 ( .A(n_232), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g411 ( .A(n_232), .B(n_408), .Y(n_411) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx4_ASAP7_75t_L g270 ( .A(n_233), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_233), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g340 ( .A(n_233), .Y(n_340) );
OR2x2_ASAP7_75t_L g346 ( .A(n_233), .B(n_260), .Y(n_346) );
AND2x4_ASAP7_75t_L g360 ( .A(n_233), .B(n_321), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_233), .B(n_329), .Y(n_361) );
OR2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_245), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g405 ( .A(n_244), .B(n_324), .Y(n_405) );
BUFx2_ASAP7_75t_L g457 ( .A(n_244), .Y(n_457) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g488 ( .A(n_246), .B(n_400), .Y(n_488) );
INVx2_ASAP7_75t_L g282 ( .A(n_247), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_249), .B(n_255), .Y(n_248) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_269), .Y(n_257) );
AND2x2_ASAP7_75t_L g304 ( .A(n_258), .B(n_305), .Y(n_304) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_SL g289 ( .A(n_259), .B(n_279), .Y(n_289) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g277 ( .A(n_260), .Y(n_277) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_260), .Y(n_383) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_260), .Y(n_450) );
INVx1_ASAP7_75t_L g490 ( .A(n_260), .Y(n_490) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B(n_268), .Y(n_260) );
AO21x2_ASAP7_75t_L g582 ( .A1(n_261), .A2(n_583), .B(n_589), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
BUFx2_ASAP7_75t_L g404 ( .A(n_269), .Y(n_404) );
NOR2x1_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
AND2x4_ASAP7_75t_L g320 ( .A(n_270), .B(n_321), .Y(n_320) );
NOR2xp67_ASAP7_75t_SL g352 ( .A(n_270), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g425 ( .A(n_270), .B(n_408), .Y(n_425) );
AND2x4_ASAP7_75t_SL g428 ( .A(n_270), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g477 ( .A(n_270), .B(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g344 ( .A(n_271), .Y(n_344) );
INVx4_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g339 ( .A(n_272), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_272), .B(n_337), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_272), .B(n_397), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_272), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2x1_ASAP7_75t_L g274 ( .A(n_275), .B(n_278), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g422 ( .A(n_276), .B(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g338 ( .A(n_277), .Y(n_338) );
NAND2x1p5_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
AND2x2_ASAP7_75t_L g456 ( .A(n_281), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g464 ( .A(n_281), .B(n_393), .Y(n_464) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g333 ( .A(n_282), .B(n_318), .Y(n_333) );
AND2x4_ASAP7_75t_L g366 ( .A(n_282), .B(n_300), .Y(n_366) );
INVx1_ASAP7_75t_L g483 ( .A(n_282), .Y(n_483) );
AND2x2_ASAP7_75t_L g369 ( .A(n_284), .B(n_309), .Y(n_369) );
INVx2_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g390 ( .A(n_285), .B(n_325), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_294), .B1(n_303), .B2(n_306), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .B(n_292), .Y(n_287) );
OAI22xp5_ASAP7_75t_SL g469 ( .A1(n_288), .A2(n_357), .B1(n_465), .B2(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_289), .B(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g358 ( .A(n_289), .B(n_290), .Y(n_358) );
AND2x2_ASAP7_75t_SL g388 ( .A(n_289), .B(n_360), .Y(n_388) );
AOI211xp5_ASAP7_75t_SL g476 ( .A1(n_289), .A2(n_477), .B(n_479), .C(n_480), .Y(n_476) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_290), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_290), .B(n_336), .Y(n_462) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g367 ( .A(n_292), .Y(n_367) );
INVx2_ASAP7_75t_L g423 ( .A(n_293), .Y(n_423) );
AND2x2_ASAP7_75t_L g497 ( .A(n_293), .B(n_490), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_294), .A2(n_446), .B(n_452), .Y(n_445) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_299), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g432 ( .A(n_296), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g442 ( .A(n_296), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g349 ( .A(n_297), .B(n_302), .Y(n_349) );
NOR2xp67_ASAP7_75t_L g351 ( .A(n_297), .B(n_318), .Y(n_351) );
AND2x2_ASAP7_75t_L g393 ( .A(n_297), .B(n_318), .Y(n_393) );
INVx2_ASAP7_75t_L g310 ( .A(n_298), .Y(n_310) );
AND2x4_ASAP7_75t_L g316 ( .A(n_298), .B(n_317), .Y(n_316) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx3_ASAP7_75t_L g308 ( .A(n_300), .Y(n_308) );
INVx3_ASAP7_75t_L g314 ( .A(n_301), .Y(n_314) );
BUFx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_305), .A2(n_411), .B(n_487), .Y(n_491) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g323 ( .A(n_308), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_308), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_308), .B(n_383), .Y(n_398) );
OR2x2_ASAP7_75t_L g413 ( .A(n_308), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g420 ( .A(n_308), .B(n_324), .Y(n_420) );
AND2x2_ASAP7_75t_L g376 ( .A(n_309), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g392 ( .A(n_309), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g409 ( .A(n_309), .B(n_378), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_319), .B1(n_322), .B2(n_326), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NOR2xp67_ASAP7_75t_L g386 ( .A(n_314), .B(n_315), .Y(n_386) );
NOR2xp67_ASAP7_75t_SL g424 ( .A(n_314), .B(n_332), .Y(n_424) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2x1_ASAP7_75t_L g443 ( .A(n_318), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g327 ( .A(n_320), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g391 ( .A(n_320), .B(n_337), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_320), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g494 ( .A(n_328), .B(n_360), .Y(n_494) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NOR2x1_ASAP7_75t_L g439 ( .A(n_329), .B(n_440), .Y(n_439) );
NOR2xp67_ASAP7_75t_SL g330 ( .A(n_331), .B(n_354), .Y(n_330) );
OAI211xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B(n_341), .C(n_350), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_L g394 ( .A1(n_332), .A2(n_385), .B(n_395), .C(n_399), .Y(n_394) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g474 ( .A(n_333), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g385 ( .A(n_337), .B(n_361), .Y(n_385) );
AND2x2_ASAP7_75t_L g472 ( .A(n_337), .B(n_451), .Y(n_472) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g440 ( .A(n_340), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_347), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2x1_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_344), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g414 ( .A(n_349), .Y(n_414) );
NAND2xp33_ASAP7_75t_SL g350 ( .A(n_351), .B(n_352), .Y(n_350) );
OAI221xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_362), .B1(n_364), .B2(n_367), .C(n_368), .Y(n_354) );
NOR4xp25_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .C(n_359), .D(n_361), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g473 ( .A(n_360), .B(n_436), .Y(n_473) );
INVx2_ASAP7_75t_L g479 ( .A(n_360), .Y(n_479) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_363), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g466 ( .A(n_366), .B(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND4xp75_ASAP7_75t_L g371 ( .A(n_372), .B(n_394), .C(n_401), .D(n_410), .Y(n_371) );
OA211x2_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_375), .B(n_379), .C(n_387), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_373), .B(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g467 ( .A(n_377), .Y(n_467) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g475 ( .A(n_378), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_380), .B(n_386), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_384), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g436 ( .A(n_383), .Y(n_436) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_391), .B2(n_392), .Y(n_387) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_391), .A2(n_442), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_SL g470 ( .A(n_392), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_393), .B(n_483), .Y(n_482) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NOR2x1_ASAP7_75t_L g401 ( .A(n_402), .B(n_406), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVxp67_ASAP7_75t_L g468 ( .A(n_404), .Y(n_468) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
AND2x2_ASAP7_75t_SL g427 ( .A(n_408), .B(n_428), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_409), .A2(n_472), .B1(n_494), .B2(n_495), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND3x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_458), .C(n_471), .Y(n_416) );
NOR3x1_ASAP7_75t_L g417 ( .A(n_418), .B(n_430), .C(n_445), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_426), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_424), .B2(n_425), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_435), .B1(n_437), .B2(n_441), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g489 ( .A(n_439), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g478 ( .A(n_455), .Y(n_478) );
OAI21xp5_ASAP7_75t_SL g486 ( .A1(n_456), .A2(n_487), .B(n_489), .Y(n_486) );
NOR2x1_ASAP7_75t_L g458 ( .A(n_459), .B(n_469), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .B1(n_465), .B2(n_468), .Y(n_459) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
O2A1O1Ixp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_474), .C(n_476), .Y(n_471) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NOR2x1_ASAP7_75t_SL g484 ( .A(n_485), .B(n_492), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_491), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_493), .B(n_496), .Y(n_492) );
INVx4_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
CKINVDCx11_ASAP7_75t_R g808 ( .A(n_499), .Y(n_808) );
INVx3_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g807 ( .A(n_502), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_502), .A2(n_817), .B1(n_818), .B2(n_821), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_502), .Y(n_817) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_701), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_638), .C(n_661), .Y(n_503) );
NAND3xp33_ASAP7_75t_SL g504 ( .A(n_505), .B(n_590), .C(n_607), .Y(n_504) );
OAI31xp33_ASAP7_75t_SL g505 ( .A1(n_506), .A2(n_526), .A3(n_546), .B(n_553), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_506), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_520), .Y(n_507) );
AND2x4_ASAP7_75t_L g593 ( .A(n_508), .B(n_520), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_508), .B(n_537), .Y(n_622) );
AND2x4_ASAP7_75t_L g624 ( .A(n_508), .B(n_618), .Y(n_624) );
AND2x2_ASAP7_75t_L g755 ( .A(n_508), .B(n_550), .Y(n_755) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g600 ( .A(n_509), .Y(n_600) );
OAI21x1_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_513), .B(n_518), .Y(n_509) );
INVx1_ASAP7_75t_L g519 ( .A(n_512), .Y(n_519) );
AND2x2_ASAP7_75t_L g536 ( .A(n_520), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_SL g691 ( .A(n_520), .B(n_599), .Y(n_691) );
AND2x2_ASAP7_75t_L g697 ( .A(n_520), .B(n_538), .Y(n_697) );
AND2x2_ASAP7_75t_L g786 ( .A(n_520), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_SL g768 ( .A(n_526), .Y(n_768) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_536), .Y(n_526) );
BUFx2_ASAP7_75t_L g597 ( .A(n_527), .Y(n_597) );
AND2x2_ASAP7_75t_L g631 ( .A(n_527), .B(n_537), .Y(n_631) );
AND2x2_ASAP7_75t_L g680 ( .A(n_527), .B(n_538), .Y(n_680) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g637 ( .A(n_528), .B(n_538), .Y(n_637) );
INVxp67_ASAP7_75t_L g649 ( .A(n_528), .Y(n_649) );
BUFx3_ASAP7_75t_L g694 ( .A(n_528), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_534), .Y(n_529) );
OAI31xp33_ASAP7_75t_L g590 ( .A1(n_536), .A2(n_591), .A3(n_596), .B(n_601), .Y(n_590) );
AND2x2_ASAP7_75t_L g598 ( .A(n_537), .B(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g617 ( .A(n_538), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_540), .B(n_544), .Y(n_539) );
AOI322xp5_ASAP7_75t_L g791 ( .A1(n_546), .A2(n_666), .A3(n_695), .B1(n_700), .B2(n_792), .C1(n_795), .C2(n_796), .Y(n_791) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_547), .B(n_637), .Y(n_642) );
NAND2x1_ASAP7_75t_L g679 ( .A(n_547), .B(n_680), .Y(n_679) );
AND2x4_ASAP7_75t_L g723 ( .A(n_547), .B(n_627), .Y(n_723) );
INVx1_ASAP7_75t_SL g737 ( .A(n_547), .Y(n_737) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g618 ( .A(n_548), .Y(n_618) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_548), .Y(n_761) );
AND2x2_ASAP7_75t_L g690 ( .A(n_549), .B(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_549), .B(n_737), .Y(n_736) );
AND2x4_ASAP7_75t_SL g549 ( .A(n_550), .B(n_551), .Y(n_549) );
BUFx2_ASAP7_75t_L g595 ( .A(n_550), .Y(n_595) );
INVx1_ASAP7_75t_L g787 ( .A(n_550), .Y(n_787) );
OR2x2_ASAP7_75t_L g654 ( .A(n_551), .B(n_599), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_551), .B(n_624), .Y(n_688) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g627 ( .A(n_552), .B(n_599), .Y(n_627) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_573), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g683 ( .A(n_555), .Y(n_683) );
OR2x2_ASAP7_75t_L g710 ( .A(n_555), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_566), .Y(n_555) );
NOR2x1_ASAP7_75t_SL g604 ( .A(n_556), .B(n_574), .Y(n_604) );
AND2x2_ASAP7_75t_L g611 ( .A(n_556), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g783 ( .A(n_556), .B(n_645), .Y(n_783) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_564), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_557), .B(n_565), .Y(n_564) );
AO21x2_ASAP7_75t_L g660 ( .A1(n_557), .A2(n_558), .B(n_564), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_563), .Y(n_558) );
OR2x2_ASAP7_75t_L g605 ( .A(n_566), .B(n_606), .Y(n_605) );
BUFx3_ASAP7_75t_L g614 ( .A(n_566), .Y(n_614) );
INVx2_ASAP7_75t_L g645 ( .A(n_566), .Y(n_645) );
INVx1_ASAP7_75t_L g686 ( .A(n_566), .Y(n_686) );
AND2x2_ASAP7_75t_L g717 ( .A(n_566), .B(n_574), .Y(n_717) );
AND2x2_ASAP7_75t_L g748 ( .A(n_566), .B(n_675), .Y(n_748) );
AND2x2_ASAP7_75t_L g644 ( .A(n_573), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_573), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_SL g747 ( .A(n_573), .B(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g752 ( .A(n_573), .B(n_614), .Y(n_752) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_582), .Y(n_573) );
INVx5_ASAP7_75t_L g612 ( .A(n_574), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_574), .B(n_606), .Y(n_684) );
BUFx2_ASAP7_75t_L g744 ( .A(n_574), .Y(n_744) );
OR2x6_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx4_ASAP7_75t_L g606 ( .A(n_582), .Y(n_606) );
AND2x2_ASAP7_75t_L g729 ( .A(n_582), .B(n_612), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_588), .Y(n_583) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OAI221xp5_ASAP7_75t_L g718 ( .A1(n_592), .A2(n_719), .B1(n_722), .B2(n_724), .C(n_725), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g740 ( .A(n_593), .B(n_631), .Y(n_740) );
INVx1_ASAP7_75t_SL g766 ( .A(n_593), .Y(n_766) );
AND2x2_ASAP7_75t_L g751 ( .A(n_594), .B(n_723), .Y(n_751) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_595), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AND2x2_ASAP7_75t_L g620 ( .A(n_597), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g626 ( .A(n_597), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g650 ( .A(n_598), .Y(n_650) );
AND2x2_ASAP7_75t_L g708 ( .A(n_598), .B(n_636), .Y(n_708) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx2_ASAP7_75t_L g633 ( .A(n_600), .Y(n_633) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g629 ( .A(n_605), .Y(n_629) );
OR2x2_ASAP7_75t_L g797 ( .A(n_605), .B(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g613 ( .A(n_606), .Y(n_613) );
AND2x4_ASAP7_75t_L g669 ( .A(n_606), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_606), .B(n_674), .Y(n_673) );
NAND2x1p5_ASAP7_75t_L g711 ( .A(n_606), .B(n_612), .Y(n_711) );
AND2x2_ASAP7_75t_L g771 ( .A(n_606), .B(n_674), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_615), .B1(n_628), .B2(n_630), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_608), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND3x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .C(n_614), .Y(n_610) );
AND2x4_ASAP7_75t_L g628 ( .A(n_611), .B(n_629), .Y(n_628) );
INVx4_ASAP7_75t_L g668 ( .A(n_612), .Y(n_668) );
AND2x2_ASAP7_75t_SL g801 ( .A(n_612), .B(n_669), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_613), .B(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g713 ( .A(n_614), .Y(n_713) );
AOI322xp5_ASAP7_75t_L g778 ( .A1(n_614), .A2(n_743), .A3(n_779), .B1(n_781), .B2(n_784), .C1(n_788), .C2(n_789), .Y(n_778) );
NAND4xp25_ASAP7_75t_SL g615 ( .A(n_616), .B(n_619), .C(n_623), .D(n_625), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_SL g745 ( .A(n_617), .B(n_633), .Y(n_745) );
BUFx2_ASAP7_75t_L g636 ( .A(n_618), .Y(n_636) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g760 ( .A(n_621), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g774 ( .A(n_622), .B(n_649), .Y(n_774) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g640 ( .A(n_624), .B(n_641), .Y(n_640) );
OAI211xp5_ASAP7_75t_L g692 ( .A1(n_624), .A2(n_693), .B(n_695), .C(n_698), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_624), .B(n_631), .Y(n_750) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_626), .A2(n_708), .B1(n_709), .B2(n_712), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_627), .A2(n_663), .B1(n_667), .B2(n_671), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_627), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_627), .B(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_627), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g794 ( .A(n_627), .Y(n_794) );
INVx1_ASAP7_75t_L g733 ( .A(n_628), .Y(n_733) );
OAI21xp33_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_632), .B(n_634), .Y(n_630) );
INVx1_ASAP7_75t_L g641 ( .A(n_631), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_631), .B(n_636), .Y(n_790) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g726 ( .A(n_633), .B(n_637), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_635), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g793 ( .A(n_636), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g767 ( .A(n_637), .Y(n_767) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_642), .B(n_643), .C(n_646), .Y(n_638) );
INVxp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp33_ASAP7_75t_SL g753 ( .A1(n_641), .A2(n_672), .B1(n_719), .B2(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_645), .B(n_668), .Y(n_676) );
OR2x2_ASAP7_75t_L g705 ( .A(n_645), .B(n_706), .Y(n_705) );
OAI21xp5_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_651), .B(n_655), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g666 ( .A(n_649), .Y(n_666) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI211xp5_ASAP7_75t_SL g704 ( .A1(n_652), .A2(n_705), .B(n_707), .C(n_715), .Y(n_704) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp67_ASAP7_75t_SL g738 ( .A(n_657), .B(n_684), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_657), .Y(n_741) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_659), .B(n_668), .Y(n_798) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g670 ( .A(n_660), .Y(n_670) );
INVx2_ASAP7_75t_L g675 ( .A(n_660), .Y(n_675) );
NAND4xp25_ASAP7_75t_L g661 ( .A(n_662), .B(n_677), .C(n_689), .D(n_692), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g796 ( .A1(n_665), .A2(n_797), .B1(n_799), .B2(n_800), .Y(n_796) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
AND2x4_ASAP7_75t_L g764 ( .A(n_668), .B(n_694), .Y(n_764) );
AND2x2_ASAP7_75t_L g685 ( .A(n_669), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g706 ( .A(n_669), .Y(n_706) );
AND2x2_ASAP7_75t_L g716 ( .A(n_669), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_676), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_675), .Y(n_730) );
INVx1_ASAP7_75t_L g720 ( .A(n_676), .Y(n_720) );
AOI32xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_681), .A3(n_684), .B1(n_685), .B2(n_687), .Y(n_677) );
OAI21xp33_ASAP7_75t_L g725 ( .A1(n_678), .A2(n_726), .B(n_727), .Y(n_725) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g757 ( .A1(n_681), .A2(n_758), .B1(n_760), .B2(n_762), .C(n_765), .Y(n_757) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g742 ( .A(n_683), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g700 ( .A(n_684), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_685), .A2(n_723), .B1(n_773), .B2(n_775), .Y(n_772) );
INVx1_ASAP7_75t_L g699 ( .A(n_686), .Y(n_699) );
AND2x2_ASAP7_75t_L g777 ( .A(n_686), .B(n_730), .Y(n_777) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g780 ( .A(n_693), .B(n_745), .Y(n_780) );
INVx1_ASAP7_75t_L g799 ( .A(n_693), .Y(n_799) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
NOR2xp67_ASAP7_75t_L g701 ( .A(n_702), .B(n_756), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_746), .Y(n_702) );
NOR3xp33_ASAP7_75t_SL g703 ( .A(n_704), .B(n_718), .C(n_731), .Y(n_703) );
INVx1_ASAP7_75t_L g721 ( .A(n_706), .Y(n_721) );
INVx1_ASAP7_75t_SL g732 ( .A(n_708), .Y(n_732) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g714 ( .A(n_711), .Y(n_714) );
INVx2_ASAP7_75t_L g724 ( .A(n_712), .Y(n_724) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
AND2x4_ASAP7_75t_L g770 ( .A(n_713), .B(n_771), .Y(n_770) );
AND2x4_ASAP7_75t_L g788 ( .A(n_717), .B(n_771), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .Y(n_727) );
AOI32xp33_ASAP7_75t_L g739 ( .A1(n_728), .A2(n_740), .A3(n_741), .B1(n_742), .B2(n_745), .Y(n_739) );
NOR2xp33_ASAP7_75t_SL g758 ( .A(n_728), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g759 ( .A(n_730), .Y(n_759) );
OAI211xp5_ASAP7_75t_SL g731 ( .A1(n_732), .A2(n_733), .B(n_734), .C(n_739), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_738), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g795 ( .A(n_743), .B(n_783), .Y(n_795) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_744), .B(n_783), .Y(n_782) );
AOI221xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_749), .B1(n_751), .B2(n_752), .C(n_753), .Y(n_746) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
CKINVDCx16_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
NAND4xp25_ASAP7_75t_L g756 ( .A(n_757), .B(n_772), .C(n_778), .D(n_791), .Y(n_756) );
INVxp33_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
O2A1O1Ixp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_767), .B(n_768), .C(n_769), .Y(n_765) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx3_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g821 ( .A(n_818), .Y(n_821) );
INVx1_ASAP7_75t_SL g822 ( .A(n_823), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_SL g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g835 ( .A(n_827), .Y(n_835) );
NAND2xp5_ASAP7_75t_SL g827 ( .A(n_828), .B(n_830), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .Y(n_833) );
endmodule