module fake_jpeg_25729_n_223 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_223);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_223;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_24),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_26),
.B1(n_27),
.B2(n_18),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_43),
.A2(n_41),
.B1(n_38),
.B2(n_35),
.Y(n_81)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_54),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_18),
.B1(n_27),
.B2(n_25),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_41),
.B1(n_38),
.B2(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_58),
.B(n_59),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_48),
.B1(n_35),
.B2(n_33),
.Y(n_92)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_72),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_21),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_78),
.Y(n_89)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_74),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_80),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_28),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_28),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_66),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_67),
.B1(n_63),
.B2(n_38),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_40),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_107),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_36),
.B1(n_32),
.B2(n_17),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_49),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_37),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_40),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_109),
.B(n_115),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_62),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_118),
.C(n_122),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_62),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_117),
.B(n_124),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_59),
.Y(n_113)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_72),
.Y(n_116)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_89),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_22),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_17),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_121),
.Y(n_149)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_24),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_127),
.B1(n_100),
.B2(n_69),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_129),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_82),
.B1(n_69),
.B2(n_60),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_32),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_98),
.B(n_74),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_96),
.B(n_44),
.Y(n_132)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_141),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_97),
.B(n_102),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_112),
.B(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_92),
.B1(n_97),
.B2(n_102),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_33),
.B1(n_108),
.B2(n_88),
.Y(n_161)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_147),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_100),
.B1(n_33),
.B2(n_60),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_108),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_154),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_112),
.B(n_114),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_88),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_114),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_156),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_122),
.B(n_111),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_118),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_160),
.Y(n_175)
);

OAI322xp33_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_21),
.A3(n_16),
.B1(n_30),
.B2(n_14),
.C1(n_15),
.C2(n_9),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_164),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_137),
.B(n_136),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_151),
.B1(n_139),
.B2(n_146),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_170),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_44),
.C(n_30),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_30),
.C(n_16),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_172),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_0),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_178),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_144),
.B1(n_133),
.B2(n_141),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_177),
.A2(n_166),
.B1(n_173),
.B2(n_172),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_157),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_137),
.B1(n_171),
.B2(n_167),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_182),
.A2(n_135),
.B(n_140),
.Y(n_196)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_177),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_162),
.B(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_191),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_158),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_193),
.Y(n_198)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_173),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_136),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_196),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_200),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_138),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_204),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_183),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_205),
.Y(n_209)
);

OAI322xp33_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_175),
.A3(n_168),
.B1(n_183),
.B2(n_181),
.C1(n_13),
.C2(n_11),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_181),
.C(n_175),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_194),
.B1(n_186),
.B2(n_11),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_202),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_0),
.B(n_2),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_2),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_213),
.A2(n_215),
.B1(n_209),
.B2(n_4),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_206),
.B(n_198),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_2),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_211),
.C(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

AOI322xp5_ASAP7_75t_L g221 ( 
.A1(n_219),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_209),
.C1(n_216),
.C2(n_211),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_221),
.A2(n_220),
.B1(n_217),
.B2(n_5),
.Y(n_222)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_222),
.Y(n_223)
);


endmodule