module fake_ariane_1765_n_14789 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_14789);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_14789;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_9872;
wire n_14741;
wire n_9604;
wire n_10943;
wire n_10453;
wire n_12407;
wire n_7329;
wire n_4030;
wire n_12343;
wire n_13909;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_14469;
wire n_11913;
wire n_8165;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_12760;
wire n_11172;
wire n_12018;
wire n_14470;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_10678;
wire n_5402;
wire n_11190;
wire n_13957;
wire n_6581;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_11458;
wire n_2680;
wire n_7277;
wire n_11999;
wire n_3264;
wire n_1250;
wire n_10649;
wire n_13176;
wire n_5717;
wire n_10794;
wire n_12945;
wire n_2993;
wire n_4283;
wire n_9297;
wire n_11627;
wire n_2879;
wire n_4403;
wire n_10557;
wire n_13125;
wire n_8139;
wire n_11453;
wire n_416;
wire n_4962;
wire n_1430;
wire n_14456;
wire n_7832;
wire n_8438;
wire n_2002;
wire n_12806;
wire n_12244;
wire n_11306;
wire n_1238;
wire n_11135;
wire n_2729;
wire n_4302;
wire n_14658;
wire n_12589;
wire n_5791;
wire n_7127;
wire n_13109;
wire n_4547;
wire n_14209;
wire n_13718;
wire n_5090;
wire n_3765;
wire n_8321;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_10000;
wire n_2376;
wire n_12103;
wire n_7922;
wire n_7805;
wire n_9807;
wire n_2790;
wire n_7542;
wire n_12354;
wire n_2207;
wire n_11783;
wire n_7053;
wire n_11614;
wire n_9892;
wire n_5712;
wire n_11143;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_10704;
wire n_14334;
wire n_11431;
wire n_11799;
wire n_462;
wire n_8699;
wire n_9263;
wire n_9734;
wire n_1131;
wire n_8037;
wire n_5479;
wire n_2646;
wire n_8257;
wire n_737;
wire n_2653;
wire n_4610;
wire n_11377;
wire n_11246;
wire n_10213;
wire n_6058;
wire n_232;
wire n_13029;
wire n_3115;
wire n_9886;
wire n_4028;
wire n_5263;
wire n_10904;
wire n_9096;
wire n_5565;
wire n_6358;
wire n_8546;
wire n_6293;
wire n_8997;
wire n_13215;
wire n_14066;
wire n_2482;
wire n_9985;
wire n_9665;
wire n_1682;
wire n_14300;
wire n_12233;
wire n_11349;
wire n_7001;
wire n_10169;
wire n_10903;
wire n_13875;
wire n_11906;
wire n_958;
wire n_6129;
wire n_13755;
wire n_14335;
wire n_2554;
wire n_14473;
wire n_13910;
wire n_4321;
wire n_10574;
wire n_13066;
wire n_1985;
wire n_5590;
wire n_10468;
wire n_2621;
wire n_14226;
wire n_9241;
wire n_146;
wire n_6524;
wire n_9286;
wire n_4853;
wire n_8744;
wire n_338;
wire n_9592;
wire n_1909;
wire n_5229;
wire n_12574;
wire n_6313;
wire n_12260;
wire n_7464;
wire n_8449;
wire n_9683;
wire n_10380;
wire n_10968;
wire n_4260;
wire n_13491;
wire n_903;
wire n_7626;
wire n_9939;
wire n_3348;
wire n_239;
wire n_12315;
wire n_10688;
wire n_3261;
wire n_9358;
wire n_1761;
wire n_9466;
wire n_8953;
wire n_11756;
wire n_7965;
wire n_13636;
wire n_7368;
wire n_9787;
wire n_1690;
wire n_8399;
wire n_2807;
wire n_6664;
wire n_8598;
wire n_10276;
wire n_7562;
wire n_11604;
wire n_9997;
wire n_7534;
wire n_13196;
wire n_1018;
wire n_7428;
wire n_12581;
wire n_4512;
wire n_6190;
wire n_8460;
wire n_12085;
wire n_4132;
wire n_13980;
wire n_1364;
wire n_8068;
wire n_2390;
wire n_7373;
wire n_6891;
wire n_4500;
wire n_9318;
wire n_10281;
wire n_13715;
wire n_12089;
wire n_625;
wire n_2322;
wire n_8734;
wire n_12671;
wire n_1107;
wire n_14592;
wire n_8720;
wire n_331;
wire n_559;
wire n_2663;
wire n_10528;
wire n_8097;
wire n_5481;
wire n_6539;
wire n_12993;
wire n_13120;
wire n_495;
wire n_8114;
wire n_4824;
wire n_8422;
wire n_12728;
wire n_7467;
wire n_14572;
wire n_350;
wire n_8126;
wire n_381;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_7392;
wire n_9714;
wire n_14405;
wire n_14598;
wire n_10399;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_7526;
wire n_8664;
wire n_10131;
wire n_11721;
wire n_14378;
wire n_561;
wire n_11736;
wire n_4143;
wire n_14430;
wire n_10634;
wire n_4273;
wire n_507;
wire n_11444;
wire n_901;
wire n_11891;
wire n_13058;
wire n_4136;
wire n_14094;
wire n_9809;
wire n_11492;
wire n_3144;
wire n_14636;
wire n_2359;
wire n_9613;
wire n_9354;
wire n_1519;
wire n_5896;
wire n_7338;
wire n_4567;
wire n_12647;
wire n_9897;
wire n_786;
wire n_9295;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_10595;
wire n_11767;
wire n_13180;
wire n_6253;
wire n_9119;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_9058;
wire n_6197;
wire n_8326;
wire n_7200;
wire n_11807;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_11944;
wire n_2301;
wire n_13090;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_11474;
wire n_11819;
wire n_8504;
wire n_3015;
wire n_5744;
wire n_8920;
wire n_3870;
wire n_12080;
wire n_6808;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_277;
wire n_5691;
wire n_7937;
wire n_8985;
wire n_3482;
wire n_7490;
wire n_13069;
wire n_6295;
wire n_11409;
wire n_5403;
wire n_823;
wire n_11692;
wire n_1900;
wire n_620;
wire n_13138;
wire n_12599;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_587;
wire n_863;
wire n_6992;
wire n_303;
wire n_3960;
wire n_10644;
wire n_12863;
wire n_2433;
wire n_352;
wire n_899;
wire n_3975;
wire n_8035;
wire n_11856;
wire n_5830;
wire n_9516;
wire n_365;
wire n_2004;
wire n_13996;
wire n_13064;
wire n_4018;
wire n_1495;
wire n_8660;
wire n_334;
wire n_192;
wire n_3325;
wire n_6681;
wire n_661;
wire n_4227;
wire n_5158;
wire n_9917;
wire n_12185;
wire n_5152;
wire n_8939;
wire n_11737;
wire n_533;
wire n_11652;
wire n_11038;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_13991;
wire n_1924;
wire n_6542;
wire n_13466;
wire n_9202;
wire n_13689;
wire n_13896;
wire n_11925;
wire n_1811;
wire n_14115;
wire n_6161;
wire n_3612;
wire n_273;
wire n_4505;
wire n_11974;
wire n_12457;
wire n_6452;
wire n_10426;
wire n_1840;
wire n_5247;
wire n_9512;
wire n_9923;
wire n_8469;
wire n_8715;
wire n_5464;
wire n_7306;
wire n_10070;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_12792;
wire n_579;
wire n_7507;
wire n_13458;
wire n_844;
wire n_1267;
wire n_8176;
wire n_9677;
wire n_2956;
wire n_5210;
wire n_7215;
wire n_149;
wire n_1213;
wire n_2382;
wire n_7441;
wire n_7379;
wire n_237;
wire n_780;
wire n_5292;
wire n_1918;
wire n_12556;
wire n_8327;
wire n_8991;
wire n_7438;
wire n_11200;
wire n_8855;
wire n_4119;
wire n_4443;
wire n_9811;
wire n_4000;
wire n_13762;
wire n_9508;
wire n_13441;
wire n_13532;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_1140;
wire n_14236;
wire n_3458;
wire n_570;
wire n_11597;
wire n_5843;
wire n_7874;
wire n_11309;
wire n_14156;
wire n_8539;
wire n_13118;
wire n_8630;
wire n_9308;
wire n_14587;
wire n_8533;
wire n_13830;
wire n_11233;
wire n_11047;
wire n_3511;
wire n_2077;
wire n_9638;
wire n_1121;
wire n_7108;
wire n_11068;
wire n_490;
wire n_3012;
wire n_13912;
wire n_1947;
wire n_13768;
wire n_4529;
wire n_3850;
wire n_575;
wire n_11476;
wire n_8435;
wire n_7695;
wire n_10245;
wire n_6156;
wire n_11611;
wire n_13111;
wire n_1216;
wire n_4908;
wire n_8098;
wire n_3754;
wire n_11957;
wire n_8204;
wire n_5060;
wire n_13290;
wire n_12509;
wire n_12663;
wire n_9199;
wire n_12155;
wire n_13379;
wire n_7162;
wire n_4432;
wire n_11210;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_9808;
wire n_7331;
wire n_10457;
wire n_5913;
wire n_8958;
wire n_13838;
wire n_4530;
wire n_11333;
wire n_11682;
wire n_9821;
wire n_1432;
wire n_2245;
wire n_13692;
wire n_5614;
wire n_5452;
wire n_5391;
wire n_10715;
wire n_11381;
wire n_3359;
wire n_7944;
wire n_3841;
wire n_11922;
wire n_5249;
wire n_13126;
wire n_249;
wire n_14762;
wire n_851;
wire n_12068;
wire n_444;
wire n_10579;
wire n_3900;
wire n_3413;
wire n_7850;
wire n_5076;
wire n_10707;
wire n_3539;
wire n_5757;
wire n_9265;
wire n_6872;
wire n_12332;
wire n_12858;
wire n_6644;
wire n_11352;
wire n_9143;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_12641;
wire n_930;
wire n_4912;
wire n_12140;
wire n_9845;
wire n_4226;
wire n_10112;
wire n_14505;
wire n_10556;
wire n_14150;
wire n_4311;
wire n_3284;
wire n_8542;
wire n_8572;
wire n_5046;
wire n_7607;
wire n_14292;
wire n_13330;
wire n_7642;
wire n_8373;
wire n_8424;
wire n_13417;
wire n_8442;
wire n_1386;
wire n_9304;
wire n_14492;
wire n_6236;
wire n_8147;
wire n_7104;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_11152;
wire n_13505;
wire n_1842;
wire n_7397;
wire n_4993;
wire n_3678;
wire n_7205;
wire n_10080;
wire n_366;
wire n_2791;
wire n_1661;
wire n_555;
wire n_3212;
wire n_11022;
wire n_4871;
wire n_11025;
wire n_12517;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_11251;
wire n_966;
wire n_992;
wire n_3549;
wire n_13821;
wire n_3914;
wire n_10766;
wire n_13787;
wire n_6398;
wire n_11222;
wire n_5586;
wire n_14065;
wire n_7461;
wire n_8519;
wire n_1692;
wire n_11650;
wire n_14310;
wire n_2611;
wire n_8075;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_7638;
wire n_10781;
wire n_2398;
wire n_11091;
wire n_13243;
wire n_4233;
wire n_4791;
wire n_8642;
wire n_6319;
wire n_5971;
wire n_11713;
wire n_8648;
wire n_10217;
wire n_7224;
wire n_6966;
wire n_9791;
wire n_5056;
wire n_9449;
wire n_9934;
wire n_9149;
wire n_9686;
wire n_13063;
wire n_1178;
wire n_2015;
wire n_13186;
wire n_14639;
wire n_13463;
wire n_7259;
wire n_8556;
wire n_7838;
wire n_5984;
wire n_12961;
wire n_14039;
wire n_11398;
wire n_9844;
wire n_5204;
wire n_6724;
wire n_6705;
wire n_12389;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_11208;
wire n_203;
wire n_9458;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_150;
wire n_2930;
wire n_7840;
wire n_8585;
wire n_9717;
wire n_11858;
wire n_12595;
wire n_11487;
wire n_14194;
wire n_2745;
wire n_8455;
wire n_2087;
wire n_8444;
wire n_13237;
wire n_619;
wire n_9128;
wire n_14788;
wire n_10638;
wire n_14559;
wire n_14255;
wire n_2161;
wire n_11745;
wire n_10239;
wire n_746;
wire n_12368;
wire n_13353;
wire n_6624;
wire n_1357;
wire n_7888;
wire n_8560;
wire n_292;
wire n_12816;
wire n_14730;
wire n_11525;
wire n_6710;
wire n_1787;
wire n_6883;
wire n_9558;
wire n_8108;
wire n_1389;
wire n_8158;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_10464;
wire n_13054;
wire n_3747;
wire n_10446;
wire n_6553;
wire n_9715;
wire n_14166;
wire n_4905;
wire n_10219;
wire n_9016;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_6659;
wire n_9399;
wire n_6261;
wire n_428;
wire n_7351;
wire n_3614;
wire n_7256;
wire n_959;
wire n_12967;
wire n_2257;
wire n_14458;
wire n_1101;
wire n_1343;
wire n_12907;
wire n_14353;
wire n_3116;
wire n_12020;
wire n_4141;
wire n_13877;
wire n_3784;
wire n_6893;
wire n_12377;
wire n_3891;
wire n_3372;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_12007;
wire n_13272;
wire n_11087;
wire n_8814;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_2435;
wire n_10394;
wire n_6337;
wire n_6210;
wire n_1932;
wire n_7583;
wire n_5680;
wire n_1780;
wire n_14368;
wire n_2825;
wire n_5685;
wire n_13394;
wire n_5974;
wire n_10776;
wire n_14032;
wire n_14375;
wire n_10917;
wire n_5723;
wire n_542;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_1087;
wire n_13536;
wire n_632;
wire n_9094;
wire n_2388;
wire n_13524;
wire n_2273;
wire n_8130;
wire n_1911;
wire n_11483;
wire n_14075;
wire n_3496;
wire n_14093;
wire n_4364;
wire n_3493;
wire n_12944;
wire n_14705;
wire n_9510;
wire n_11049;
wire n_7488;
wire n_3700;
wire n_7690;
wire n_12706;
wire n_12973;
wire n_12319;
wire n_6076;
wire n_4307;
wire n_14178;
wire n_2795;
wire n_14053;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_12388;
wire n_6206;
wire n_7893;
wire n_2954;
wire n_11031;
wire n_382;
wire n_9429;
wire n_489;
wire n_11599;
wire n_4438;
wire n_11292;
wire n_6538;
wire n_11568;
wire n_7966;
wire n_251;
wire n_974;
wire n_506;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_9653;
wire n_4367;
wire n_5134;
wire n_11468;
wire n_13815;
wire n_2467;
wire n_7599;
wire n_9648;
wire n_7231;
wire n_14626;
wire n_10240;
wire n_4195;
wire n_7007;
wire n_7717;
wire n_6579;
wire n_12470;
wire n_12711;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_1447;
wire n_8675;
wire n_1220;
wire n_12216;
wire n_9095;
wire n_7900;
wire n_11203;
wire n_2019;
wire n_5708;
wire n_8123;
wire n_698;
wire n_9048;
wire n_9003;
wire n_12879;
wire n_14228;
wire n_13801;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_14472;
wire n_13659;
wire n_307;
wire n_1209;
wire n_4254;
wire n_10578;
wire n_11206;
wire n_646;
wire n_12649;
wire n_12093;
wire n_13473;
wire n_8913;
wire n_9932;
wire n_3438;
wire n_8220;
wire n_12165;
wire n_404;
wire n_2625;
wire n_11779;
wire n_13497;
wire n_9309;
wire n_8355;
wire n_12724;
wire n_9661;
wire n_14557;
wire n_9799;
wire n_12447;
wire n_5373;
wire n_7403;
wire n_1578;
wire n_6665;
wire n_8883;
wire n_3147;
wire n_13822;
wire n_299;
wire n_3661;
wire n_7168;
wire n_10427;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_11609;
wire n_11927;
wire n_10626;
wire n_11676;
wire n_1029;
wire n_2649;
wire n_6033;
wire n_6461;
wire n_10138;
wire n_1247;
wire n_6860;
wire n_9063;
wire n_522;
wire n_1568;
wire n_2919;
wire n_10364;
wire n_7322;
wire n_6060;
wire n_10532;
wire n_3108;
wire n_5788;
wire n_5983;
wire n_9895;
wire n_10288;
wire n_367;
wire n_6709;
wire n_11602;
wire n_13843;
wire n_2632;
wire n_11865;
wire n_12566;
wire n_5557;
wire n_12383;
wire n_6914;
wire n_8816;
wire n_4314;
wire n_8418;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_7287;
wire n_7789;
wire n_12035;
wire n_3239;
wire n_2631;
wire n_12212;
wire n_11427;
wire n_3311;
wire n_9110;
wire n_3516;
wire n_11613;
wire n_4442;
wire n_424;
wire n_10668;
wire n_4857;
wire n_8739;
wire n_9969;
wire n_11375;
wire n_8927;
wire n_10398;
wire n_1651;
wire n_3087;
wire n_6009;
wire n_7221;
wire n_5523;
wire n_11870;
wire n_12053;
wire n_2697;
wire n_13250;
wire n_4637;
wire n_1263;
wire n_1817;
wire n_8243;
wire n_3704;
wire n_8798;
wire n_13228;
wire n_7963;
wire n_13893;
wire n_6382;
wire n_8423;
wire n_13869;
wire n_14326;
wire n_9028;
wire n_670;
wire n_2677;
wire n_4296;
wire n_14699;
wire n_379;
wire n_138;
wire n_162;
wire n_13100;
wire n_9654;
wire n_10683;
wire n_14232;
wire n_2483;
wire n_10249;
wire n_7938;
wire n_5088;
wire n_6615;
wire n_9810;
wire n_441;
wire n_7294;
wire n_6192;
wire n_5773;
wire n_7414;
wire n_1032;
wire n_12852;
wire n_12123;
wire n_1592;
wire n_9701;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_9270;
wire n_11373;
wire n_11878;
wire n_3589;
wire n_6418;
wire n_1743;
wire n_8548;
wire n_9437;
wire n_8996;
wire n_13185;
wire n_207;
wire n_9483;
wire n_720;
wire n_6263;
wire n_1943;
wire n_14593;
wire n_6731;
wire n_8156;
wire n_5138;
wire n_8845;
wire n_4588;
wire n_6048;
wire n_13738;
wire n_10229;
wire n_7185;
wire n_194;
wire n_12268;
wire n_5149;
wire n_9256;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_10889;
wire n_11070;
wire n_6234;
wire n_4153;
wire n_8992;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_7141;
wire n_11107;
wire n_2373;
wire n_14116;
wire n_3881;
wire n_13195;
wire n_12298;
wire n_12930;
wire n_6224;
wire n_8510;
wire n_5089;
wire n_11394;
wire n_5775;
wire n_9854;
wire n_2099;
wire n_3759;
wire n_9737;
wire n_8961;
wire n_12890;
wire n_14551;
wire n_9964;
wire n_11154;
wire n_3323;
wire n_4643;
wire n_9719;
wire n_6142;
wire n_10826;
wire n_2617;
wire n_6119;
wire n_10358;
wire n_12301;
wire n_13886;
wire n_6619;
wire n_808;
wire n_2476;
wire n_11973;
wire n_13200;
wire n_2814;
wire n_4133;
wire n_11073;
wire n_13876;
wire n_2636;
wire n_1439;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_1665;
wire n_7092;
wire n_7233;
wire n_2122;
wire n_4543;
wire n_14442;
wire n_4337;
wire n_9679;
wire n_9669;
wire n_11186;
wire n_12382;
wire n_5082;
wire n_12996;
wire n_10835;
wire n_13095;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_10416;
wire n_3465;
wire n_12661;
wire n_8402;
wire n_8978;
wire n_14097;
wire n_7191;
wire n_2117;
wire n_14279;
wire n_6189;
wire n_1053;
wire n_5796;
wire n_13907;
wire n_9105;
wire n_13085;
wire n_14411;
wire n_9699;
wire n_11360;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_14304;
wire n_9673;
wire n_2194;
wire n_10860;
wire n_11823;
wire n_4780;
wire n_4640;
wire n_8685;
wire n_1828;
wire n_10997;
wire n_9240;
wire n_1304;
wire n_7202;
wire n_14033;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_7445;
wire n_5858;
wire n_9212;
wire n_13889;
wire n_5985;
wire n_8595;
wire n_10602;
wire n_604;
wire n_12088;
wire n_478;
wire n_11181;
wire n_9040;
wire n_1349;
wire n_9478;
wire n_10261;
wire n_10817;
wire n_12062;
wire n_12277;
wire n_14045;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_9742;
wire n_11806;
wire n_3477;
wire n_7868;
wire n_10124;
wire n_13386;
wire n_3370;
wire n_874;
wire n_7654;
wire n_3949;
wire n_2286;
wire n_8779;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_10132;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_8520;
wire n_4583;
wire n_14305;
wire n_8555;
wire n_12421;
wire n_10730;
wire n_9456;
wire n_6366;
wire n_1015;
wire n_11321;
wire n_1162;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_9146;
wire n_11702;
wire n_688;
wire n_7176;
wire n_14233;
wire n_636;
wire n_8565;
wire n_8334;
wire n_13605;
wire n_1490;
wire n_5552;
wire n_6074;
wire n_7547;
wire n_12133;
wire n_442;
wire n_11970;
wire n_3764;
wire n_1553;
wire n_13283;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_13596;
wire n_3025;
wire n_9573;
wire n_3051;
wire n_11286;
wire n_986;
wire n_1104;
wire n_2802;
wire n_8030;
wire n_8513;
wire n_14511;
wire n_887;
wire n_13746;
wire n_13327;
wire n_14550;
wire n_9379;
wire n_10948;
wire n_9219;
wire n_13534;
wire n_2125;
wire n_14056;
wire n_10927;
wire n_11496;
wire n_1156;
wire n_14151;
wire n_13149;
wire n_4974;
wire n_5123;
wire n_6689;
wire n_2861;
wire n_8245;
wire n_13727;
wire n_13992;
wire n_7942;
wire n_4344;
wire n_5242;
wire n_12186;
wire n_3130;
wire n_8753;
wire n_1188;
wire n_1498;
wire n_7527;
wire n_9706;
wire n_4856;
wire n_2618;
wire n_7948;
wire n_7096;
wire n_11863;
wire n_4216;
wire n_957;
wire n_1242;
wire n_9206;
wire n_2707;
wire n_14139;
wire n_8485;
wire n_6482;
wire n_5596;
wire n_10118;
wire n_8106;
wire n_2849;
wire n_1489;
wire n_8325;
wire n_2756;
wire n_3781;
wire n_14619;
wire n_2217;
wire n_10875;
wire n_4864;
wire n_11225;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_10731;
wire n_4313;
wire n_14071;
wire n_11355;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_9434;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_13198;
wire n_5536;
wire n_13097;
wire n_4798;
wire n_10350;
wire n_10654;
wire n_1500;
wire n_616;
wire n_7293;
wire n_9874;
wire n_11261;
wire n_11862;
wire n_13369;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_12579;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_10564;
wire n_3424;
wire n_12342;
wire n_13653;
wire n_3356;
wire n_14691;
wire n_11584;
wire n_9082;
wire n_7144;
wire n_12877;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_12256;
wire n_2516;
wire n_4991;
wire n_11893;
wire n_10262;
wire n_13360;
wire n_11500;
wire n_11044;
wire n_7316;
wire n_7508;
wire n_13785;
wire n_9596;
wire n_3070;
wire n_1005;
wire n_8677;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_11109;
wire n_12909;
wire n_13044;
wire n_3245;
wire n_12859;
wire n_10729;
wire n_2894;
wire n_9559;
wire n_9709;
wire n_10973;
wire n_2452;
wire n_4182;
wire n_8626;
wire n_12822;
wire n_2827;
wire n_7869;
wire n_13217;
wire n_3214;
wire n_13943;
wire n_10069;
wire n_10810;
wire n_12468;
wire n_9356;
wire n_8166;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_12267;
wire n_3710;
wire n_12170;
wire n_12426;
wire n_1844;
wire n_6943;
wire n_10791;
wire n_1957;
wire n_1953;
wire n_12900;
wire n_10553;
wire n_1219;
wire n_14555;
wire n_710;
wire n_6631;
wire n_5889;
wire n_12846;
wire n_8602;
wire n_9609;
wire n_7151;
wire n_10284;
wire n_3944;
wire n_7762;
wire n_13469;
wire n_13840;
wire n_13836;
wire n_5632;
wire n_12855;
wire n_11501;
wire n_4729;
wire n_8002;
wire n_6728;
wire n_13569;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_7472;
wire n_9342;
wire n_14229;
wire n_4800;
wire n_14425;
wire n_1373;
wire n_7075;
wire n_13076;
wire n_1540;
wire n_5427;
wire n_12234;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_6770;
wire n_14317;
wire n_5450;
wire n_7611;
wire n_11437;
wire n_7796;
wire n_6508;
wire n_14682;
wire n_832;
wire n_7989;
wire n_13082;
wire n_8047;
wire n_12120;
wire n_13320;
wire n_744;
wire n_2821;
wire n_3696;
wire n_9233;
wire n_10474;
wire n_7936;
wire n_10694;
wire n_215;
wire n_10529;
wire n_13117;
wire n_1331;
wire n_4781;
wire n_12042;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_14328;
wire n_5124;
wire n_655;
wire n_4237;
wire n_8751;
wire n_5297;
wire n_11722;
wire n_4828;
wire n_3333;
wire n_12568;
wire n_12149;
wire n_14444;
wire n_8800;
wire n_4652;
wire n_12278;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_7655;
wire n_10622;
wire n_1007;
wire n_9435;
wire n_1580;
wire n_3135;
wire n_13318;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_2448;
wire n_9557;
wire n_11639;
wire n_2211;
wire n_8955;
wire n_9551;
wire n_6365;
wire n_951;
wire n_8039;
wire n_8193;
wire n_12231;
wire n_12116;
wire n_9073;
wire n_13677;
wire n_7546;
wire n_8432;
wire n_14422;
wire n_5904;
wire n_11997;
wire n_6628;
wire n_5318;
wire n_8684;
wire n_10270;
wire n_2424;
wire n_5374;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_722;
wire n_13158;
wire n_7407;
wire n_12014;
wire n_13230;
wire n_9388;
wire n_3277;
wire n_10463;
wire n_9721;
wire n_11731;
wire n_14061;
wire n_4863;
wire n_10880;
wire n_11610;
wire n_12097;
wire n_14612;
wire n_12363;
wire n_13115;
wire n_13427;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_6328;
wire n_11498;
wire n_12008;
wire n_6929;
wire n_11509;
wire n_4859;
wire n_4568;
wire n_8628;
wire n_14401;
wire n_14034;
wire n_13559;
wire n_3617;
wire n_6012;
wire n_704;
wire n_2958;
wire n_7481;
wire n_11447;
wire n_1044;
wire n_1714;
wire n_4429;
wire n_5435;
wire n_6484;
wire n_11706;
wire n_3340;
wire n_5053;
wire n_7182;
wire n_11055;
wire n_14498;
wire n_10689;
wire n_9507;
wire n_5476;
wire n_5483;
wire n_12534;
wire n_9539;
wire n_8617;
wire n_14297;
wire n_14517;
wire n_7605;
wire n_8591;
wire n_8090;
wire n_1243;
wire n_9268;
wire n_5511;
wire n_9718;
wire n_8661;
wire n_13512;
wire n_10068;
wire n_3486;
wire n_6639;
wire n_11258;
wire n_358;
wire n_608;
wire n_9672;
wire n_12748;
wire n_11168;
wire n_9890;
wire n_12272;
wire n_9187;
wire n_2457;
wire n_9572;
wire n_12148;
wire n_2992;
wire n_10363;
wire n_6124;
wire n_12142;
wire n_12615;
wire n_13201;
wire n_9527;
wire n_317;
wire n_3197;
wire n_11234;
wire n_9949;
wire n_13388;
wire n_14484;
wire n_7423;
wire n_13674;
wire n_3256;
wire n_1878;
wire n_7375;
wire n_7076;
wire n_7689;
wire n_6344;
wire n_8189;
wire n_8811;
wire n_13858;
wire n_266;
wire n_9952;
wire n_11612;
wire n_7736;
wire n_6435;
wire n_13949;
wire n_10888;
wire n_12714;
wire n_13782;
wire n_14486;
wire n_3646;
wire n_14759;
wire n_5829;
wire n_2520;
wire n_14580;
wire n_7419;
wire n_811;
wire n_13612;
wire n_6600;
wire n_14087;
wire n_13681;
wire n_7010;
wire n_13700;
wire n_14421;
wire n_14193;
wire n_791;
wire n_10277;
wire n_5881;
wire n_9798;
wire n_3864;
wire n_4694;
wire n_11895;
wire n_8192;
wire n_9251;
wire n_1025;
wire n_4664;
wire n_6201;
wire n_10537;
wire n_14684;
wire n_3450;
wire n_14653;
wire n_8573;
wire n_14703;
wire n_687;
wire n_4633;
wire n_13770;
wire n_2026;
wire n_10807;
wire n_4050;
wire n_3173;
wire n_480;
wire n_14048;
wire n_13920;
wire n_7918;
wire n_642;
wire n_9546;
wire n_10331;
wire n_1406;
wire n_5073;
wire n_6555;
wire n_4306;
wire n_6360;
wire n_13130;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_9602;
wire n_9181;
wire n_12812;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_13377;
wire n_11455;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_474;
wire n_4098;
wire n_2691;
wire n_10981;
wire n_5894;
wire n_13750;
wire n_9635;
wire n_11868;
wire n_4511;
wire n_3422;
wire n_12189;
wire n_12639;
wire n_14063;
wire n_14343;
wire n_14521;
wire n_4675;
wire n_13701;
wire n_695;
wire n_11934;
wire n_13518;
wire n_2991;
wire n_5419;
wire n_8339;
wire n_14737;
wire n_386;
wire n_1596;
wire n_11969;
wire n_13668;
wire n_4289;
wire n_4972;
wire n_11571;
wire n_197;
wire n_2723;
wire n_1476;
wire n_7346;
wire n_9405;
wire n_6036;
wire n_2016;
wire n_3925;
wire n_12428;
wire n_12069;
wire n_14384;
wire n_4689;
wire n_5165;
wire n_8775;
wire n_678;
wire n_10780;
wire n_10158;
wire n_11481;
wire n_651;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_6102;
wire n_14276;
wire n_12057;
wire n_3780;
wire n_12050;
wire n_1657;
wire n_13587;
wire n_9726;
wire n_13488;
wire n_8804;
wire n_9577;
wire n_6650;
wire n_10024;
wire n_6573;
wire n_11774;
wire n_6904;
wire n_12214;
wire n_3753;
wire n_6329;
wire n_13805;
wire n_7385;
wire n_9802;
wire n_1488;
wire n_6244;
wire n_4846;
wire n_9250;
wire n_1330;
wire n_906;
wire n_9540;
wire n_13365;
wire n_13767;
wire n_13972;
wire n_14357;
wire n_6204;
wire n_12381;
wire n_10191;
wire n_2295;
wire n_5225;
wire n_283;
wire n_7295;
wire n_4076;
wire n_7824;
wire n_12157;
wire n_7148;
wire n_13938;
wire n_3142;
wire n_9171;
wire n_7169;
wire n_3129;
wire n_13443;
wire n_9350;
wire n_374;
wire n_3495;
wire n_3843;
wire n_11257;
wire n_12330;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_9441;
wire n_7600;
wire n_9124;
wire n_10675;
wire n_2386;
wire n_5826;
wire n_8697;
wire n_11598;
wire n_9626;
wire n_14011;
wire n_14645;
wire n_4822;
wire n_11327;
wire n_6946;
wire n_12926;
wire n_7947;
wire n_8645;
wire n_8820;
wire n_9408;
wire n_8146;
wire n_5931;
wire n_1829;
wire n_14712;
wire n_4635;
wire n_7847;
wire n_8154;
wire n_1450;
wire n_12824;
wire n_12392;
wire n_13094;
wire n_5532;
wire n_14545;
wire n_7311;
wire n_3740;
wire n_6804;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_14103;
wire n_6059;
wire n_1815;
wire n_7039;
wire n_8027;
wire n_7807;
wire n_1493;
wire n_2911;
wire n_515;
wire n_8063;
wire n_3313;
wire n_13798;
wire n_14677;
wire n_8406;
wire n_2354;
wire n_6427;
wire n_14474;
wire n_14459;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_12070;
wire n_3726;
wire n_8480;
wire n_11265;
wire n_14037;
wire n_11788;
wire n_14112;
wire n_9754;
wire n_10477;
wire n_4419;
wire n_14296;
wire n_11904;
wire n_8849;
wire n_13071;
wire n_5405;
wire n_9750;
wire n_10296;
wire n_7660;
wire n_13676;
wire n_13735;
wire n_14127;
wire n_1256;
wire n_5365;
wire n_9529;
wire n_3560;
wire n_3345;
wire n_9566;
wire n_11901;
wire n_10339;
wire n_12848;
wire n_5772;
wire n_6442;
wire n_10307;
wire n_8241;
wire n_140;
wire n_10606;
wire n_6188;
wire n_12161;
wire n_3421;
wire n_1448;
wire n_10066;
wire n_11755;
wire n_1009;
wire n_230;
wire n_3548;
wire n_4906;
wire n_11754;
wire n_6846;
wire n_13825;
wire n_10054;
wire n_4630;
wire n_8261;
wire n_10343;
wire n_6840;
wire n_142;
wire n_6645;
wire n_8535;
wire n_8348;
wire n_13985;
wire n_4829;
wire n_6749;
wire n_12238;
wire n_6915;
wire n_12956;
wire n_12320;
wire n_7831;
wire n_8138;
wire n_13342;
wire n_2612;
wire n_11413;
wire n_13953;
wire n_10652;
wire n_13040;
wire n_5259;
wire n_3236;
wire n_8702;
wire n_11601;
wire n_1995;
wire n_7455;
wire n_8273;
wire n_14250;
wire n_10944;
wire n_1397;
wire n_6247;
wire n_10367;
wire n_5921;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_11129;
wire n_11710;
wire n_833;
wire n_4966;
wire n_14602;
wire n_2250;
wire n_8235;
wire n_13685;
wire n_1117;
wire n_6104;
wire n_3321;
wire n_9940;
wire n_8294;
wire n_1303;
wire n_12476;
wire n_4188;
wire n_10016;
wire n_2001;
wire n_9036;
wire n_9165;
wire n_7509;
wire n_9283;
wire n_6205;
wire n_2506;
wire n_11010;
wire n_8349;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_10036;
wire n_9822;
wire n_2626;
wire n_9443;
wire n_9607;
wire n_7497;
wire n_10749;
wire n_7315;
wire n_10166;
wire n_8429;
wire n_13765;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_10419;
wire n_7887;
wire n_2804;
wire n_9298;
wire n_5884;
wire n_5006;
wire n_14200;
wire n_4882;
wire n_3206;
wire n_10006;
wire n_5728;
wire n_1035;
wire n_13334;
wire n_3475;
wire n_4878;
wire n_8486;
wire n_11240;
wire n_9052;
wire n_2070;
wire n_426;
wire n_6706;
wire n_13123;
wire n_12154;
wire n_7431;
wire n_8140;
wire n_398;
wire n_11734;
wire n_14450;
wire n_3842;
wire n_12645;
wire n_1367;
wire n_14477;
wire n_4202;
wire n_6909;
wire n_13933;
wire n_2044;
wire n_5679;
wire n_6487;
wire n_166;
wire n_8117;
wire n_12668;
wire n_3886;
wire n_10348;
wire n_13884;
wire n_825;
wire n_732;
wire n_2619;
wire n_7521;
wire n_10058;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_8129;
wire n_1291;
wire n_10355;
wire n_11156;
wire n_7253;
wire n_5208;
wire n_9535;
wire n_13511;
wire n_5113;
wire n_10304;
wire n_12928;
wire n_3987;
wire n_11955;
wire n_5205;
wire n_4249;
wire n_9943;
wire n_7569;
wire n_12538;
wire n_13745;
wire n_12151;
wire n_3160;
wire n_10966;
wire n_14697;
wire n_13112;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_13646;
wire n_12130;
wire n_14608;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_12409;
wire n_13031;
wire n_6551;
wire n_3386;
wire n_12350;
wire n_400;
wire n_7972;
wire n_8672;
wire n_13455;
wire n_7505;
wire n_13993;
wire n_3921;
wire n_282;
wire n_14280;
wire n_467;
wire n_2177;
wire n_13946;
wire n_6516;
wire n_14567;
wire n_2766;
wire n_10060;
wire n_7524;
wire n_13931;
wire n_4196;
wire n_1197;
wire n_11270;
wire n_8934;
wire n_11020;
wire n_7318;
wire n_2613;
wire n_9977;
wire n_10722;
wire n_7411;
wire n_13314;
wire n_7326;
wire n_13378;
wire n_5667;
wire n_168;
wire n_9555;
wire n_1517;
wire n_13618;
wire n_10957;
wire n_2647;
wire n_14277;
wire n_8847;
wire n_8005;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_11344;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_6500;
wire n_11303;
wire n_5027;
wire n_1048;
wire n_2343;
wire n_775;
wire n_12847;
wire n_667;
wire n_3380;
wire n_14340;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_9030;
wire n_869;
wire n_11216;
wire n_846;
wire n_1398;
wire n_1921;
wire n_8221;
wire n_13638;
wire n_7573;
wire n_6630;
wire n_5629;
wire n_5759;
wire n_10409;
wire n_2411;
wire n_13167;
wire n_4631;
wire n_8191;
wire n_6798;
wire n_13758;
wire n_5999;
wire n_1504;
wire n_9590;
wire n_2110;
wire n_14646;
wire n_11511;
wire n_7498;
wire n_7895;
wire n_6421;
wire n_10322;
wire n_11339;
wire n_11346;
wire n_11829;
wire n_12680;
wire n_5377;
wire n_6180;
wire n_12530;
wire n_11581;
wire n_8225;
wire n_3822;
wire n_889;
wire n_4355;
wire n_7453;
wire n_3818;
wire n_12163;
wire n_14131;
wire n_7932;
wire n_9651;
wire n_7890;
wire n_5599;
wire n_10825;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_9583;
wire n_9763;
wire n_9944;
wire n_10349;
wire n_13709;
wire n_13035;
wire n_1948;
wire n_6652;
wire n_9888;
wire n_7183;
wire n_10040;
wire n_810;
wire n_4278;
wire n_10636;
wire n_10844;
wire n_4710;
wire n_12738;
wire n_4155;
wire n_1959;
wire n_6275;
wire n_6403;
wire n_3497;
wire n_6395;
wire n_9862;
wire n_14622;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_4326;
wire n_9966;
wire n_2121;
wire n_10242;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_9936;
wire n_565;
wire n_3927;
wire n_6141;
wire n_8559;
wire n_11165;
wire n_2068;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_1194;
wire n_9617;
wire n_10727;
wire n_4060;
wire n_1647;
wire n_9341;
wire n_6194;
wire n_1454;
wire n_2459;
wire n_941;
wire n_8689;
wire n_11231;
wire n_3396;
wire n_9749;
wire n_5517;
wire n_9629;
wire n_13654;
wire n_5807;
wire n_11448;
wire n_12227;
wire n_5426;
wire n_6475;
wire n_12525;
wire n_10679;
wire n_4093;
wire n_11132;
wire n_452;
wire n_10524;
wire n_12282;
wire n_5693;
wire n_13426;
wire n_5695;
wire n_12932;
wire n_4123;
wire n_13799;
wire n_14207;
wire n_4294;
wire n_8330;
wire n_10011;
wire n_1521;
wire n_12037;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_10030;
wire n_6944;
wire n_11410;
wire n_14365;
wire n_4452;
wire n_284;
wire n_3887;
wire n_3195;
wire n_8304;
wire n_9349;
wire n_13480;
wire n_11267;
wire n_4722;
wire n_5587;
wire n_13780;
wire n_6318;
wire n_10119;
wire n_11348;
wire n_11940;
wire n_13613;
wire n_10845;
wire n_8163;
wire n_6805;
wire n_11947;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_5030;
wire n_7240;
wire n_8907;
wire n_409;
wire n_2963;
wire n_14227;
wire n_5674;
wire n_2561;
wire n_7499;
wire n_9423;
wire n_1056;
wire n_526;
wire n_5584;
wire n_674;
wire n_12424;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_6075;
wire n_10063;
wire n_12942;
wire n_6559;
wire n_4088;
wire n_9038;
wire n_8777;
wire n_11149;
wire n_2669;
wire n_8698;
wire n_10709;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_12236;
wire n_4366;
wire n_1584;
wire n_6248;
wire n_6541;
wire n_11436;
wire n_9034;
wire n_848;
wire n_5125;
wire n_4922;
wire n_11909;
wire n_12547;
wire n_13554;
wire n_6066;
wire n_6080;
wire n_14372;
wire n_629;
wire n_13421;
wire n_4733;
wire n_7927;
wire n_161;
wire n_8928;
wire n_13967;
wire n_1814;
wire n_13150;
wire n_13014;
wire n_7219;
wire n_2441;
wire n_10526;
wire n_11439;
wire n_8081;
wire n_12192;
wire n_4041;
wire n_12747;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_216;
wire n_11462;
wire n_6638;
wire n_6150;
wire n_14564;
wire n_7063;
wire n_7402;
wire n_9676;
wire n_6351;
wire n_4509;
wire n_4935;
wire n_2073;
wire n_7382;
wire n_8384;
wire n_10861;
wire n_4004;
wire n_5238;
wire n_750;
wire n_13795;
wire n_834;
wire n_8650;
wire n_14729;
wire n_3630;
wire n_1612;
wire n_11272;
wire n_800;
wire n_14044;
wire n_12989;
wire n_1910;
wire n_5906;
wire n_7767;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_11759;
wire n_10494;
wire n_14431;
wire n_2602;
wire n_11061;
wire n_10478;
wire n_5780;
wire n_724;
wire n_11653;
wire n_2931;
wire n_3433;
wire n_8284;
wire n_10534;
wire n_8374;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_13662;
wire n_13864;
wire n_5743;
wire n_6481;
wire n_10078;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_11478;
wire n_7510;
wire n_12273;
wire n_5633;
wire n_9041;
wire n_3786;
wire n_875;
wire n_9995;
wire n_12200;
wire n_6991;
wire n_10629;
wire n_13863;
wire n_2828;
wire n_6022;
wire n_7434;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_9035;
wire n_13926;
wire n_9011;
wire n_1715;
wire n_14240;
wire n_4204;
wire n_7691;
wire n_296;
wire n_3553;
wire n_5323;
wire n_7745;
wire n_11748;
wire n_14165;
wire n_9135;
wire n_6744;
wire n_3645;
wire n_9776;
wire n_793;
wire n_5705;
wire n_12660;
wire n_11867;
wire n_14192;
wire n_6927;
wire n_14678;
wire n_7335;
wire n_12400;
wire n_13072;
wire n_14708;
wire n_10472;
wire n_10695;
wire n_10286;
wire n_9413;
wire n_4996;
wire n_9107;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_7735;
wire n_8531;
wire n_6116;
wire n_9548;
wire n_8074;
wire n_14246;
wire n_494;
wire n_3550;
wire n_8780;
wire n_7956;
wire n_5510;
wire n_7651;
wire n_7495;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_9775;
wire n_13857;
wire n_12922;
wire n_1805;
wire n_13033;
wire n_8580;
wire n_4068;
wire n_5440;
wire n_12193;
wire n_9288;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_185;
wire n_5011;
wire n_6757;
wire n_7536;
wire n_1554;
wire n_3279;
wire n_12243;
wire n_5513;
wire n_10218;
wire n_5875;
wire n_14671;
wire n_8358;
wire n_972;
wire n_7734;
wire n_4262;
wire n_2923;
wire n_10441;
wire n_164;
wire n_2843;
wire n_3714;
wire n_9305;
wire n_9093;
wire n_184;
wire n_11764;
wire n_7671;
wire n_13696;
wire n_12950;
wire n_10043;
wire n_4832;
wire n_8033;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_13041;
wire n_5848;
wire n_1679;
wire n_5834;
wire n_14269;
wire n_7926;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_11882;
wire n_5784;
wire n_13418;
wire n_3125;
wire n_12250;
wire n_5128;
wire n_10628;
wire n_13498;
wire n_14290;
wire n_8643;
wire n_2356;
wire n_11787;
wire n_12403;
wire n_5618;
wire n_11539;
wire n_10440;
wire n_10134;
wire n_12904;
wire n_6495;
wire n_7528;
wire n_14669;
wire n_12444;
wire n_11163;
wire n_6209;
wire n_4672;
wire n_8094;
wire n_2564;
wire n_3558;
wire n_11695;
wire n_9425;
wire n_13489;
wire n_14520;
wire n_13373;
wire n_3034;
wire n_10317;
wire n_13739;
wire n_11730;
wire n_13101;
wire n_11916;
wire n_13723;
wire n_3502;
wire n_783;
wire n_13000;
wire n_13556;
wire n_4053;
wire n_11311;
wire n_1127;
wire n_14525;
wire n_7413;
wire n_14435;
wire n_7993;
wire n_11980;
wire n_7821;
wire n_160;
wire n_11151;
wire n_14238;
wire n_7620;
wire n_1008;
wire n_3963;
wire n_13153;
wire n_12837;
wire n_12356;
wire n_581;
wire n_3091;
wire n_13091;
wire n_13937;
wire n_13032;
wire n_6274;
wire n_1024;
wire n_176;
wire n_5157;
wire n_12764;
wire n_14654;
wire n_4496;
wire n_9347;
wire n_12269;
wire n_14556;
wire n_2518;
wire n_12079;
wire n_14687;
wire n_936;
wire n_13508;
wire n_10706;
wire n_4596;
wire n_5178;
wire n_9420;
wire n_13350;
wire n_13901;
wire n_12972;
wire n_3105;
wire n_6237;
wire n_13635;
wire n_1525;
wire n_4628;
wire n_6802;
wire n_13224;
wire n_7343;
wire n_8477;
wire n_5982;
wire n_1775;
wire n_908;
wire n_13306;
wire n_1036;
wire n_9344;
wire n_14657;
wire n_12438;
wire n_7109;
wire n_8028;
wire n_14245;
wire n_14254;
wire n_12125;
wire n_341;
wire n_4083;
wire n_1270;
wire n_12554;
wire n_10297;
wire n_1272;
wire n_549;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_7506;
wire n_3940;
wire n_9530;
wire n_10160;
wire n_11296;
wire n_6099;
wire n_10849;
wire n_3225;
wire n_10605;
wire n_6809;
wire n_13259;
wire n_8530;
wire n_14217;
wire n_10379;
wire n_9446;
wire n_3621;
wire n_5529;
wire n_244;
wire n_7561;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_11081;
wire n_8500;
wire n_13278;
wire n_6716;
wire n_8713;
wire n_12860;
wire n_3565;
wire n_7885;
wire n_14554;
wire n_8297;
wire n_14100;
wire n_6905;
wire n_8926;
wire n_9865;
wire n_8456;
wire n_7722;
wire n_5388;
wire n_7470;
wire n_11230;
wire n_5824;
wire n_8025;
wire n_10282;
wire n_5354;
wire n_2453;
wire n_11357;
wire n_7898;
wire n_3331;
wire n_11027;
wire n_13179;
wire n_1788;
wire n_10458;
wire n_12206;
wire n_11393;
wire n_6203;
wire n_12947;
wire n_2138;
wire n_6407;
wire n_14468;
wire n_3040;
wire n_4230;
wire n_11892;
wire n_6899;
wire n_7980;
wire n_7817;
wire n_6413;
wire n_445;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_7070;
wire n_9025;
wire n_2000;
wire n_5276;
wire n_11105;
wire n_4037;
wire n_9713;
wire n_11160;
wire n_13043;
wire n_3804;
wire n_14675;
wire n_4659;
wire n_13962;
wire n_8293;
wire n_3211;
wire n_7299;
wire n_917;
wire n_5196;
wire n_2440;
wire n_2096;
wire n_2556;
wire n_10382;
wire n_8029;
wire n_2215;
wire n_13468;
wire n_9314;
wire n_3847;
wire n_12270;
wire n_6960;
wire n_4073;
wire n_14235;
wire n_8880;
wire n_1261;
wire n_7249;
wire n_9660;
wire n_5763;
wire n_3633;
wire n_857;
wire n_13018;
wire n_363;
wire n_12739;
wire n_6061;
wire n_1235;
wire n_13831;
wire n_9769;
wire n_2584;
wire n_4001;
wire n_8471;
wire n_1462;
wire n_5701;
wire n_7002;
wire n_14529;
wire n_1064;
wire n_633;
wire n_1446;
wire n_12906;
wire n_12490;
wire n_9902;
wire n_1701;
wire n_6273;
wire n_14424;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_12751;
wire n_11397;
wire n_8726;
wire n_10640;
wire n_731;
wire n_8977;
wire n_1813;
wire n_315;
wire n_2997;
wire n_7018;
wire n_11897;
wire n_10522;
wire n_1573;
wire n_6746;
wire n_3258;
wire n_10691;
wire n_758;
wire n_12650;
wire n_10764;
wire n_10244;
wire n_10914;
wire n_13348;
wire n_3691;
wire n_2252;
wire n_8316;
wire n_6174;
wire n_10272;
wire n_6545;
wire n_7773;
wire n_6763;
wire n_14690;
wire n_1996;
wire n_1106;
wire n_13415;
wire n_2009;
wire n_5907;
wire n_784;
wire n_4339;
wire n_7297;
wire n_7730;
wire n_10980;
wire n_12279;
wire n_13265;
wire n_8134;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_9588;
wire n_2651;
wire n_753;
wire n_9410;
wire n_12242;
wire n_2733;
wire n_2445;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_8610;
wire n_4023;
wire n_10071;
wire n_4253;
wire n_7637;
wire n_2522;
wire n_3632;
wire n_12588;
wire n_309;
wire n_1344;
wire n_485;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_13382;
wire n_10176;
wire n_435;
wire n_9740;
wire n_1141;
wire n_3457;
wire n_6113;
wire n_14767;
wire n_5384;
wire n_6477;
wire n_7486;
wire n_840;
wire n_2324;
wire n_6575;
wire n_11719;
wire n_5283;
wire n_9910;
wire n_3454;
wire n_5961;
wire n_7544;
wire n_2139;
wire n_7613;
wire n_9061;
wire n_7995;
wire n_9941;
wire n_8113;
wire n_9579;
wire n_2521;
wire n_5686;
wire n_10254;
wire n_6391;
wire n_2740;
wire n_14446;
wire n_1991;
wire n_8724;
wire n_14121;
wire n_10332;
wire n_7140;
wire n_12775;
wire n_614;
wire n_12173;
wire n_4066;
wire n_10938;
wire n_10257;
wire n_9668;
wire n_6252;
wire n_6426;
wire n_14031;
wire n_4681;
wire n_11956;
wire n_12167;
wire n_8253;
wire n_9258;
wire n_9228;
wire n_3303;
wire n_13461;
wire n_7910;
wire n_6592;
wire n_4414;
wire n_10214;
wire n_11874;
wire n_2541;
wire n_5094;
wire n_10195;
wire n_3232;
wire n_13979;
wire n_1113;
wire n_9598;
wire n_10354;
wire n_248;
wire n_7741;
wire n_12060;
wire n_3768;
wire n_4295;
wire n_10436;
wire n_1615;
wire n_11450;
wire n_4100;
wire n_228;
wire n_11723;
wire n_6668;
wire n_9311;
wire n_11982;
wire n_1265;
wire n_14062;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_11822;
wire n_12179;
wire n_14448;
wire n_11522;
wire n_4087;
wire n_8232;
wire n_12842;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_8803;
wire n_10866;
wire n_1673;
wire n_4473;
wire n_14715;
wire n_4619;
wire n_12499;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_7679;
wire n_3018;
wire n_8818;
wire n_12693;
wire n_10811;
wire n_7698;
wire n_1875;
wire n_10073;
wire n_6962;
wire n_14187;
wire n_2429;
wire n_6779;
wire n_9608;
wire n_5286;
wire n_10164;
wire n_4449;
wire n_14779;
wire n_13172;
wire n_3285;
wire n_4607;
wire n_10205;
wire n_1039;
wire n_5676;
wire n_14716;
wire n_5949;
wire n_5040;
wire n_10515;
wire n_12326;
wire n_1150;
wire n_7800;
wire n_6901;
wire n_4266;
wire n_6336;
wire n_13713;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_7835;
wire n_1136;
wire n_12542;
wire n_13650;
wire n_458;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_11499;
wire n_3628;
wire n_14390;
wire n_9818;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_11034;
wire n_7415;
wire n_14747;
wire n_8823;
wire n_5399;
wire n_8536;
wire n_9433;
wire n_14004;
wire n_11746;
wire n_658;
wire n_11698;
wire n_362;
wire n_8795;
wire n_2846;
wire n_3371;
wire n_10430;
wire n_12934;
wire n_10338;
wire n_11560;
wire n_9599;
wire n_8674;
wire n_9186;
wire n_14054;
wire n_4918;
wire n_13941;
wire n_8016;
wire n_5856;
wire n_3872;
wire n_5760;
wire n_12483;
wire n_7747;
wire n_9935;
wire n_14263;
wire n_12404;
wire n_12258;
wire n_4415;
wire n_5110;
wire n_8966;
wire n_11871;
wire n_14694;
wire n_1964;
wire n_3659;
wire n_7552;
wire n_3928;
wire n_10018;
wire n_9537;
wire n_10500;
wire n_1777;
wire n_9552;
wire n_9421;
wire n_3366;
wire n_6998;
wire n_7395;
wire n_13209;
wire n_5844;
wire n_10359;
wire n_6298;
wire n_8132;
wire n_7650;
wire n_3441;
wire n_199;
wire n_3020;
wire n_12823;
wire n_4146;
wire n_4947;
wire n_7535;
wire n_14775;
wire n_708;
wire n_6609;
wire n_10548;
wire n_2545;
wire n_2513;
wire n_7635;
wire n_4408;
wire n_12905;
wire n_10291;
wire n_2115;
wire n_8567;
wire n_8259;
wire n_2017;
wire n_10667;
wire n_1810;
wire n_12274;
wire n_12849;
wire n_1347;
wire n_11167;
wire n_11297;
wire n_4976;
wire n_9473;
wire n_860;
wire n_6525;
wire n_10208;
wire n_11183;
wire n_3555;
wire n_9469;
wire n_11285;
wire n_5938;
wire n_14270;
wire n_7274;
wire n_3534;
wire n_450;
wire n_11740;
wire n_8578;
wire n_10757;
wire n_4548;
wire n_7819;
wire n_8495;
wire n_14679;
wire n_2670;
wire n_13975;
wire n_6494;
wire n_3556;
wire n_896;
wire n_4574;
wire n_8160;
wire n_8980;
wire n_2644;
wire n_10631;
wire n_6132;
wire n_10864;
wire n_11136;
wire n_4557;
wire n_3071;
wire n_11434;
wire n_8336;
wire n_11133;
wire n_1698;
wire n_14710;
wire n_14781;
wire n_13711;
wire n_1337;
wire n_774;
wire n_2148;
wire n_5548;
wire n_7788;
wire n_6974;
wire n_13477;
wire n_1168;
wire n_10748;
wire n_14783;
wire n_4663;
wire n_219;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_9909;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_656;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_12303;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_12002;
wire n_8600;
wire n_8229;
wire n_12442;
wire n_415;
wire n_4686;
wire n_9751;
wire n_9236;
wire n_2384;
wire n_10751;
wire n_14649;
wire n_7794;
wire n_1705;
wire n_13579;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_10434;
wire n_9369;
wire n_3149;
wire n_3934;
wire n_13634;
wire n_4338;
wire n_13987;
wire n_12597;
wire n_5917;
wire n_9757;
wire n_12419;
wire n_6965;
wire n_11886;
wire n_2058;
wire n_3231;
wire n_14210;
wire n_8761;
wire n_1846;
wire n_14316;
wire n_7630;
wire n_11804;
wire n_13262;
wire n_4161;
wire n_304;
wire n_14673;
wire n_9076;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6951;
wire n_6963;
wire n_1581;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_375;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_5355;
wire n_9729;
wire n_11531;
wire n_12943;
wire n_13543;
wire n_6284;
wire n_998;
wire n_3592;
wire n_12039;
wire n_10663;
wire n_14393;
wire n_5321;
wire n_14144;
wire n_7454;
wire n_2536;
wire n_10263;
wire n_12295;
wire n_1604;
wire n_3399;
wire n_8473;
wire n_9366;
wire n_4772;
wire n_11883;
wire n_6931;
wire n_6521;
wire n_8351;
wire n_5915;
wire n_7276;
wire n_174;
wire n_11792;
wire n_6379;
wire n_9647;
wire n_12410;
wire n_1368;
wire n_963;
wire n_7085;
wire n_6306;
wire n_12938;
wire n_4120;
wire n_925;
wire n_7753;
wire n_12891;
wire n_13493;
wire n_12304;
wire n_6834;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_1115;
wire n_8948;
wire n_13166;
wire n_14760;
wire n_13541;
wire n_1339;
wire n_12572;
wire n_10318;
wire n_13551;
wire n_1051;
wire n_14356;
wire n_5116;
wire n_3771;
wire n_10740;
wire n_7225;
wire n_719;
wire n_11634;
wire n_7541;
wire n_3158;
wire n_11039;
wire n_3221;
wire n_10062;
wire n_2316;
wire n_10128;
wire n_7913;
wire n_8020;
wire n_7946;
wire n_8944;
wire n_1010;
wire n_2830;
wire n_10717;
wire n_11965;
wire n_5500;
wire n_13890;
wire n_9275;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_9520;
wire n_6949;
wire n_6471;
wire n_11477;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_9493;
wire n_5621;
wire n_6760;
wire n_2940;
wire n_548;
wire n_3427;
wire n_8875;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_9102;
wire n_5966;
wire n_14128;
wire n_5515;
wire n_11588;
wire n_11818;
wire n_6589;
wire n_11592;
wire n_3083;
wire n_4570;
wire n_10721;
wire n_7014;
wire n_10945;
wire n_12290;
wire n_9801;
wire n_11742;
wire n_2491;
wire n_13902;
wire n_12718;
wire n_7920;
wire n_11312;
wire n_1931;
wire n_5559;
wire n_8649;
wire n_2259;
wire n_5337;
wire n_849;
wire n_11235;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_14185;
wire n_1820;
wire n_7841;
wire n_9424;
wire n_10013;
wire n_7324;
wire n_7160;
wire n_9333;
wire n_8205;
wire n_11505;
wire n_12469;
wire n_6046;
wire n_11673;
wire n_7054;
wire n_1233;
wire n_4493;
wire n_8975;
wire n_6055;
wire n_7161;
wire n_9004;
wire n_1808;
wire n_6364;
wire n_8919;
wire n_6091;
wire n_6348;
wire n_9987;
wire n_1635;
wire n_8440;
wire n_11555;
wire n_1704;
wire n_13917;
wire n_4896;
wire n_8041;
wire n_4851;
wire n_6848;
wire n_2479;
wire n_9860;
wire n_10565;
wire n_886;
wire n_14327;
wire n_7837;
wire n_359;
wire n_9670;
wire n_13548;
wire n_6788;
wire n_1308;
wire n_13903;
wire n_11241;
wire n_6144;
wire n_10389;
wire n_1451;
wire n_1487;
wire n_675;
wire n_9200;
wire n_5528;
wire n_7806;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_12336;
wire n_1938;
wire n_13080;
wire n_9417;
wire n_11059;
wire n_6896;
wire n_2484;
wire n_5753;
wire n_8076;
wire n_5358;
wire n_12248;
wire n_12931;
wire n_1469;
wire n_14047;
wire n_11066;
wire n_4901;
wire n_3480;
wire n_8757;
wire n_1355;
wire n_10020;
wire n_7201;
wire n_13408;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_9386;
wire n_12713;
wire n_8897;
wire n_12810;
wire n_7676;
wire n_8177;
wire n_11683;
wire n_13733;
wire n_2334;
wire n_14311;
wire n_5467;
wire n_7241;
wire n_1169;
wire n_789;
wire n_3181;
wire n_14147;
wire n_5493;
wire n_9207;
wire n_13592;
wire n_1916;
wire n_6285;
wire n_10356;
wire n_12717;
wire n_610;
wire n_13915;
wire n_7644;
wire n_9276;
wire n_4602;
wire n_1713;
wire n_7816;
wire n_8829;
wire n_12119;
wire n_14186;
wire n_1436;
wire n_2818;
wire n_14149;
wire n_4900;
wire n_10110;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_11275;
wire n_7430;
wire n_14540;
wire n_13589;
wire n_3487;
wire n_3668;
wire n_11329;
wire n_2011;
wire n_8638;
wire n_1515;
wire n_817;
wire n_14272;
wire n_13189;
wire n_13260;
wire n_5901;
wire n_9980;
wire n_1566;
wire n_2837;
wire n_11923;
wire n_717;
wire n_952;
wire n_11718;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_7724;
wire n_5360;
wire n_10501;
wire n_7269;
wire n_12003;
wire n_7047;
wire n_2671;
wire n_12292;
wire n_2702;
wire n_10908;
wire n_9176;
wire n_6937;
wire n_4363;
wire n_12405;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_214;
wire n_9728;
wire n_11809;
wire n_4103;
wire n_10777;
wire n_2529;
wire n_8101;
wire n_2374;
wire n_13712;
wire n_5439;
wire n_8687;
wire n_6115;
wire n_1225;
wire n_3154;
wire n_9866;
wire n_137;
wire n_14685;
wire n_8721;
wire n_1366;
wire n_8749;
wire n_12780;
wire n_13349;
wire n_9465;
wire n_13277;
wire n_3938;
wire n_11975;
wire n_8937;
wire n_2278;
wire n_6272;
wire n_7067;
wire n_12087;
wire n_13233;
wire n_13808;
wire n_14478;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_5250;
wire n_4842;
wire n_12662;
wire n_10965;
wire n_4416;
wire n_7879;
wire n_8730;
wire n_11441;
wire n_12416;
wire n_9702;
wire n_10998;
wire n_13503;
wire n_6607;
wire n_12854;
wire n_4439;
wire n_520;
wire n_870;
wire n_4985;
wire n_12936;
wire n_9000;
wire n_13056;
wire n_3382;
wire n_13300;
wire n_11743;
wire n_12765;
wire n_3930;
wire n_3808;
wire n_13087;
wire n_9610;
wire n_5471;
wire n_2248;
wire n_7117;
wire n_813;
wire n_10082;
wire n_8503;
wire n_10870;
wire n_12796;
wire n_4660;
wire n_11914;
wire n_3081;
wire n_6446;
wire n_10756;
wire n_5497;
wire n_9139;
wire n_13287;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_12028;
wire n_8315;
wire n_11175;
wire n_1961;
wire n_10411;
wire n_1535;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_871;
wire n_6807;
wire n_2844;
wire n_11753;
wire n_8197;
wire n_13726;
wire n_11790;
wire n_402;
wire n_1979;
wire n_9407;
wire n_6616;
wire n_6719;
wire n_12294;
wire n_14621;
wire n_10423;
wire n_829;
wire n_4814;
wire n_8019;
wire n_8801;
wire n_12190;
wire n_14396;
wire n_339;
wire n_6178;
wire n_11249;
wire n_8707;
wire n_6677;
wire n_11791;
wire n_2221;
wire n_12786;
wire n_7875;
wire n_5502;
wire n_8962;
wire n_13665;
wire n_8931;
wire n_8248;
wire n_14177;
wire n_1283;
wire n_7550;
wire n_14533;
wire n_8554;
wire n_2317;
wire n_2838;
wire n_13242;
wire n_1736;
wire n_11879;
wire n_13900;
wire n_10782;
wire n_13837;
wire n_2200;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_12386;
wire n_13121;
wire n_13679;
wire n_13680;
wire n_9357;
wire n_2442;
wire n_9477;
wire n_11911;
wire n_13734;
wire n_14591;
wire n_7238;
wire n_6862;
wire n_8501;
wire n_3657;
wire n_5706;
wire n_11842;
wire n_12746;
wire n_14023;
wire n_2634;
wire n_13047;
wire n_11320;
wire n_11304;
wire n_2746;
wire n_7292;
wire n_242;
wire n_645;
wire n_13146;
wire n_7804;
wire n_10251;
wire n_12128;
wire n_11776;
wire n_14544;
wire n_11471;
wire n_5098;
wire n_13475;
wire n_721;
wire n_1084;
wire n_6000;
wire n_6774;
wire n_9289;
wire n_11794;
wire n_6443;
wire n_9828;
wire n_1276;
wire n_8263;
wire n_5145;
wire n_6072;
wire n_13236;
wire n_2878;
wire n_7248;
wire n_10737;
wire n_3830;
wire n_10475;
wire n_3252;
wire n_6647;
wire n_11198;
wire n_8040;
wire n_13336;
wire n_5466;
wire n_14465;
wire n_1528;
wire n_7239;
wire n_9797;
wire n_6941;
wire n_6552;
wire n_7826;
wire n_10665;
wire n_9981;
wire n_3315;
wire n_6094;
wire n_14482;
wire n_3523;
wire n_12113;
wire n_8102;
wire n_3999;
wire n_14440;
wire n_10541;
wire n_13393;
wire n_14765;
wire n_9793;
wire n_518;
wire n_11419;
wire n_14214;
wire n_13202;
wire n_8196;
wire n_11171;
wire n_12017;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_8822;
wire n_7112;
wire n_3474;
wire n_5738;
wire n_14483;
wire n_9514;
wire n_2458;
wire n_7971;
wire n_12139;
wire n_8885;
wire n_11564;
wire n_5592;
wire n_11078;
wire n_5620;
wire n_12802;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_10633;
wire n_12592;
wire n_4782;
wire n_9825;
wire n_1539;
wire n_2859;
wire n_10573;
wire n_5216;
wire n_3412;
wire n_11218;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_8474;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_10258;
wire n_6886;
wire n_7078;
wire n_1636;
wire n_4597;
wire n_12791;
wire n_9501;
wire n_12352;
wire n_13811;
wire n_12296;
wire n_11459;
wire n_9043;
wire n_8152;
wire n_12491;
wire n_11998;
wire n_8269;
wire n_4546;
wire n_11775;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_11288;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_12454;
wire n_10042;
wire n_12162;
wire n_10570;
wire n_13151;
wire n_3073;
wire n_6531;
wire n_9481;
wire n_3571;
wire n_11768;
wire n_238;
wire n_4576;
wire n_7577;
wire n_12992;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_11456;
wire n_14706;
wire n_11708;
wire n_14330;
wire n_12960;
wire n_8144;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_11662;
wire n_13617;
wire n_7513;
wire n_10098;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_7812;
wire n_5330;
wire n_9351;
wire n_9766;
wire n_13935;
wire n_13930;
wire n_6935;
wire n_1560;
wire n_2899;
wire n_10106;
wire n_6984;
wire n_12046;
wire n_8058;
wire n_11877;
wire n_6778;
wire n_8909;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_12074;
wire n_14380;
wire n_3817;
wire n_6345;
wire n_9242;
wire n_10754;
wire n_6386;
wire n_2722;
wire n_3728;
wire n_6596;
wire n_12749;
wire n_612;
wire n_333;
wire n_14630;
wire n_5107;
wire n_7165;
wire n_512;
wire n_9777;
wire n_4680;
wire n_5067;
wire n_11932;
wire n_11821;
wire n_12485;
wire n_14464;
wire n_9522;
wire n_14560;
wire n_6830;
wire n_1012;
wire n_2685;
wire n_2061;
wire n_9748;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_12488;
wire n_14028;
wire n_12252;
wire n_10851;
wire n_12090;
wire n_9005;
wire n_11395;
wire n_2788;
wire n_10387;
wire n_9666;
wire n_6291;
wire n_6642;
wire n_6510;
wire n_1443;
wire n_10615;
wire n_5264;
wire n_14081;
wire n_14281;
wire n_2595;
wire n_10790;
wire n_1465;
wire n_3084;
wire n_10028;
wire n_705;
wire n_10555;
wire n_12896;
wire n_7667;
wire n_6781;
wire n_4593;
wire n_11532;
wire n_8024;
wire n_7123;
wire n_14670;
wire n_4562;
wire n_3860;
wire n_10222;
wire n_2909;
wire n_461;
wire n_3554;
wire n_12868;
wire n_6509;
wire n_10671;
wire n_2717;
wire n_6376;
wire n_1391;
wire n_8107;
wire n_9605;
wire n_2981;
wire n_10498;
wire n_225;
wire n_13959;
wire n_9947;
wire n_1006;
wire n_546;
wire n_9930;
wire n_14755;
wire n_13292;
wire n_4995;
wire n_1159;
wire n_6514;
wire n_10420;
wire n_4498;
wire n_5873;
wire n_772;
wire n_6741;
wire n_10083;
wire n_1245;
wire n_10520;
wire n_6434;
wire n_9662;
wire n_5741;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_9768;
wire n_1675;
wire n_2466;
wire n_6593;
wire n_676;
wire n_7827;
wire n_3758;
wire n_7631;
wire n_12583;
wire n_8748;
wire n_14420;
wire n_8452;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_10255;
wire n_8742;
wire n_3777;
wire n_8393;
wire n_9835;
wire n_11117;
wire n_11494;
wire n_1872;
wire n_9656;
wire n_1585;
wire n_11643;
wire n_14613;
wire n_3767;
wire n_12462;
wire n_12618;
wire n_14090;
wire n_14604;
wire n_6056;
wire n_9475;
wire n_5866;
wire n_5926;
wire n_212;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_14347;
wire n_2216;
wire n_11475;
wire n_8122;
wire n_11004;
wire n_9724;
wire n_2426;
wire n_652;
wire n_6947;
wire n_8403;
wire n_8912;
wire n_10612;
wire n_4850;
wire n_10007;
wire n_9154;
wire n_12127;
wire n_13651;
wire n_1260;
wire n_3716;
wire n_11223;
wire n_11570;
wire n_7157;
wire n_2926;
wire n_10937;
wire n_4937;
wire n_798;
wire n_8740;
wire n_10493;
wire n_13631;
wire n_5574;
wire n_13264;
wire n_13678;
wire n_8310;
wire n_3391;
wire n_5877;
wire n_14406;
wire n_912;
wire n_10104;
wire n_6375;
wire n_460;
wire n_11212;
wire n_10552;
wire n_7781;
wire n_13294;
wire n_4786;
wire n_6042;
wire n_14746;
wire n_8238;
wire n_5203;
wire n_7908;
wire n_10295;
wire n_8296;
wire n_10954;
wire n_7091;
wire n_9833;
wire n_9788;
wire n_4354;
wire n_9589;
wire n_4235;
wire n_6429;
wire n_3159;
wire n_6315;
wire n_7855;
wire n_14590;
wire n_8850;
wire n_9861;
wire n_2855;
wire n_794;
wire n_2848;
wire n_7886;
wire n_14740;
wire n_7675;
wire n_11122;
wire n_6775;
wire n_8943;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_8993;
wire n_11159;
wire n_12329;
wire n_9205;
wire n_11631;
wire n_9418;
wire n_9946;
wire n_288;
wire n_10376;
wire n_1292;
wire n_7774;
wire n_8634;
wire n_12611;
wire n_11715;
wire n_13625;
wire n_8831;
wire n_6970;
wire n_13034;
wire n_1026;
wire n_9979;
wire n_12205;
wire n_13122;
wire n_6948;
wire n_3460;
wire n_14324;
wire n_13210;
wire n_1610;
wire n_5155;
wire n_8676;
wire n_14337;
wire n_2202;
wire n_11889;
wire n_14509;
wire n_306;
wire n_3530;
wire n_2952;
wire n_6133;
wire n_10341;
wire n_2693;
wire n_7409;
wire n_10087;
wire n_5408;
wire n_11278;
wire n_12606;
wire n_6920;
wire n_14692;
wire n_8758;
wire n_11671;
wire n_5812;
wire n_9973;
wire n_5540;
wire n_11782;
wire n_7381;
wire n_5804;
wire n_9007;
wire n_8544;
wire n_3240;
wire n_7999;
wire n_5066;
wire n_14253;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_967;
wire n_9020;
wire n_10027;
wire n_9260;
wire n_5130;
wire n_14212;
wire n_4175;
wire n_10154;
wire n_6241;
wire n_13597;
wire n_9619;
wire n_14392;
wire n_13510;
wire n_1079;
wire n_5200;
wire n_9235;
wire n_3393;
wire n_10161;
wire n_13003;
wire n_8652;
wire n_9112;
wire n_12365;
wire n_2836;
wire n_12423;
wire n_7873;
wire n_12843;
wire n_2864;
wire n_4456;
wire n_11372;
wire n_1717;
wire n_9691;
wire n_5992;
wire n_8646;
wire n_13573;
wire n_2172;
wire n_2601;
wire n_12518;
wire n_12861;
wire n_2365;
wire n_1880;
wire n_9133;
wire n_5684;
wire n_1399;
wire n_13708;
wire n_7228;
wire n_5981;
wire n_7784;
wire n_9752;
wire n_1855;
wire n_6632;
wire n_2333;
wire n_8999;
wire n_3629;
wire n_4948;
wire n_10902;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_7713;
wire n_6623;
wire n_9395;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_1226;
wire n_2224;
wire n_6933;
wire n_1970;
wire n_10294;
wire n_3724;
wire n_9353;
wire n_11155;
wire n_3287;
wire n_11714;
wire n_12293;
wire n_2167;
wire n_13947;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_8031;
wire n_3257;
wire n_11590;
wire n_9804;
wire n_12450;
wire n_5737;
wire n_9125;
wire n_8015;
wire n_8412;
wire n_425;
wire n_3730;
wire n_8439;
wire n_8575;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_13648;
wire n_5097;
wire n_10323;
wire n_2695;
wire n_7084;
wire n_11976;
wire n_13274;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_9397;
wire n_10969;
wire n_8499;
wire n_13015;
wire n_13472;
wire n_13322;
wire n_13870;
wire n_7640;
wire n_12000;
wire n_6390;
wire n_2302;
wire n_6799;
wire n_8772;
wire n_10806;
wire n_9767;
wire n_12903;
wire n_3014;
wire n_7912;
wire n_2294;
wire n_6278;
wire n_11430;
wire n_2274;
wire n_7195;
wire n_12309;
wire n_5640;
wire n_3342;
wire n_13401;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_8557;
wire n_13891;
wire n_3796;
wire n_9384;
wire n_3884;
wire n_4492;
wire n_13850;
wire n_3625;
wire n_13835;
wire n_5550;
wire n_397;
wire n_3375;
wire n_2768;
wire n_351;
wire n_10666;
wire n_12895;
wire n_155;
wire n_3760;
wire n_5661;
wire n_7641;
wire n_4975;
wire n_11638;
wire n_3515;
wire n_2363;
wire n_12687;
wire n_12023;
wire n_14460;
wire n_5306;
wire n_5905;
wire n_13908;
wire n_8815;
wire n_7949;
wire n_6112;
wire n_11659;
wire n_2728;
wire n_9906;
wire n_2025;
wire n_8679;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_11948;
wire n_4022;
wire n_7115;
wire n_1020;
wire n_9310;
wire n_11843;
wire n_10659;
wire n_11689;
wire n_7764;
wire n_8446;
wire n_9163;
wire n_172;
wire n_11535;
wire n_2495;
wire n_12022;
wire n_1058;
wire n_12624;
wire n_4336;
wire n_11808;
wire n_8789;
wire n_8128;
wire n_7520;
wire n_5314;
wire n_9322;
wire n_12719;
wire n_7616;
wire n_14493;
wire n_10793;
wire n_14491;
wire n_8359;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_1279;
wire n_6271;
wire n_11108;
wire n_9377;
wire n_7235;
wire n_2511;
wire n_564;
wire n_6572;
wire n_9224;
wire n_10211;
wire n_10837;
wire n_3981;
wire n_14381;
wire n_12664;
wire n_13020;
wire n_11577;
wire n_7271;
wire n_9055;
wire n_13749;
wire n_13311;
wire n_2681;
wire n_7222;
wire n_8678;
wire n_9971;
wire n_1689;
wire n_8605;
wire n_2535;
wire n_12981;
wire n_13945;
wire n_1255;
wire n_3031;
wire n_345;
wire n_10976;
wire n_9624;
wire n_14766;
wire n_6930;
wire n_10045;
wire n_14172;
wire n_2335;
wire n_10289;
wire n_5482;
wire n_9145;
wire n_12716;
wire n_10232;
wire n_13079;
wire n_11098;
wire n_3215;
wire n_8443;
wire n_8525;
wire n_12166;
wire n_12507;
wire n_1401;
wire n_3138;
wire n_8312;
wire n_10819;
wire n_776;
wire n_2860;
wire n_8901;
wire n_2041;
wire n_13786;
wire n_1933;
wire n_13645;
wire n_6584;
wire n_4494;
wire n_9887;
wire n_12044;
wire n_6387;
wire n_466;
wire n_9373;
wire n_4201;
wire n_346;
wire n_14374;
wire n_6470;
wire n_7206;
wire n_8869;
wire n_552;
wire n_11279;
wire n_11729;
wire n_14012;
wire n_9770;
wire n_11514;
wire n_5287;
wire n_8272;
wire n_4719;
wire n_5651;
wire n_264;
wire n_3577;
wire n_6625;
wire n_14569;
wire n_4074;
wire n_7383;
wire n_12430;
wire n_3994;
wire n_4636;
wire n_11606;
wire n_4983;
wire n_3185;
wire n_6826;
wire n_10306;
wire n_12902;
wire n_12257;
wire n_1217;
wire n_11727;
wire n_13299;
wire n_10103;
wire n_14664;
wire n_11337;
wire n_327;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_10183;
wire n_1231;
wire n_12839;
wire n_13693;
wire n_5623;
wire n_11778;
wire n_12925;
wire n_11658;
wire n_10710;
wire n_8870;
wire n_9753;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_10931;
wire n_9468;
wire n_11433;
wire n_8178;
wire n_5524;
wire n_7854;
wire n_9517;
wire n_926;
wire n_9544;
wire n_2296;
wire n_5735;
wire n_7959;
wire n_14338;
wire n_14728;
wire n_8234;
wire n_6363;
wire n_13434;
wire n_6588;
wire n_11369;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_7897;
wire n_12759;
wire n_11720;
wire n_14418;
wire n_186;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_13500;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_1501;
wire n_8488;
wire n_11840;
wire n_2241;
wire n_6865;
wire n_11284;
wire n_12553;
wire n_13113;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_9774;
wire n_2531;
wire n_7132;
wire n_12016;
wire n_11987;
wire n_12496;
wire n_1570;
wire n_7533;
wire n_9586;
wire n_11052;
wire n_10670;
wire n_13655;
wire n_10150;
wire n_3377;
wire n_6722;
wire n_9780;
wire n_1518;
wire n_13476;
wire n_11177;
wire n_6420;
wire n_10004;
wire n_4907;
wire n_11169;
wire n_3961;
wire n_5153;
wire n_7766;
wire n_855;
wire n_8862;
wire n_13229;
wire n_2059;
wire n_14092;
wire n_8184;
wire n_13950;
wire n_4713;
wire n_6911;
wire n_5787;
wire n_11221;
wire n_14219;
wire n_13344;
wire n_10353;
wire n_10151;
wire n_1287;
wire n_11095;
wire n_10187;
wire n_1611;
wire n_10171;
wire n_11211;
wire n_7129;
wire n_12138;
wire n_7080;
wire n_3374;
wire n_4870;
wire n_7776;
wire n_6981;
wire n_4818;
wire n_8001;
wire n_10406;
wire n_8695;
wire n_12230;
wire n_12521;
wire n_11236;
wire n_11931;
wire n_7436;
wire n_8767;
wire n_11036;
wire n_12562;
wire n_8571;
wire n_7020;
wire n_11600;
wire n_5935;
wire n_8064;
wire n_14117;
wire n_14588;
wire n_6696;
wire n_13721;
wire n_4916;
wire n_8472;
wire n_13302;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_529;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_12217;
wire n_13535;
wire n_14261;
wire n_3508;
wire n_6300;
wire n_13704;
wire n_6653;
wire n_6372;
wire n_13969;
wire n_4129;
wire n_7120;
wire n_11114;
wire n_10479;
wire n_7978;
wire n_10033;
wire n_5488;
wire n_9099;
wire n_1105;
wire n_6900;
wire n_10034;
wire n_5727;
wire n_11336;
wire n_3599;
wire n_6660;
wire n_8787;
wire n_11009;
wire n_9543;
wire n_8131;
wire n_5988;
wire n_6424;
wire n_10696;
wire n_14633;
wire n_11480;
wire n_5646;
wire n_14538;
wire n_7448;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_6787;
wire n_7694;
wire n_8771;
wire n_9245;
wire n_5832;
wire n_13269;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_983;
wire n_7142;
wire n_10360;
wire n_6423;
wire n_6526;
wire n_699;
wire n_3542;
wire n_301;
wire n_3263;
wire n_8150;
wire n_5891;
wire n_2523;
wire n_1945;
wire n_9168;
wire n_11423;
wire n_12691;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_9074;
wire n_12159;
wire n_3222;
wire n_325;
wire n_1740;
wire n_4616;
wire n_6011;
wire n_12259;
wire n_11665;
wire n_12975;
wire n_5016;
wire n_9330;
wire n_9367;
wire n_7465;
wire n_11556;
wire n_11685;
wire n_13402;
wire n_14231;
wire n_5470;
wire n_10230;
wire n_11801;
wire n_12117;
wire n_8917;
wire n_12587;
wire n_1092;
wire n_11573;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_9300;
wire n_14489;
wire n_13619;
wire n_14663;
wire n_3868;
wire n_11589;
wire n_11667;
wire n_14395;
wire n_729;
wire n_8230;
wire n_10414;
wire n_6222;
wire n_13110;
wire n_2218;
wire n_12422;
wire n_8352;
wire n_1122;
wire n_7760;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_9918;
wire n_12977;
wire n_13060;
wire n_390;
wire n_6969;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_9496;
wire n_13177;
wire n_8914;
wire n_10953;
wire n_14082;
wire n_8821;
wire n_11446;
wire n_13853;
wire n_8465;
wire n_6587;
wire n_6688;
wire n_8360;
wire n_6505;
wire n_13586;
wire n_9837;
wire n_12772;
wire n_5362;
wire n_8209;
wire n_388;
wire n_8986;
wire n_14701;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_1218;
wire n_3611;
wire n_11633;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_11011;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_7629;
wire n_12145;
wire n_10787;
wire n_6987;
wire n_877;
wire n_3995;
wire n_7567;
wire n_11342;
wire n_8743;
wire n_8963;
wire n_9191;
wire n_3908;
wire n_11812;
wire n_6453;
wire n_9114;
wire n_11142;
wire n_6308;
wire n_13074;
wire n_1055;
wire n_10896;
wire n_8396;
wire n_1395;
wire n_3892;
wire n_13773;
wire n_1346;
wire n_8514;
wire n_12196;
wire n_13482;
wire n_8550;
wire n_1089;
wire n_7449;
wire n_11959;
wire n_8151;
wire n_13927;
wire n_14688;
wire n_1502;
wire n_3501;
wire n_12889;
wire n_1478;
wire n_13096;
wire n_2555;
wire n_3568;
wire n_3216;
wire n_12493;
wire n_9913;
wire n_2708;
wire n_6187;
wire n_735;
wire n_11626;
wire n_6597;
wire n_13810;
wire n_11178;
wire n_12440;
wire n_4844;
wire n_9329;
wire n_13684;
wire n_6220;
wire n_14452;
wire n_12608;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_10598;
wire n_845;
wire n_13008;
wire n_13800;
wire n_7479;
wire n_7882;
wire n_13607;
wire n_1649;
wire n_2470;
wire n_11750;
wire n_13742;
wire n_7517;
wire n_1297;
wire n_9627;
wire n_3551;
wire n_417;
wire n_13412;
wire n_1708;
wire n_11283;
wire n_10271;
wire n_11338;
wire n_5037;
wire n_11295;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_5189;
wire n_4677;
wire n_8070;
wire n_4525;
wire n_8866;
wire n_10402;
wire n_6149;
wire n_11191;
wire n_10064;
wire n_3364;
wire n_11661;
wire n_13329;
wire n_10137;
wire n_2643;
wire n_755;
wire n_9585;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_7878;
wire n_9376;
wire n_4369;
wire n_12515;
wire n_3826;
wire n_5648;
wire n_278;
wire n_2266;
wire n_11644;
wire n_12249;
wire n_6439;
wire n_4324;
wire n_11354;
wire n_842;
wire n_148;
wire n_13537;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_8797;
wire n_14247;
wire n_14462;
wire n_6547;
wire n_13075;
wire n_11126;
wire n_9524;
wire n_7177;
wire n_7902;
wire n_11408;
wire n_12623;
wire n_742;
wire n_5160;
wire n_12971;
wire n_1719;
wire n_2742;
wire n_13051;
wire n_769;
wire n_3671;
wire n_12674;
wire n_2366;
wire n_9606;
wire n_5762;
wire n_1753;
wire n_14419;
wire n_10800;
wire n_5484;
wire n_1372;
wire n_476;
wire n_12026;
wire n_13038;
wire n_14514;
wire n_13812;
wire n_14733;
wire n_10019;
wire n_10762;
wire n_14135;
wire n_1895;
wire n_7353;
wire n_4104;
wire n_11935;
wire n_8054;
wire n_982;
wire n_3791;
wire n_915;
wire n_10047;
wire n_6478;
wire n_11037;
wire n_2008;
wire n_454;
wire n_298;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_13977;
wire n_3199;
wire n_8841;
wire n_11396;
wire n_9084;
wire n_2127;
wire n_14681;
wire n_7050;
wire n_3151;
wire n_7590;
wire n_14453;
wire n_6906;
wire n_403;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_1319;
wire n_3669;
wire n_3367;
wire n_10995;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_606;
wire n_4528;
wire n_2772;
wire n_14036;
wire n_1700;
wire n_10597;
wire n_659;
wire n_1332;
wire n_10561;
wire n_7818;
wire n_509;
wire n_12345;
wire n_7645;
wire n_5385;
wire n_7482;
wire n_1747;
wire n_3990;
wire n_13841;
wire n_14312;
wire n_11726;
wire n_12346;
wire n_5622;
wire n_14522;
wire n_14110;
wire n_10523;
wire n_8618;
wire n_10377;
wire n_1171;
wire n_10243;
wire n_5635;
wire n_4069;
wire n_8538;
wire n_3582;
wire n_8590;
wire n_13883;
wire n_7907;
wire n_9204;
wire n_8970;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_8791;
wire n_14739;
wire n_13724;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_521;
wire n_5910;
wire n_2140;
wire n_10165;
wire n_14776;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_9616;
wire n_9708;
wire n_1400;
wire n_7862;
wire n_10153;
wire n_9130;
wire n_9988;
wire n_3735;
wire n_8703;
wire n_12265;
wire n_7565;
wire n_7410;
wire n_6422;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_12147;
wire n_7721;
wire n_4524;
wire n_9209;
wire n_8061;
wire n_2831;
wire n_10775;
wire n_10173;
wire n_10585;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_12075;
wire n_8754;
wire n_8864;
wire n_5941;
wire n_10985;
wire n_11300;
wire n_4891;
wire n_14294;
wire n_8837;
wire n_12108;
wire n_10999;
wire n_13425;
wire n_2629;
wire n_3369;
wire n_13791;
wire n_8915;
wire n_1257;
wire n_10587;
wire n_1954;
wire n_8784;
wire n_11219;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_11857;
wire n_5597;
wire n_11735;
wire n_2486;
wire n_11986;
wire n_9086;
wire n_1897;
wire n_8768;
wire n_6999;
wire n_8086;
wire n_8072;
wire n_9014;
wire n_12102;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_7539;
wire n_14611;
wire n_9010;
wire n_11637;
wire n_13925;
wire n_6440;
wire n_4977;
wire n_8774;
wire n_14417;
wire n_2492;
wire n_6976;
wire n_7608;
wire n_7234;
wire n_11072;
wire n_12183;
wire n_2939;
wire n_3425;
wire n_13432;
wire n_4876;
wire n_241;
wire n_5021;
wire n_1449;
wire n_12519;
wire n_2900;
wire n_12955;
wire n_797;
wire n_9044;
wire n_2912;
wire n_13538;
wire n_14176;
wire n_5936;
wire n_14650;
wire n_8307;
wire n_595;
wire n_1405;
wire n_3813;
wire n_13774;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_9694;
wire n_1757;
wire n_11421;
wire n_13323;
wire n_10718;
wire n_13214;
wire n_10951;
wire n_10412;
wire n_8470;
wire n_1950;
wire n_2264;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_7830;
wire n_8050;
wire n_3124;
wire n_3811;
wire n_295;
wire n_10310;
wire n_4200;
wire n_190;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_10655;
wire n_9633;
wire n_6165;
wire n_10133;
wire n_12793;
wire n_3463;
wire n_11989;
wire n_10942;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_463;
wire n_1524;
wire n_13192;
wire n_2928;
wire n_13392;
wire n_5505;
wire n_13433;
wire n_12865;
wire n_1118;
wire n_14662;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_469;
wire n_9261;
wire n_11331;
wire n_12285;
wire n_726;
wire n_5504;
wire n_878;
wire n_7348;
wire n_9345;
wire n_11953;
wire n_4118;
wire n_6829;
wire n_11820;
wire n_12478;
wire n_3857;
wire n_3110;
wire n_9375;
wire n_4239;
wire n_9472;
wire n_9764;
wire n_10509;
wire n_8010;
wire n_3157;
wire n_13059;
wire n_12522;
wire n_13451;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_9448;
wire n_6464;
wire n_8802;
wire n_8950;
wire n_5129;
wire n_13199;
wire n_806;
wire n_1350;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_8603;
wire n_9487;
wire n_10639;
wire n_13588;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_11358;
wire n_12413;
wire n_6838;
wire n_13191;
wire n_2700;
wire n_6368;
wire n_14133;
wire n_10690;
wire n_12369;
wire n_12681;
wire n_1616;
wire n_7935;
wire n_2416;
wire n_11118;
wire n_8143;
wire n_11844;
wire n_2064;
wire n_3640;
wire n_9271;
wire n_5663;
wire n_12084;
wire n_5161;
wire n_14132;
wire n_7933;
wire n_12152;
wire n_12726;
wire n_12784;
wire n_1557;
wire n_6640;
wire n_7155;
wire n_9851;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_349;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_12520;
wire n_12511;
wire n_12705;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_11861;
wire n_12761;
wire n_7743;
wire n_13899;
wire n_4990;
wire n_2986;
wire n_8584;
wire n_14443;
wire n_11370;
wire n_13017;
wire n_949;
wire n_2454;
wire n_9101;
wire n_6550;
wire n_6656;
wire n_8153;
wire n_6972;
wire n_3591;
wire n_8574;
wire n_198;
wire n_12832;
wire n_2760;
wire n_4919;
wire n_13422;
wire n_1208;
wire n_7043;
wire n_7986;
wire n_3317;
wire n_8049;
wire n_9927;
wire n_12207;
wire n_13666;
wire n_12782;
wire n_13042;
wire n_7266;
wire n_10621;
wire n_11884;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_554;
wire n_4420;
wire n_7996;
wire n_14513;
wire n_12970;
wire n_10789;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_354;
wire n_5266;
wire n_10496;
wire n_4559;
wire n_4742;
wire n_12384;
wire n_12605;
wire n_5038;
wire n_14724;
wire n_3566;
wire n_10319;
wire n_5800;
wire n_14021;
wire n_8509;
wire n_12408;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_9850;
wire n_4162;
wire n_5766;
wire n_10499;
wire n_14223;
wire n_11717;
wire n_5293;
wire n_10224;
wire n_13234;
wire n_779;
wire n_4790;
wire n_594;
wire n_7035;
wire n_10970;
wire n_4173;
wire n_8354;
wire n_12651;
wire n_5309;
wire n_6047;
wire n_9432;
wire n_3573;
wire n_2943;
wire n_12160;
wire n_13829;
wire n_11464;
wire n_3319;
wire n_11243;
wire n_2247;
wire n_2230;
wire n_9824;
wire n_422;
wire n_14582;
wire n_1269;
wire n_8277;
wire n_7442;
wire n_4727;
wire n_10827;
wire n_1547;
wire n_1438;
wire n_6568;
wire n_3654;
wire n_11473;
wire n_14508;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_10055;
wire n_12638;
wire n_12698;
wire n_4008;
wire n_11654;
wire n_13878;
wire n_10783;
wire n_2158;
wire n_14562;
wire n_8583;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_8681;
wire n_6258;
wire n_1288;
wire n_8644;
wire n_10148;
wire n_7939;
wire n_9884;
wire n_7715;
wire n_11534;
wire n_2173;
wire n_3982;
wire n_10465;
wire n_14040;
wire n_14361;
wire n_11749;
wire n_7350;
wire n_3647;
wire n_7314;
wire n_6026;
wire n_10610;
wire n_8609;
wire n_13955;
wire n_1143;
wire n_9144;
wire n_3973;
wire n_12481;
wire n_8052;
wire n_4799;
wire n_8733;
wire n_9758;
wire n_12078;
wire n_8082;
wire n_5882;
wire n_6700;
wire n_12815;
wire n_7136;
wire n_4534;
wire n_12129;
wire n_5636;
wire n_4960;
wire n_9931;
wire n_7699;
wire n_11546;
wire n_9693;
wire n_12502;
wire n_10830;
wire n_1153;
wire n_9273;
wire n_271;
wire n_465;
wire n_9196;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_10086;
wire n_9029;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_13763;
wire n_562;
wire n_2020;
wire n_7580;
wire n_5606;
wire n_11785;
wire n_6727;
wire n_2310;
wire n_510;
wire n_5911;
wire n_12697;
wire n_7340;
wire n_8080;
wire n_256;
wire n_13437;
wire n_3600;
wire n_10279;
wire n_7303;
wire n_1023;
wire n_10932;
wire n_11440;
wire n_9967;
wire n_12908;
wire n_8819;
wire n_914;
wire n_7870;
wire n_689;
wire n_7568;
wire n_6139;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_7387;
wire n_3190;
wire n_8487;
wire n_13293;
wire n_3027;
wire n_11545;
wire n_11697;
wire n_4011;
wire n_6454;
wire n_3695;
wire n_13487;
wire n_3800;
wire n_13555;
wire n_13239;
wire n_3462;
wire n_10487;
wire n_14579;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_9881;
wire n_2820;
wire n_497;
wire n_3733;
wire n_1165;
wire n_11645;
wire n_3967;
wire n_12512;
wire n_11263;
wire n_12199;
wire n_6333;
wire n_11937;
wire n_7004;
wire n_12584;
wire n_455;
wire n_13854;
wire n_588;
wire n_13361;
wire n_638;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_10910;
wire n_5058;
wire n_8382;
wire n_1417;
wire n_9733;
wire n_3096;
wire n_8517;
wire n_7207;
wire n_8827;
wire n_13558;
wire n_9075;
wire n_11324;
wire n_13954;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_11763;
wire n_13803;
wire n_7167;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_11853;
wire n_2431;
wire n_3322;
wire n_12988;
wire n_14537;
wire n_8906;
wire n_1603;
wire n_5841;
wire n_10109;
wire n_7146;
wire n_7030;
wire n_14542;
wire n_10857;
wire n_4478;
wire n_8203;
wire n_413;
wire n_2935;
wire n_9442;
wire n_4246;
wire n_715;
wire n_7618;
wire n_14625;
wire n_1066;
wire n_2863;
wire n_13244;
wire n_2331;
wire n_4632;
wire n_13305;
wire n_12284;
wire n_11364;
wire n_11941;
wire n_685;
wire n_9630;
wire n_4061;
wire n_11359;
wire n_12031;
wire n_14203;
wire n_9898;
wire n_11323;
wire n_11504;
wire n_11704;
wire n_2920;
wire n_11587;
wire n_1712;
wire n_11620;
wire n_13697;
wire n_3344;
wire n_8340;
wire n_4754;
wire n_12652;
wire n_9582;
wire n_1534;
wire n_8268;
wire n_10865;
wire n_8171;
wire n_1290;
wire n_4375;
wire n_12850;
wire n_617;
wire n_9877;
wire n_14578;
wire n_10179;
wire n_12969;
wire n_2396;
wire n_10925;
wire n_12379;
wire n_12607;
wire n_3368;
wire n_9986;
wire n_13743;
wire n_1559;
wire n_13951;
wire n_14222;
wire n_13695;
wire n_8008;
wire n_7633;
wire n_10246;
wire n_9636;
wire n_3117;
wire n_4684;
wire n_10439;
wire n_743;
wire n_13376;
wire n_14377;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_8553;
wire n_2592;
wire n_8824;
wire n_11902;
wire n_3490;
wire n_7280;
wire n_8369;
wire n_962;
wire n_5043;
wire n_12701;
wire n_14008;
wire n_7339;
wire n_7597;
wire n_8884;
wire n_12898;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_9225;
wire n_4183;
wire n_7768;
wire n_918;
wire n_1968;
wire n_11282;
wire n_5645;
wire n_639;
wire n_5020;
wire n_673;
wire n_6455;
wire n_13639;
wire n_2842;
wire n_7615;
wire n_2196;
wire n_12475;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_10182;
wire n_8271;
wire n_9091;
wire n_3720;
wire n_6183;
wire n_13772;
wire n_14643;
wire n_12027;
wire n_8392;
wire n_8309;
wire n_6107;
wire n_12218;
wire n_10795;
wire n_13602;
wire n_6476;
wire n_5232;
wire n_10046;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_9412;
wire n_11834;
wire n_8874;
wire n_8228;
wire n_12174;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_11405;
wire n_11028;
wire n_3037;
wire n_11663;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_8483;
wire n_6003;
wire n_5443;
wire n_8133;
wire n_7612;
wire n_12385;
wire n_1166;
wire n_2007;
wire n_14407;
wire n_3363;
wire n_6636;
wire n_9525;
wire n_1158;
wire n_11071;
wire n_12289;
wire n_11625;
wire n_1803;
wire n_872;
wire n_11187;
wire n_12041;
wire n_12565;
wire n_3522;
wire n_12882;
wire n_13736;
wire n_13254;
wire n_12819;
wire n_8172;
wire n_4455;
wire n_13341;
wire n_3241;
wire n_3899;
wire n_6554;
wire n_9575;
wire n_5631;
wire n_3481;
wire n_280;
wire n_10456;
wire n_11566;
wire n_10413;
wire n_12164;
wire n_7401;
wire n_11271;
wire n_12433;
wire n_6994;
wire n_11649;
wire n_12224;
wire n_13061;
wire n_5101;
wire n_9738;
wire n_10735;
wire n_6020;
wire n_2236;
wire n_13328;
wire n_9252;
wire n_12550;
wire n_6185;
wire n_8344;
wire n_12800;
wire n_14568;
wire n_692;
wire n_14259;
wire n_7594;
wire n_7711;
wire n_7321;
wire n_4457;
wire n_12561;
wire n_223;
wire n_2150;
wire n_8936;
wire n_8738;
wire n_10822;
wire n_9739;
wire n_6785;
wire n_1816;
wire n_2803;
wire n_9727;
wire n_2887;
wire n_10508;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_13281;
wire n_7574;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_8226;
wire n_6695;
wire n_7529;
wire n_3354;
wire n_5608;
wire n_6501;
wire n_2204;
wire n_11308;
wire n_11739;
wire n_11593;
wire n_9148;
wire n_10858;
wire n_1481;
wire n_2040;
wire n_6466;
wire n_10736;
wire n_11828;
wire n_9958;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_6467;
wire n_9323;
wire n_2231;
wire n_14138;
wire n_4212;
wire n_622;
wire n_4584;
wire n_7522;
wire n_7188;
wire n_9779;
wire n_8088;
wire n_5702;
wire n_14244;
wire n_9545;
wire n_9155;
wire n_8930;
wire n_12563;
wire n_8662;
wire n_13114;
wire n_11291;
wire n_3574;
wire n_11425;
wire n_13566;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_9046;
wire n_9430;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_9625;
wire n_11890;
wire n_13621;
wire n_8783;
wire n_12398;
wire n_13624;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_8663;
wire n_14015;
wire n_10928;
wire n_5277;
wire n_792;
wire n_1262;
wire n_6507;
wire n_10842;
wire n_1942;
wire n_12941;
wire n_6618;
wire n_9447;
wire n_13407;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_13404;
wire n_6213;
wire n_1579;
wire n_8364;
wire n_9485;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_8981;
wire n_9129;
wire n_229;
wire n_8490;
wire n_923;
wire n_12461;
wire n_1124;
wire n_11832;
wire n_7872;
wire n_1326;
wire n_3969;
wire n_6873;
wire n_7958;
wire n_2282;
wire n_4605;
wire n_8118;
wire n_981;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_8671;
wire n_7101;
wire n_12095;
wire n_14191;
wire n_8785;
wire n_11294;
wire n_11470;
wire n_10210;
wire n_1204;
wire n_11744;
wire n_13994;
wire n_7843;
wire n_12998;
wire n_994;
wire n_2428;
wire n_9047;
wire n_13219;
wire n_10057;
wire n_1360;
wire n_6063;
wire n_13737;
wire n_2858;
wire n_12630;
wire n_11641;
wire n_3076;
wire n_7578;
wire n_12789;
wire n_12679;
wire n_14146;
wire n_3410;
wire n_13372;
wire n_5415;
wire n_14084;
wire n_856;
wire n_7261;
wire n_8982;
wire n_10739;
wire n_4592;
wire n_4999;
wire n_1564;
wire n_12327;
wire n_6993;
wire n_9745;
wire n_14288;
wire n_12038;
wire n_508;
wire n_13932;
wire n_10533;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_13978;
wire n_11875;
wire n_8100;
wire n_1858;
wire n_10878;
wire n_353;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_10988;
wire n_1482;
wire n_8522;
wire n_13563;
wire n_1361;
wire n_13141;
wire n_12338;
wire n_10993;
wire n_13249;
wire n_8381;
wire n_9320;
wire n_8835;
wire n_6767;
wire n_11014;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_12030;
wire n_14553;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_6558;
wire n_13517;
wire n_9457;
wire n_9108;
wire n_6755;
wire n_9907;
wire n_10959;
wire n_6153;
wire n_11310;
wire n_3536;
wire n_1721;
wire n_11062;
wire n_7263;
wire n_3782;
wire n_10940;
wire n_12067;
wire n_13783;
wire n_1317;
wire n_12675;
wire n_6608;
wire n_11400;
wire n_11040;
wire n_6202;
wire n_6780;
wire n_7688;
wire n_13968;
wire n_12870;
wire n_14038;
wire n_3594;
wire n_12291;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_7925;
wire n_7245;
wire n_7310;
wire n_9567;
wire n_294;
wire n_6359;
wire n_11773;
wire n_14385;
wire n_5690;
wire n_10583;
wire n_14027;
wire n_11332;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_7585;
wire n_8356;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_13279;
wire n_13731;
wire n_12013;
wire n_13007;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_9852;
wire n_10881;
wire n_12395;
wire n_3855;
wire n_7418;
wire n_14049;
wire n_6353;
wire n_13160;
wire n_2985;
wire n_11943;
wire n_5218;
wire n_10544;
wire n_12933;
wire n_2630;
wire n_7772;
wire n_6577;
wire n_13895;
wire n_14403;
wire n_13213;
wire n_8736;
wire n_2028;
wire n_919;
wire n_3114;
wire n_10491;
wire n_12131;
wire n_2092;
wire n_13507;
wire n_6082;
wire n_11144;
wire n_13385;
wire n_10926;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_11841;
wire n_8918;
wire n_11766;
wire n_2402;
wire n_1458;
wire n_12766;
wire n_679;
wire n_10839;
wire n_220;
wire n_3047;
wire n_10603;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_9022;
wire n_13790;
wire n_7514;
wire n_1550;
wire n_12399;
wire n_1358;
wire n_8616;
wire n_1200;
wire n_6105;
wire n_387;
wire n_12762;
wire n_10400;
wire n_11518;
wire n_826;
wire n_5512;
wire n_13567;
wire n_7738;
wire n_14346;
wire n_2808;
wire n_14787;
wire n_2344;
wire n_8838;
wire n_8908;
wire n_13687;
wire n_3520;
wire n_11960;
wire n_2392;
wire n_7609;
wire n_13580;
wire n_9161;
wire n_3272;
wire n_12241;
wire n_10792;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_11274;
wire n_6548;
wire n_8607;
wire n_13779;
wire n_607;
wire n_8213;
wire n_14487;
wire n_13722;
wire n_13225;
wire n_14615;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_10994;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_13514;
wire n_1268;
wire n_13806;
wire n_2676;
wire n_9903;
wire n_9831;
wire n_14595;
wire n_10032;
wire n_8436;
wire n_7282;
wire n_372;
wire n_13261;
wire n_8551;
wire n_14638;
wire n_13039;
wire n_2770;
wire n_4550;
wire n_14717;
wire n_9238;
wire n_12137;
wire n_14167;
wire n_4347;
wire n_11624;
wire n_10580;
wire n_7921;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_10512;
wire n_9248;
wire n_12495;
wire n_5514;
wire n_11917;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_12790;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_9867;
wire n_12106;
wire n_1282;
wire n_11130;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_10005;
wire n_11053;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_11872;
wire n_5188;
wire n_12434;
wire n_6674;
wire n_13669;
wire n_5049;
wire n_12710;
wire n_2212;
wire n_7489;
wire n_9056;
wire n_6331;
wire n_5308;
wire n_9106;
wire n_311;
wire n_4434;
wire n_13303;
wire n_5068;
wire n_12881;
wire n_7863;
wire n_6493;
wire n_7363;
wire n_14496;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_10596;
wire n_12920;
wire n_4019;
wire n_4199;
wire n_14260;
wire n_7968;
wire n_11220;
wire n_10061;
wire n_10507;
wire n_6023;
wire n_7820;
wire n_8437;
wire n_269;
wire n_816;
wire n_7833;
wire n_12086;
wire n_1322;
wire n_11887;
wire n_3829;
wire n_14189;
wire n_12281;
wire n_12991;
wire n_4510;
wire n_14552;
wire n_7750;
wire n_5057;
wire n_446;
wire n_9071;
wire n_6196;
wire n_12995;
wire n_5425;
wire n_5273;
wire n_10136;
wire n_5839;
wire n_2469;
wire n_7588;
wire n_1125;
wire n_10967;
wire n_11551;
wire n_2358;
wire n_1710;
wire n_14339;
wire n_13368;
wire n_10369;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_10025;
wire n_10708;
wire n_11703;
wire n_7697;
wire n_5887;
wire n_13948;
wire n_7808;
wire n_3068;
wire n_9519;
wire n_1629;
wire n_9027;
wire n_7603;
wire n_13598;
wire n_1094;
wire n_6321;
wire n_14180;
wire n_5683;
wire n_1510;
wire n_8704;
wire n_14341;
wire n_3002;
wire n_8984;
wire n_9786;
wire n_10194;
wire n_7192;
wire n_1099;
wire n_12807;
wire n_5248;
wire n_4899;
wire n_11153;
wire n_10833;
wire n_3146;
wire n_10685;
wire n_3038;
wire n_759;
wire n_10513;
wire n_567;
wire n_4156;
wire n_8613;
wire n_13611;
wire n_1727;
wire n_11030;
wire n_14704;
wire n_3693;
wire n_13178;
wire n_14293;
wire n_10223;
wire n_5880;
wire n_13495;
wire n_8012;
wire n_12012;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_8881;
wire n_5531;
wire n_9404;
wire n_831;
wire n_13777;
wire n_3681;
wire n_5666;
wire n_13301;
wire n_3970;
wire n_11368;
wire n_778;
wire n_2351;
wire n_1619;
wire n_12098;
wire n_7988;
wire n_12025;
wire n_550;
wire n_12669;
wire n_13205;
wire n_3188;
wire n_4448;
wire n_10410;
wire n_13049;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_8763;
wire n_6450;
wire n_9370;
wire n_1152;
wire n_6995;
wire n_2447;
wire n_13009;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_6347;
wire n_13748;
wire n_13338;
wire n_6496;
wire n_13747;
wire n_4776;
wire n_671;
wire n_8387;
wire n_9352;
wire n_11716;
wire n_14083;
wire n_8105;
wire n_10984;
wire n_13485;
wire n_10144;
wire n_12019;
wire n_2704;
wire n_1334;
wire n_6745;
wire n_7943;
wire n_3729;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_13416;
wire n_11967;
wire n_12255;
wire n_7377;
wire n_8900;
wire n_4392;
wire n_3103;
wire n_488;
wire n_6064;
wire n_9681;
wire n_14439;
wire n_8353;
wire n_12503;
wire n_505;
wire n_9051;
wire n_2048;
wire n_7723;
wire n_498;
wire n_3028;
wire n_4691;
wire n_7904;
wire n_3775;
wire n_3148;
wire n_5682;
wire n_684;
wire n_5461;
wire n_9098;
wire n_12415;
wire n_7296;
wire n_3966;
wire n_4397;
wire n_8323;
wire n_13053;
wire n_13752;
wire n_10459;
wire n_12951;
wire n_14125;
wire n_6164;
wire n_11426;
wire n_8711;
wire n_13273;
wire n_3616;
wire n_11628;
wire n_4753;
wire n_12704;
wire n_9484;
wire n_4803;
wire n_8731;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_10155;
wire n_11367;
wire n_6292;
wire n_7759;
wire n_6743;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_11418;
wire n_2852;
wire n_8597;
wire n_2515;
wire n_6330;
wire n_1600;
wire n_1144;
wire n_7178;
wire n_838;
wire n_11026;
wire n_1941;
wire n_7045;
wire n_11576;
wire n_175;
wire n_3637;
wire n_9853;
wire n_8534;
wire n_1017;
wire n_9210;
wire n_8655;
wire n_12884;
wire n_734;
wire n_6923;
wire n_13324;
wire n_4893;
wire n_10915;
wire n_13414;
wire n_13894;
wire n_2240;
wire n_10949;
wire n_7777;
wire n_12339;
wire n_8302;
wire n_14616;
wire n_4258;
wire n_5756;
wire n_14784;
wire n_14695;
wire n_14455;
wire n_310;
wire n_12911;
wire n_8496;
wire n_7693;
wire n_11150;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2432;
wire n_2085;
wire n_10156;
wire n_5033;
wire n_11123;
wire n_14414;
wire n_10248;
wire n_6015;
wire n_1686;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_8078;
wire n_14449;
wire n_2097;
wire n_662;
wire n_11733;
wire n_3461;
wire n_10215;
wire n_10624;
wire n_12915;
wire n_7682;
wire n_10152;
wire n_939;
wire n_1410;
wire n_2297;
wire n_6861;
wire n_12888;
wire n_7300;
wire n_4203;
wire n_12105;
wire n_9756;
wire n_5789;
wire n_12034;
wire n_5400;
wire n_1325;
wire n_7558;
wire n_1223;
wire n_5347;
wire n_14744;
wire n_2957;
wire n_572;
wire n_11188;
wire n_9166;
wire n_8103;
wire n_8719;
wire n_1983;
wire n_10877;
wire n_7798;
wire n_9778;
wire n_8879;
wire n_13906;
wire n_4767;
wire n_8969;
wire n_9141;
wire n_4569;
wire n_11209;
wire n_948;
wire n_448;
wire n_6528;
wire n_14441;
wire n_13159;
wire n_9700;
wire n_10316;
wire n_8896;
wire n_3820;
wire n_5144;
wire n_11503;
wire n_6895;
wire n_3072;
wire n_10385;
wire n_14769;
wire n_14732;
wire n_8335;
wire n_2961;
wire n_13337;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_7400;
wire n_14230;
wire n_11699;
wire n_13145;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_8116;
wire n_12549;
wire n_6523;
wire n_11817;
wire n_5169;
wire n_4885;
wire n_7475;
wire n_14618;
wire n_1479;
wire n_11469;
wire n_9363;
wire n_11971;
wire n_4698;
wire n_14199;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_14722;
wire n_5349;
wire n_14101;
wire n_6472;
wire n_3763;
wire n_9532;
wire n_10823;
wire n_12237;
wire n_933;
wire n_14001;
wire n_6389;
wire n_14586;
wire n_3499;
wire n_14623;
wire n_14635;
wire n_10680;
wire n_5534;
wire n_1821;
wire n_9307;
wire n_13922;
wire n_9876;
wire n_12220;
wire n_3910;
wire n_3947;
wire n_12564;
wire n_492;
wire n_10814;
wire n_12375;
wire n_13333;
wire n_252;
wire n_5183;
wire n_2585;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_8462;
wire n_9959;
wire n_3228;
wire n_8834;
wire n_9989;
wire n_10651;
wire n_14495;
wire n_8417;
wire n_8286;
wire n_2164;
wire n_1732;
wire n_13872;
wire n_12809;
wire n_2678;
wire n_8964;
wire n_10611;
wire n_1186;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_10549;
wire n_10370;
wire n_11621;
wire n_7672;
wire n_10770;
wire n_14171;
wire n_4556;
wire n_6137;
wire n_9467;
wire n_2205;
wire n_2183;
wire n_11558;
wire n_389;
wire n_12043;
wire n_1724;
wire n_3088;
wire n_12513;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_12337;
wire n_1126;
wire n_10393;
wire n_5079;
wire n_8247;
wire n_2761;
wire n_2357;
wire n_10089;
wire n_9406;
wire n_11113;
wire n_14182;
wire n_4520;
wire n_10543;
wire n_895;
wire n_13355;
wire n_8639;
wire n_12504;
wire n_1639;
wire n_11301;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_9160;
wire n_5751;
wire n_11051;
wire n_12489;
wire n_626;
wire n_10321;
wire n_12886;
wire n_13308;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_7712;
wire n_7681;
wire n_6885;
wire n_5039;
wire n_1818;
wire n_6613;
wire n_6580;
wire n_8566;
wire n_8727;
wire n_4265;
wire n_8482;
wire n_13923;
wire n_6120;
wire n_3557;
wire n_13905;
wire n_1598;
wire n_11018;
wire n_6404;
wire n_2269;
wire n_10259;
wire n_7491;
wire n_12836;
wire n_265;
wire n_1583;
wire n_14243;
wire n_13936;
wire n_10909;
wire n_10094;
wire n_8599;
wire n_4612;
wire n_14386;
wire n_5997;
wire n_10302;
wire n_11328;
wire n_8781;
wire n_11276;
wire n_5438;
wire n_9167;
wire n_5375;
wire n_7150;
wire n_7954;
wire n_7974;
wire n_1264;
wire n_6602;
wire n_6530;
wire n_7915;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_6135;
wire n_246;
wire n_12655;
wire n_10623;
wire n_8839;
wire n_11326;
wire n_13627;
wire n_14359;
wire n_14786;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_13882;
wire n_12779;
wire n_8365;
wire n_1102;
wire n_13144;
wire n_14085;
wire n_2239;
wire n_6942;
wire n_7860;
wire n_14108;
wire n_6892;
wire n_1296;
wire n_4730;
wire n_7357;
wire n_8112;
wire n_8489;
wire n_13364;
wire n_8859;
wire n_8060;
wire n_9290;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_882;
wire n_8244;
wire n_2304;
wire n_13134;
wire n_13340;
wire n_2514;
wire n_6977;
wire n_7229;
wire n_12688;
wire n_11732;
wire n_5604;
wire n_10485;
wire n_8096;
wire n_11946;
wire n_7336;
wire n_11334;
wire n_5932;
wire n_289;
wire n_6598;
wire n_10105;
wire n_6795;
wire n_6121;
wire n_11855;
wire n_12321;
wire n_457;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_8346;
wire n_3489;
wire n_5012;
wire n_11781;
wire n_6506;
wire n_13310;
wire n_6614;
wire n_14548;
wire n_14306;
wire n_11080;
wire n_2079;
wire n_9705;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_8367;
wire n_9113;
wire n_10761;
wire n_12104;
wire n_3484;
wire n_6001;
wire n_13445;
wire n_411;
wire n_14043;
wire n_4971;
wire n_9521;
wire n_9682;
wire n_2095;
wire n_14676;
wire n_7493;
wire n_9278;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_14355;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_357;
wire n_3041;
wire n_412;
wire n_5823;
wire n_8898;
wire n_9222;
wire n_1421;
wire n_2423;
wire n_2208;
wire n_5422;
wire n_8905;
wire n_8658;
wire n_5944;
wire n_6989;
wire n_8145;
wire n_8237;
wire n_6299;
wire n_11445;
wire n_12643;
wire n_10592;
wire n_9813;
wire n_7424;
wire n_10216;
wire n_5246;
wire n_8562;
wire n_4376;
wire n_9863;
wire n_3832;
wire n_10616;
wire n_11350;
wire n_14527;
wire n_12799;
wire n_3525;
wire n_13833;
wire n_3712;
wire n_12202;
wire n_12694;
wire n_11057;
wire n_9394;
wire n_10170;
wire n_11182;
wire n_1069;
wire n_4305;
wire n_11140;
wire n_2037;
wire n_2953;
wire n_573;
wire n_2823;
wire n_11082;
wire n_7273;
wire n_9663;
wire n_7901;
wire n_3684;
wire n_14371;
wire n_5725;
wire n_10146;
wire n_5404;
wire n_913;
wire n_10175;
wire n_1681;
wire n_11949;
wire n_13576;
wire n_12055;
wire n_4834;
wire n_9994;
wire n_1507;
wire n_5332;
wire n_9723;
wire n_7149;
wire n_589;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_11693;
wire n_12506;
wire n_8211;
wire n_3268;
wire n_2559;
wire n_8537;
wire n_8946;
wire n_5616;
wire n_1383;
wire n_603;
wire n_8055;
wire n_10848;
wire n_373;
wire n_4259;
wire n_5870;
wire n_7909;
wire n_12788;
wire n_12894;
wire n_2030;
wire n_6053;
wire n_11024;
wire n_850;
wire n_6233;
wire n_10450;
wire n_10918;
wire n_12333;
wire n_13502;
wire n_4299;
wire n_13131;
wire n_5625;
wire n_245;
wire n_13238;
wire n_14597;
wire n_319;
wire n_6758;
wire n_2407;
wire n_690;
wire n_5367;
wire n_9069;
wire n_525;
wire n_2243;
wire n_12866;
wire n_6629;
wire n_5288;
wire n_13247;
wire n_11158;
wire n_2694;
wire n_6356;
wire n_8332;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_7601;
wire n_8998;
wire n_13391;
wire n_14190;
wire n_11046;
wire n_1837;
wire n_7033;
wire n_4178;
wire n_6010;
wire n_11390;
wire n_12551;
wire n_11224;
wire n_13970;
wire n_10536;
wire n_14696;
wire n_189;
wire n_8157;
wire n_2006;
wire n_9284;
wire n_4953;
wire n_10990;
wire n_8484;
wire n_4813;
wire n_3352;
wire n_12223;
wire n_12390;
wire n_12627;
wire n_2367;
wire n_7147;
wire n_7596;
wire n_9556;
wire n_12226;
wire n_14546;
wire n_5294;
wire n_11380;
wire n_8161;
wire n_5570;
wire n_11101;
wire n_6411;
wire n_11578;
wire n_9337;
wire n_2731;
wire n_3703;
wire n_5670;
wire n_5411;
wire n_1246;
wire n_13256;
wire n_11015;
wire n_11214;
wire n_9211;
wire n_12378;
wire n_5265;
wire n_7549;
wire n_5955;
wire n_10278;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_10482;
wire n_14174;
wire n_6032;
wire n_1196;
wire n_10996;
wire n_5733;
wire n_8692;
wire n_3435;
wire n_12794;
wire n_410;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_9243;
wire n_14046;
wire n_12436;
wire n_6918;
wire n_1298;
wire n_10733;
wire n_1745;
wire n_9773;
wire n_14158;
wire n_4674;
wire n_8812;
wire n_14218;
wire n_568;
wire n_11033;
wire n_8682;
wire n_13170;
wire n_4796;
wire n_8290;
wire n_1088;
wire n_7138;
wire n_13664;
wire n_766;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_7976;
wire n_377;
wire n_9928;
wire n_10975;
wire n_2750;
wire n_11950;
wire n_8890;
wire n_10484;
wire n_2547;
wire n_12962;
wire n_8747;
wire n_7617;
wire n_12094;
wire n_279;
wire n_945;
wire n_4575;
wire n_9784;
wire n_10641;
wire n_11115;
wire n_12964;
wire n_3665;
wire n_3063;
wire n_8062;
wire n_14120;
wire n_3281;
wire n_7137;
wire n_3535;
wire n_5061;
wire n_14652;
wire n_2288;
wire n_14412;
wire n_3858;
wire n_14499;
wire n_4653;
wire n_7700;
wire n_11709;
wire n_8275;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_10584;
wire n_14609;
wire n_8667;
wire n_3220;
wire n_4581;
wire n_9192;
wire n_10365;
wire n_14427;
wire n_6008;
wire n_500;
wire n_665;
wire n_10778;
wire n_4625;
wire n_11607;
wire n_11542;
wire n_7098;
wire n_6181;
wire n_14668;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_13105;
wire n_4148;
wire n_9134;
wire n_12838;
wire n_13964;
wire n_3679;
wire n_738;
wire n_5575;
wire n_6654;
wire n_11491;
wire n_7661;
wire n_672;
wire n_4968;
wire n_7801;
wire n_8807;
wire n_9975;
wire n_13766;
wire n_9765;
wire n_11896;
wire n_13525;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_11371;
wire n_11939;
wire n_5316;
wire n_7876;
wire n_2735;
wire n_953;
wire n_14332;
wire n_4214;
wire n_13081;
wire n_10378;
wire n_143;
wire n_1888;
wire n_5290;
wire n_13057;
wire n_1224;
wire n_10324;
wire n_11563;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_557;
wire n_3419;
wire n_7323;
wire n_13861;
wire n_989;
wire n_10850;
wire n_5048;
wire n_11565;
wire n_2233;
wire n_13129;
wire n_13257;
wire n_5363;
wire n_14583;
wire n_11164;
wire n_12633;
wire n_5665;
wire n_6517;
wire n_11401;
wire n_11414;
wire n_795;
wire n_4892;
wire n_6339;
wire n_10330;
wire n_12514;
wire n_14408;
wire n_14659;
wire n_1936;
wire n_9564;
wire n_14267;
wire n_9127;
wire n_11199;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_8048;
wire n_821;
wire n_770;
wire n_14370;
wire n_5607;
wire n_1514;
wire n_7929;
wire n_14516;
wire n_486;
wire n_2782;
wire n_569;
wire n_3929;
wire n_11319;
wire n_9306;
wire n_971;
wire n_4353;
wire n_2201;
wire n_8212;
wire n_4950;
wire n_10442;
wire n_1650;
wire n_7755;
wire n_6504;
wire n_9891;
wire n_13865;
wire n_13135;
wire n_10962;
wire n_10022;
wire n_13973;
wire n_4176;
wire n_9078;
wire n_7556;
wire n_222;
wire n_11415;
wire n_13553;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_10972;
wire n_7216;
wire n_13248;
wire n_6814;
wire n_4488;
wire n_10127;
wire n_5278;
wire n_14278;
wire n_2779;
wire n_3627;
wire n_10824;
wire n_3596;
wire n_5214;
wire n_11128;
wire n_9332;
wire n_12262;
wire n_3756;
wire n_12391;
wire n_8223;
wire n_8043;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_8159;
wire n_5845;
wire n_8868;
wire n_9889;
wire n_4608;
wire n_9294;
wire n_12731;
wire n_6691;
wire n_13623;
wire n_432;
wire n_293;
wire n_13775;
wire n_12235;
wire n_3948;
wire n_4839;
wire n_9174;
wire n_1074;
wire n_5969;
wire n_10375;
wire n_1765;
wire n_9132;
wire n_13464;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_11669;
wire n_4184;
wire n_206;
wire n_2332;
wire n_9547;
wire n_2391;
wire n_12406;
wire n_6343;
wire n_6005;
wire n_611;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_6686;
wire n_4032;
wire n_12929;
wire n_2571;
wire n_136;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_14067;
wire n_2874;
wire n_6536;
wire n_6029;
wire n_6684;
wire n_4117;
wire n_300;
wire n_6025;
wire n_12229;
wire n_3049;
wire n_8434;
wire n_14264;
wire n_3634;
wire n_12508;
wire n_5436;
wire n_7962;
wire n_2341;
wire n_1654;
wire n_6697;
wire n_11262;
wire n_12271;
wire n_3066;
wire n_11110;
wire n_12803;
wire n_2045;
wire n_13084;
wire n_14451;
wire n_14614;
wire n_10122;
wire n_10898;
wire n_6085;
wire n_3913;
wire n_14785;
wire n_9762;
wire n_11849;
wire n_5341;
wire n_8608;
wire n_2575;
wire n_13583;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_376;
wire n_13470;
wire n_1597;
wire n_12245;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_14394;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_8656;
wire n_3861;
wire n_5096;
wire n_9183;
wire n_2043;
wire n_11287;
wire n_7905;
wire n_6771;
wire n_4171;
wire n_11247;
wire n_5847;
wire n_7204;
wire n_12376;
wire n_9461;
wire n_9117;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_12773;
wire n_4665;
wire n_6877;
wire n_7308;
wire n_10116;
wire n_7476;
wire n_10590;
wire n_10991;
wire n_11945;
wire n_5639;
wire n_14743;
wire n_11769;
wire n_4884;
wire n_3580;
wire n_12720;
wire n_1437;
wire n_12736;
wire n_8249;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_9062;
wire n_209;
wire n_5240;
wire n_5503;
wire n_1461;
wire n_7208;
wire n_9915;
wire n_10265;
wire n_7718;
wire n_5718;
wire n_13006;
wire n_11277;
wire n_1876;
wire n_1830;
wire n_12459;
wire n_11075;
wire n_5001;
wire n_12708;
wire n_6567;
wire n_11919;
wire n_503;
wire n_12387;
wire n_13705;
wire n_5658;
wire n_1112;
wire n_700;
wire n_4174;
wire n_9001;
wire n_13599;
wire n_6868;
wire n_13077;
wire n_5131;
wire n_7290;
wire n_9081;
wire n_6813;
wire n_7756;
wire n_9156;
wire n_5546;
wire n_6294;
wire n_7795;
wire n_7822;
wire n_8717;
wire n_10159;
wire n_5174;
wire n_9024;
wire n_9198;
wire n_10178;
wire n_2145;
wire n_4801;
wire n_10571;
wire n_6079;
wire n_6260;
wire n_680;
wire n_4582;
wire n_14268;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_7623;
wire n_13892;
wire n_380;
wire n_14251;
wire n_12239;
wire n_14136;
wire n_12636;
wire n_14002;
wire n_3119;
wire n_6671;
wire n_11085;
wire n_9335;
wire n_4740;
wire n_1108;
wire n_10550;
wire n_9488;
wire n_1274;
wire n_7632;
wire n_4394;
wire n_257;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_11510;
wire n_9725;
wire n_8842;
wire n_475;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_8073;
wire n_10185;
wire n_12648;
wire n_9526;
wire n_4920;
wire n_3909;
wire n_10809;
wire n_13316;
wire n_4220;
wire n_2703;
wire n_13140;
wire n_5069;
wire n_5541;
wire n_13162;
wire n_10660;
wire n_6314;
wire n_12501;
wire n_577;
wire n_5610;
wire n_407;
wire n_9962;
wire n_8576;
wire n_916;
wire n_2810;
wire n_12755;
wire n_6703;
wire n_5571;
wire n_1884;
wire n_14262;
wire n_1555;
wire n_10657;
wire n_10627;
wire n_8799;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_9667;
wire n_5166;
wire n_2683;
wire n_11256;
wire n_6065;
wire n_7265;
wire n_12441;
wire n_14018;
wire n_4180;
wire n_11516;
wire n_11520;
wire n_4459;
wire n_6878;
wire n_11461;
wire n_11137;
wire n_3624;
wire n_6725;
wire n_8181;
wire n_5808;
wire n_1182;
wire n_6527;
wire n_4594;
wire n_13604;
wire n_8447;
wire n_8045;
wire n_7289;
wire n_7538;
wire n_14029;
wire n_13157;
wire n_2748;
wire n_11536;
wire n_11544;
wire n_14488;
wire n_10897;
wire n_4642;
wire n_13952;
wire n_14234;
wire n_9716;
wire n_6913;
wire n_1376;
wire n_7473;
wire n_7242;
wire n_9253;
wire n_6533;
wire n_513;
wire n_11305;
wire n_14126;
wire n_179;
wire n_7164;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_8022;
wire n_10617;
wire n_12011;
wire n_3544;
wire n_6845;
wire n_10451;
wire n_5300;
wire n_8227;
wire n_14438;
wire n_10768;
wire n_7853;
wire n_2072;
wire n_3852;
wire n_11268;
wire n_13707;
wire n_5233;
wire n_12742;
wire n_10309;
wire n_5381;
wire n_436;
wire n_9796;
wire n_5770;
wire n_7483;
wire n_13868;
wire n_8756;
wire n_5710;
wire n_10021;
wire n_324;
wire n_10053;
wire n_1491;
wire n_2628;
wire n_7389;
wire n_3219;
wire n_10315;
wire n_9953;
wire n_274;
wire n_1083;
wire n_5333;
wire n_5799;
wire n_10765;
wire n_6265;
wire n_4914;
wire n_12317;
wire n_8604;
wire n_12831;
wire n_8809;
wire n_13092;
wire n_8976;
wire n_11815;
wire n_13694;
wire n_3510;
wire n_10907;
wire n_7046;
wire n_13928;
wire n_7834;
wire n_10312;
wire n_11299;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_11273;
wire n_8940;
wire n_5008;
wire n_1312;
wire n_9077;
wire n_12872;
wire n_13147;
wire n_12871;
wire n_3871;
wire n_13212;
wire n_12590;
wire n_14503;
wire n_892;
wire n_14325;
wire n_3757;
wire n_1567;
wire n_563;
wire n_11213;
wire n_13519;
wire n_2219;
wire n_8844;
wire n_6148;
wire n_8995;
wire n_2100;
wire n_8255;
wire n_3666;
wire n_5538;
wire n_990;
wire n_6357;
wire n_867;
wire n_8216;
wire n_8693;
wire n_12785;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_13661;
wire n_9123;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_6522;
wire n_7811;
wire n_12545;
wire n_8669;
wire n_4285;
wire n_7097;
wire n_12531;
wire n_7000;
wire n_2668;
wire n_10486;
wire n_11290;
wire n_2701;
wire n_2400;
wire n_10357;
wire n_650;
wire n_3741;
wire n_9922;
wire n_5582;
wire n_2567;
wire n_9177;
wire n_14348;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_7880;
wire n_14130;
wire n_712;
wire n_8769;
wire n_9463;
wire n_909;
wire n_12916;
wire n_6713;
wire n_8149;
wire n_1392;
wire n_10067;
wire n_13163;
wire n_12953;
wire n_10698;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_7851;
wire n_13106;
wire n_13874;
wire n_2220;
wire n_13246;
wire n_7342;
wire n_7044;
wire n_7810;
wire n_10135;
wire n_13776;
wire n_6108;
wire n_12222;
wire n_10260;
wire n_7664;
wire n_12370;
wire n_6100;
wire n_14329;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_11412;
wire n_2829;
wire n_7332;
wire n_14428;
wire n_8990;
wire n_5862;
wire n_471;
wire n_7477;
wire n_1914;
wire n_14617;
wire n_10268;
wire n_8208;
wire n_2253;
wire n_7468;
wire n_11550;
wire n_12692;
wire n_13640;
wire n_5886;
wire n_9451;
wire n_7714;
wire n_7899;
wire n_8710;
wire n_12976;
wire n_6415;
wire n_8479;
wire n_6783;
wire n_14660;
wire n_2130;
wire n_4861;
wire n_13984;
wire n_12397;
wire n_2021;
wire n_8512;
wire n_14524;
wire n_13093;
wire n_9843;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_9710;
wire n_2507;
wire n_12634;
wire n_13288;
wire n_1633;
wire n_9087;
wire n_4621;
wire n_14287;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_7845;
wire n_11619;
wire n_13086;
wire n_347;
wire n_2434;
wire n_14052;
wire n_183;
wire n_14216;
wire n_1234;
wire n_3936;
wire n_479;
wire n_5564;
wire n_2261;
wire n_12613;
wire n_9956;
wire n_3082;
wire n_9079;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_12946;
wire n_5802;
wire n_9782;
wire n_10049;
wire n_4784;
wire n_14206;
wire n_13012;
wire n_13606;
wire n_2438;
wire n_12901;
wire n_13449;
wire n_10589;
wire n_3210;
wire n_6340;
wire n_13099;
wire n_14475;
wire n_9950;
wire n_11019;
wire n_14620;
wire n_7858;
wire n_11580;
wire n_3867;
wire n_3397;
wire n_13699;
wire n_12683;
wire n_6103;
wire n_1646;
wire n_6392;
wire n_6513;
wire n_11642;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_13389;
wire n_9197;
wire n_1237;
wire n_6720;
wire n_12286;
wire n_11076;
wire n_11752;
wire n_5883;
wire n_9140;
wire n_14134;
wire n_13995;
wire n_10785;
wire n_14726;
wire n_13439;
wire n_8401;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_14122;
wire n_3971;
wire n_12146;
wire n_370;
wire n_7680;
wire n_14415;
wire n_5630;
wire n_6666;
wire n_286;
wire n_9452;
wire n_9364;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_9398;
wire n_9362;
wire n_13675;
wire n_13483;
wire n_1531;
wire n_2113;
wire n_6815;
wire n_14321;
wire n_9203;
wire n_1387;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_9712;
wire n_9536;
wire n_12054;
wire n_8450;
wire n_9848;
wire n_12081;
wire n_13614;
wire n_14095;
wire n_11202;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_9460;
wire n_5929;
wire n_7710;
wire n_8788;
wire n_5394;
wire n_14080;
wire n_8324;
wire n_11227;
wire n_4751;
wire n_5975;
wire n_4242;
wire n_13814;
wire n_10381;
wire n_9841;
wire n_14502;
wire n_1951;
wire n_12557;
wire n_2490;
wire n_2558;
wire n_9772;
wire n_1496;
wire n_10147;
wire n_2812;
wire n_9057;
wire n_10554;
wire n_3300;
wire n_7061;
wire n_8104;
wire n_9068;
wire n_11860;
wire n_7066;
wire n_5496;
wire n_7485;
wire n_3104;
wire n_7174;
wire n_8014;
wire n_12213;
wire n_4122;
wire n_6661;
wire n_10919;
wire n_12646;
wire n_2132;
wire n_14750;
wire n_4522;
wire n_10228;
wire n_14159;
wire n_5991;
wire n_8623;
wire n_14077;
wire n_14518;
wire n_4952;
wire n_9634;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_9348;
wire n_11125;
wire n_3946;
wire n_5920;
wire n_13011;
wire n_12737;
wire n_2112;
wire n_2640;
wire n_8651;
wire n_10699;
wire n_5000;
wire n_6125;
wire n_4634;
wire n_9632;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_14358;
wire n_12092;
wire n_2237;
wire n_11951;
wire n_2983;
wire n_5211;
wire n_9257;
wire n_4089;
wire n_11451;
wire n_11816;
wire n_9500;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_9747;
wire n_2350;
wire n_9470;
wire n_11508;
wire n_6414;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_14467;
wire n_7783;
wire n_11232;
wire n_7662;
wire n_6057;
wire n_6936;
wire n_10188;
wire n_13531;
wire n_11138;
wire n_9591;
wire n_14373;
wire n_9049;
wire n_487;
wire n_4728;
wire n_7171;
wire n_7990;
wire n_1886;
wire n_4346;
wire n_13585;
wire n_1648;
wire n_7003;
wire n_10433;
wire n_8137;
wire n_2187;
wire n_10231;
wire n_1413;
wire n_8413;
wire n_10841;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_10929;
wire n_12642;
wire n_13142;
wire n_6916;
wire n_2327;
wire n_158;
wire n_3882;
wire n_13974;
wire n_9471;
wire n_3916;
wire n_6922;
wire n_14656;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_14070;
wire n_10582;
wire n_13494;
wire n_12601;
wire n_2841;
wire n_405;
wire n_10719;
wire n_3332;
wire n_8300;
wire n_8069;
wire n_10934;
wire n_7501;
wire n_10747;
wire n_11383;
wire n_320;
wire n_9409;
wire n_10711;
wire n_10743;
wire n_11088;
wire n_6432;
wire n_12959;
wire n_7984;
wire n_12899;
wire n_2055;
wire n_12616;
wire n_2998;
wire n_7366;
wire n_1423;
wire n_10481;
wire n_4359;
wire n_8173;
wire n_13562;
wire n_481;
wire n_1609;
wire n_13540;
wire n_12919;
wire n_2822;
wire n_2308;
wire n_1939;
wire n_2242;
wire n_7589;
wire n_13568;
wire n_13642;
wire n_4447;
wire n_14764;
wire n_2937;
wire n_4293;
wire n_218;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_9832;
wire n_4039;
wire n_12010;
wire n_12314;
wire n_5793;
wire n_14632;
wire n_6926;
wire n_1798;
wire n_8091;
wire n_13751;
wire n_3057;
wire n_1608;
wire n_12394;
wire n_12856;
wire n_5761;
wire n_13465;
wire n_6699;
wire n_12797;
wire n_547;
wire n_13683;
wire n_13630;
wire n_439;
wire n_677;
wire n_3983;
wire n_9067;
wire n_8254;
wire n_703;
wire n_8400;
wire n_10141;
wire n_11090;
wire n_14661;
wire n_10305;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_9858;
wire n_7511;
wire n_326;
wire n_10936;
wire n_12134;
wire n_227;
wire n_13824;
wire n_12730;
wire n_3773;
wire n_3494;
wire n_9482;
wire n_1278;
wire n_9033;
wire n_6957;
wire n_11429;
wire n_5074;
wire n_14624;
wire n_12735;
wire n_14510;
wire n_7917;
wire n_11908;
wire n_3788;
wire n_3939;
wire n_727;
wire n_590;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_8368;
wire n_6694;
wire n_545;
wire n_9247;
wire n_2496;
wire n_3260;
wire n_8463;
wire n_536;
wire n_9965;
wire n_10425;
wire n_3349;
wire n_6449;
wire n_10862;
wire n_12254;
wire n_14333;
wire n_4348;
wire n_1602;
wire n_7422;
wire n_9299;
wire n_13357;
wire n_3139;
wire n_8889;
wire n_427;
wire n_3801;
wire n_5681;
wire n_9785;
wire n_9244;
wire n_11298;
wire n_14667;
wire n_2338;
wire n_5261;
wire n_12427;
wire n_1080;
wire n_12124;
wire n_9195;
wire n_8322;
wire n_11353;
wire n_12494;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_8987;
wire n_13454;
wire n_3653;
wire n_3823;
wire n_9280;
wire n_3403;
wire n_7621;
wire n_9911;
wire n_12051;
wire n_8274;
wire n_13958;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_1205;
wire n_6195;
wire n_163;
wire n_2716;
wire n_10373;
wire n_6441;
wire n_11116;
wire n_7572;
wire n_7158;
wire n_13637;
wire n_11173;
wire n_314;
wire n_2944;
wire n_11660;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_7500;
wire n_1202;
wire n_4084;
wire n_627;
wire n_12355;
wire n_7985;
wire n_9687;
wire n_1371;
wire n_4240;
wire n_8657;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_11567;
wire n_233;
wire n_8954;
wire n_2774;
wire n_6354;
wire n_11881;
wire n_10563;
wire n_12458;
wire n_2799;
wire n_8311;
wire n_5748;
wire n_4393;
wire n_11363;
wire n_321;
wire n_6662;
wire n_7494;
wire n_9088;
wire n_3984;
wire n_1586;
wire n_14050;
wire n_8728;
wire n_9580;
wire n_11280;
wire n_9569;
wire n_1431;
wire n_8994;
wire n_4389;
wire n_6433;
wire n_9680;
wire n_1763;
wire n_8398;
wire n_6200;
wire n_5641;
wire n_12463;
wire n_12612;
wire n_8407;
wire n_8071;
wire n_13423;
wire n_13046;
wire n_4461;
wire n_2763;
wire n_11636;
wire n_3156;
wire n_10530;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_6902;
wire n_4615;
wire n_3492;
wire n_3044;
wire n_12798;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_8528;
wire n_14088;
wire n_9227;
wire n_13644;
wire n_5657;
wire n_12510;
wire n_11313;
wire n_14364;
wire n_8475;
wire n_297;
wire n_9951;
wire n_9855;
wire n_2379;
wire n_3579;
wire n_9072;
wire n_12635;
wire n_10102;
wire n_13545;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_12537;
wire n_4067;
wire n_13197;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_12076;
wire n_5114;
wire n_9054;
wire n_4551;
wire n_178;
wire n_10117;
wire n_551;
wire n_4521;
wire n_13252;
wire n_6956;
wire n_13139;
wire n_10126;
wire n_7587;
wire n_2284;
wire n_6451;
wire n_12874;
wire n_11920;
wire n_3005;
wire n_7704;
wire n_10604;
wire n_5420;
wire n_8511;
wire n_6497;
wire n_7865;
wire n_2283;
wire n_5206;
wire n_582;
wire n_2526;
wire n_13356;
wire n_1097;
wire n_14447;
wire n_1711;
wire n_4387;
wire n_14237;
wire n_14745;
wire n_9584;
wire n_9287;
wire n_534;
wire n_2508;
wire n_3186;
wire n_10344;
wire n_10568;
wire n_9459;
wire n_9490;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_6701;
wire n_10209;
wire n_8867;
wire n_3417;
wire n_8246;
wire n_560;
wire n_8558;
wire n_890;
wire n_9655;
wire n_13769;
wire n_9846;
wire n_3626;
wire n_12048;
wire n_451;
wire n_9593;
wire n_4598;
wire n_4464;
wire n_12072;
wire n_8925;
wire n_5106;
wire n_7881;
wire n_11317;
wire n_9147;
wire n_13339;
wire n_4789;
wire n_3180;
wire n_14433;
wire n_12829;
wire n_3423;
wire n_14672;
wire n_1081;
wire n_9678;
wire n_10803;
wire n_2119;
wire n_12132;
wire n_13626;
wire n_11903;
wire n_8641;
wire n_9658;
wire n_10299;
wire n_2493;
wire n_9560;
wire n_12528;
wire n_9578;
wire n_11813;
wire n_14195;
wire n_5080;
wire n_535;
wire n_9396;
wire n_4565;
wire n_7032;
wire n_12745;
wire n_9303;
wire n_3392;
wire n_12371;
wire n_1800;
wire n_11811;
wire n_12841;
wire n_7198;
wire n_12417;
wire n_6884;
wire n_7752;
wire n_10618;
wire n_10836;
wire n_11378;
wire n_5081;
wire n_8201;
wire n_6921;
wire n_2904;
wire n_12180;
wire n_12049;
wire n_3353;
wire n_2946;
wire n_7953;
wire n_6106;
wire n_14434;
wire n_6876;
wire n_3512;
wire n_9553;
wire n_12603;
wire n_1734;
wire n_1860;
wire n_4552;
wire n_8046;
wire n_12978;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_14575;
wire n_10930;
wire n_6172;
wire n_14005;
wire n_9942;
wire n_9805;
wire n_13686;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_12466;
wire n_13842;
wire n_4040;
wire n_8414;
wire n_3024;
wire n_5567;
wire n_8292;
wire n_9879;
wire n_9138;
wire n_5406;
wire n_8647;
wire n_11936;
wire n_6362;
wire n_9213;
wire n_12071;
wire n_4328;
wire n_12982;
wire n_8543;
wire n_14680;
wire n_13459;
wire n_1854;
wire n_666;
wire n_11543;
wire n_11184;
wire n_11795;
wire n_5191;
wire n_11391;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_11646;
wire n_6833;
wire n_4940;
wire n_9374;
wire n_785;
wire n_3161;
wire n_13649;
wire n_2389;
wire n_14720;
wire n_14497;
wire n_1309;
wire n_8331;
wire n_999;
wire n_2280;
wire n_8317;
wire n_7126;
wire n_12578;
wire n_12311;
wire n_11963;
wire n_5867;
wire n_14109;
wire n_13253;
wire n_456;
wire n_12985;
wire n_12232;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_12640;
wire n_7496;
wire n_13729;
wire n_6430;
wire n_11435;
wire n_13647;
wire n_9179;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_10014;
wire n_4112;
wire n_342;
wire n_11056;
wire n_10714;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_7196;
wire n_14241;
wire n_2614;
wire n_12101;
wire n_11120;
wire n_11185;
wire n_7360;
wire n_5428;
wire n_10895;
wire n_6325;
wire n_10916;
wire n_14693;
wire n_12197;
wire n_2494;
wire n_12497;
wire n_1538;
wire n_4865;
wire n_6678;
wire n_10838;
wire n_7982;
wire n_13002;
wire n_2128;
wire n_4071;
wire n_8929;
wire n_8174;
wire n_6564;
wire n_8187;
wire n_10108;
wire n_7268;
wire n_14069;
wire n_4436;
wire n_5822;
wire n_5786;
wire n_3586;
wire n_10661;
wire n_8846;
wire n_5817;
wire n_9277;
wire n_4160;
wire n_14754;
wire n_6109;
wire n_9611;
wire n_6385;
wire n_1668;
wire n_12571;
wire n_9744;
wire n_5798;
wire n_10123;
wire n_4137;
wire n_1078;
wire n_13022;
wire n_8032;
wire n_9504;
wire n_5417;
wire n_14118;
wire n_14445;
wire n_11147;
wire n_10048;
wire n_4545;
wire n_11194;
wire n_8200;
wire n_4758;
wire n_1161;
wire n_8036;
wire n_9285;
wire n_5713;
wire n_4840;
wire n_9905;
wire n_10963;
wire n_11016;
wire n_12228;
wire n_11146;
wire n_3097;
wire n_13088;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_10788;
wire n_14142;
wire n_9190;
wire n_8586;
wire n_8524;
wire n_618;
wire n_1191;
wire n_11924;
wire n_12540;
wire n_4535;
wire n_7518;
wire n_9639;
wire n_10422;
wire n_12001;
wire n_4385;
wire n_8828;
wire n_7779;
wire n_12059;
wire n_9664;
wire n_1215;
wire n_13275;
wire n_11830;
wire n_14577;
wire n_3748;
wire n_4731;
wire n_7575;
wire n_11489;
wire n_2337;
wire n_13026;
wire n_7073;
wire n_8092;
wire n_10471;
wire n_13760;
wire n_12479;
wire n_10979;
wire n_1786;
wire n_6309;
wire n_8370;
wire n_3732;
wire n_9109;
wire n_211;
wire n_1804;
wire n_10189;
wire n_408;
wire n_13820;
wire n_8135;
wire n_12702;
wire n_6519;
wire n_4671;
wire n_14366;
wire n_9741;
wire n_2272;
wire n_5989;
wire n_4766;
wire n_10569;
wire n_592;
wire n_4558;
wire n_13116;
wire n_13663;
wire n_14055;
wire n_10686;
wire n_1318;
wire n_14197;
wire n_8764;
wire n_14454;
wire n_1769;
wire n_1632;
wire n_7349;
wire n_1929;
wire n_9875;
wire n_10713;
wire n_11411;
wire n_8502;
wire n_4319;
wire n_9360;
wire n_6585;
wire n_12211;
wire n_14323;
wire n_7786;
wire n_10913;
wire n_9021;
wire n_8454;
wire n_2929;
wire n_12306;
wire n_4358;
wire n_11145;
wire n_9122;
wire n_1526;
wire n_7579;
wire n_10099;
wire n_12335;
wire n_12637;
wire n_7122;
wire n_10193;
wire n_14096;
wire n_4874;
wire n_180;
wire n_2656;
wire n_4904;
wire n_516;
wire n_1997;
wire n_10203;
wire n_10140;
wire n_13982;
wire n_1137;
wire n_1733;
wire n_640;
wire n_1258;
wire n_6490;
wire n_7867;
wire n_4651;
wire n_10920;
wire n_10149;
wire n_943;
wire n_11000;
wire n_11712;
wire n_14068;
wire n_4748;
wire n_3167;
wire n_14019;
wire n_7624;
wire n_13405;
wire n_9803;
wire n_13828;
wire n_14397;
wire n_1807;
wire n_1123;
wire n_8776;
wire n_10576;
wire n_2857;
wire n_8564;
wire n_12114;
wire n_8343;
wire n_7828;
wire n_14319;
wire n_1784;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_8718;
wire n_13102;
wire n_13550;
wire n_14301;
wire n_10682;
wire n_752;
wire n_985;
wire n_5506;
wire n_7543;
wire n_9659;
wire n_12204;
wire n_13643;
wire n_5475;
wire n_8042;
wire n_7727;
wire n_2412;
wire n_14774;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_9013;
wire n_5431;
wire n_9427;
wire n_12325;
wire n_8379;
wire n_643;
wire n_8034;
wire n_12143;
wire n_226;
wire n_7778;
wire n_5100;
wire n_2383;
wire n_10225;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_7019;
wire n_682;
wire n_9126;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_9474;
wire n_2907;
wire n_8441;
wire n_14026;
wire n_5752;
wire n_14362;
wire n_1429;
wire n_2353;
wire n_7702;
wire n_14114;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_686;
wire n_10368;
wire n_1154;
wire n_584;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_10237;
wire n_14504;
wire n_9538;
wire n_3718;
wire n_6685;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_8569;
wire n_9574;
wire n_10531;
wire n_12032;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_12066;
wire n_14471;
wire n_8865;
wire n_8592;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_7952;
wire n_11170;
wire n_7347;
wire n_9450;
wire n_3736;
wire n_10031;
wire n_4466;
wire n_6016;
wire n_9998;
wire n_891;
wire n_13963;
wire n_885;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_11523;
wire n_5322;
wire n_1864;
wire n_11121;
wire n_12176;
wire n_5414;
wire n_11805;
wire n_3086;
wire n_13266;
wire n_1887;
wire n_3165;
wire n_7791;
wire n_6971;
wire n_8362;
wire n_10847;
wire n_3336;
wire n_8632;
wire n_10035;
wire n_14242;
wire n_14523;
wire n_7739;
wire n_396;
wire n_12740;
wire n_7945;
wire n_9372;
wire n_9045;
wire n_8361;
wire n_9657;
wire n_7656;
wire n_11457;
wire n_5903;
wire n_7199;
wire n_10107;
wire n_3635;
wire n_11725;
wire n_3541;
wire n_2502;
wire n_10283;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_9904;
wire n_12344;
wire n_9924;
wire n_9159;
wire n_9326;
wire n_6549;
wire n_725;
wire n_8611;
wire n_8561;
wire n_8410;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_6658;
wire n_11694;
wire n_5369;
wire n_9476;
wire n_6683;
wire n_3067;
wire n_154;
wire n_3809;
wire n_4921;
wire n_473;
wire n_1852;
wire n_801;
wire n_5912;
wire n_11540;
wire n_5745;
wire n_7923;
wire n_6086;
wire n_4377;
wire n_818;
wire n_10050;
wire n_11058;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_8878;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_12203;
wire n_1877;
wire n_11403;
wire n_272;
wire n_8492;
wire n_9301;
wire n_14099;
wire n_7213;
wire n_4301;
wire n_5313;
wire n_10392;
wire n_2133;
wire n_14041;
wire n_12769;
wire n_8888;
wire n_6820;
wire n_2497;
wire n_879;
wire n_5446;
wire n_11741;
wire n_7610;
wire n_11245;
wire n_7107;
wire n_4561;
wire n_14225;
wire n_1541;
wire n_597;
wire n_3291;
wire n_7456;
wire n_9382;
wire n_11784;
wire n_8095;
wire n_11365;
wire n_13291;
wire n_14756;
wire n_9921;
wire n_7369;
wire n_1472;
wire n_9325;
wire n_1050;
wire n_9945;
wire n_9643;
wire n_7548;
wire n_11005;
wire n_13016;
wire n_2578;
wire n_12820;
wire n_152;
wire n_1201;
wire n_8735;
wire n_7598;
wire n_1185;
wire n_2475;
wire n_8808;
wire n_7250;
wire n_9201;
wire n_8902;
wire n_7823;
wire n_9771;
wire n_8833;
wire n_14605;
wire n_12869;
wire n_4715;
wire n_6157;
wire n_8796;
wire n_2715;
wire n_335;
wire n_14413;
wire n_2665;
wire n_4879;
wire n_344;
wire n_13435;
wire n_8794;
wire n_12689;
wire n_11074;
wire n_5044;
wire n_210;
wire n_1090;
wire n_3755;
wire n_4536;
wire n_9274;
wire n_9894;
wire n_11141;
wire n_12750;
wire n_14753;
wire n_8549;
wire n_14161;
wire n_6676;
wire n_4304;
wire n_10095;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_14285;
wire n_10716;
wire n_11102;
wire n_12171;
wire n_14000;
wire n_224;
wire n_10088;
wire n_11238;
wire n_11406;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_10443;
wire n_10488;
wire n_7525;
wire n_4418;
wire n_7924;
wire n_3341;
wire n_11103;
wire n_12420;
wire n_9232;
wire n_8690;
wire n_4125;
wire n_5390;
wire n_12954;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_11852;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_12500;
wire n_1511;
wire n_8593;
wire n_11837;
wire n_10912;
wire n_13501;
wire n_10469;
wire n_276;
wire n_13533;
wire n_9649;
wire n_11684;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_12112;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_538;
wire n_2845;
wire n_4412;
wire n_4151;
wire n_2036;
wire n_7649;
wire n_8195;
wire n_843;
wire n_8009;
wire n_8588;
wire n_9839;
wire n_10887;
wire n_3358;
wire n_12004;
wire n_6704;
wire n_7634;
wire n_9090;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_7406;
wire n_13520;
wire n_4682;
wire n_1128;
wire n_9346;
wire n_11012;
wire n_6673;
wire n_14480;
wire n_9696;
wire n_2419;
wire n_11041;
wire n_14181;
wire n_10742;
wire n_2330;
wire n_14024;
wire n_11798;
wire n_12614;
wire n_13165;
wire n_9996;
wire n_6534;
wire n_9968;
wire n_8805;
wire n_5078;
wire n_4810;
wire n_7659;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_6127;
wire n_10405;
wire n_9498;
wire n_9383;
wire n_1440;
wire n_6246;
wire n_10390;
wire n_11978;
wire n_1370;
wire n_10989;
wire n_305;
wire n_9836;
wire n_5005;
wire n_14570;
wire n_14702;
wire n_11827;
wire n_10328;
wire n_13315;
wire n_10692;
wire n_6126;
wire n_7372;
wire n_8596;
wire n_9938;
wire n_12912;
wire n_1549;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_10867;
wire n_6841;
wire n_11847;
wire n_10206;
wire n_7844;
wire n_5207;
wire n_7934;
wire n_11281;
wire n_361;
wire n_2658;
wire n_12957;
wire n_5624;
wire n_10092;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_7009;
wire n_3376;
wire n_11772;
wire n_181;
wire n_9743;
wire n_9121;
wire n_7371;
wire n_13448;
wire n_1362;
wire n_11237;
wire n_14752;
wire n_9509;
wire n_3123;
wire n_5447;
wire n_12153;
wire n_2692;
wire n_12005;
wire n_683;
wire n_7463;
wire n_9621;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_10738;
wire n_4308;
wire n_5700;
wire n_11851;
wire n_5755;
wire n_9158;
wire n_2862;
wire n_4325;
wire n_14239;
wire n_14501;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_6889;
wire n_2749;
wire n_12586;
wire n_11993;
wire n_5962;
wire n_660;
wire n_464;
wire n_4413;
wire n_11131;
wire n_12221;
wire n_8627;
wire n_1210;
wire n_14318;
wire n_11432;
wire n_12302;
wire n_3307;
wire n_8945;
wire n_9142;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_13628;
wire n_2833;
wire n_9216;
wire n_9189;
wire n_6723;
wire n_7398;
wire n_1038;
wire n_3723;
wire n_7941;
wire n_4135;
wire n_9563;
wire n_12757;
wire n_13010;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_13251;
wire n_14738;
wire n_8858;
wire n_12107;
wire n_414;
wire n_571;
wire n_11738;
wire n_11595;
wire n_3880;
wire n_13521;
wire n_13504;
wire n_14404;
wire n_12695;
wire n_11512;
wire n_5801;
wire n_14163;
wire n_3904;
wire n_12349;
wire n_6054;
wire n_13703;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_14758;
wire n_13161;
wire n_7011;
wire n_10813;
wire n_3405;
wire n_2313;
wire n_14076;
wire n_10986;
wire n_11603;
wire n_6393;
wire n_14291;
wire n_14761;
wire n_12380;
wire n_7074;
wire n_10853;
wire n_8916;
wire n_10899;
wire n_11707;
wire n_11728;
wire n_613;
wire n_13352;
wire n_11521;
wire n_1022;
wire n_13309;
wire n_5465;
wire n_12577;
wire n_10575;
wire n_171;
wire n_8745;
wire n_3532;
wire n_5154;
wire n_14388;
wire n_5721;
wire n_2609;
wire n_8169;
wire n_6184;
wire n_11802;
wire n_8018;
wire n_1767;
wire n_9984;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_7083;
wire n_316;
wire n_1973;
wire n_1444;
wire n_820;
wire n_8260;
wire n_12723;
wire n_10334;
wire n_14153;
wire n_12135;
wire n_254;
wire n_2882;
wire n_14674;
wire n_7143;
wire n_2303;
wire n_7701;
wire n_11688;
wire n_13484;
wire n_8688;
wire n_9794;
wire n_7969;
wire n_10726;
wire n_8279;
wire n_4384;
wire n_8793;
wire n_4639;
wire n_1664;
wire n_12864;
wire n_13486;
wire n_10388;
wire n_4577;
wire n_6312;
wire n_13478;
wire n_7683;
wire n_9550;
wire n_13108;
wire n_532;
wire n_11042;
wire n_2154;
wire n_12570;
wire n_14124;
wire n_10510;
wire n_14344;
wire n_7669;
wire n_1986;
wire n_8298;
wire n_6711;
wire n_2624;
wire n_11696;
wire n_6818;
wire n_6438;
wire n_2054;
wire n_1857;
wire n_11761;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_10635;
wire n_11681;
wire n_1552;
wire n_2938;
wire n_7209;
wire n_2498;
wire n_13429;
wire n_6193;
wire n_3992;
wire n_13897;
wire n_8023;
wire n_9319;
wire n_7330;
wire n_6007;
wire n_13374;
wire n_621;
wire n_13182;
wire n_10852;
wire n_6734;
wire n_6535;
wire n_13789;
wire n_8053;
wire n_11407;
wire n_8059;
wire n_1772;
wire n_9871;
wire n_14354;
wire n_6879;
wire n_9562;
wire n_9896;
wire n_9612;
wire n_493;
wire n_1311;
wire n_3106;
wire n_6208;
wire n_7190;
wire n_9698;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_7692;
wire n_697;
wire n_9528;
wire n_10241;
wire n_4620;
wire n_6255;
wire n_6457;
wire n_13690;
wire n_14016;
wire n_9272;
wire n_13055;
wire n_14379;
wire n_9955;
wire n_5397;
wire n_9645;
wire n_4924;
wire n_4044;
wire n_8372;
wire n_6270;
wire n_14283;
wire n_2305;
wire n_8737;
wire n_9731;
wire n_10026;
wire n_5996;
wire n_880;
wire n_13577;
wire n_5566;
wire n_9697;
wire n_3304;
wire n_7288;
wire n_10772;
wire n_4388;
wire n_13098;
wire n_10901;
wire n_7362;
wire n_7237;
wire n_7082;
wire n_8988;
wire n_3247;
wire n_10664;
wire n_7131;
wire n_6276;
wire n_739;
wire n_1028;
wire n_12328;
wire n_13839;
wire n_9642;
wire n_530;
wire n_8723;
wire n_11189;
wire n_12559;
wire n_9929;
wire n_9050;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_12056;
wire n_13898;
wire n_7042;
wire n_9859;
wire n_8419;
wire n_2809;
wire n_10767;
wire n_10320;
wire n_5652;
wire n_13380;
wire n_8893;
wire n_975;
wire n_1645;
wire n_5805;
wire n_7304;
wire n_932;
wire n_11910;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_12109;
wire n_2910;
wire n_14457;
wire n_2503;
wire n_9531;
wire n_10521;
wire n_3785;
wire n_5492;
wire n_8077;
wire n_11242;
wire n_2465;
wire n_5501;
wire n_12917;
wire n_14711;
wire n_6934;
wire n_13188;
wire n_14179;
wire n_13362;
wire n_7386;
wire n_2972;
wire n_7391;
wire n_4401;
wire n_11361;
wire n_2586;
wire n_2989;
wire n_7754;
wire n_11894;
wire n_3178;
wire n_12058;
wire n_8826;
wire n_268;
wire n_13819;
wire n_7023;
wire n_10872;
wire n_13990;
wire n_2251;
wire n_9732;
wire n_5842;
wire n_5758;
wire n_12083;
wire n_9685;
wire n_12529;
wire n_3100;
wire n_3721;
wire n_10374;
wire n_11253;
wire n_13983;
wire n_12045;
wire n_13193;
wire n_7404;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_10345;
wire n_8959;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_12471;
wire n_4973;
wire n_13781;
wire n_13802;
wire n_7981;
wire n_4792;
wire n_1601;
wire n_13037;
wire n_3537;
wire n_4402;
wire n_14252;
wire n_14736;
wire n_12188;
wire n_191;
wire n_2487;
wire n_5473;
wire n_12575;
wire n_1834;
wire n_10601;
wire n_14698;
wire n_11623;
wire n_8712;
wire n_12473;
wire n_10372;
wire n_1011;
wire n_2534;
wire n_6352;
wire n_11124;
wire n_14295;
wire n_2941;
wire n_4286;
wire n_9378;
wire n_3638;
wire n_6211;
wire n_10448;
wire n_8109;
wire n_10301;
wire n_11977;
wire n_3576;
wire n_10074;
wire n_12040;
wire n_14025;
wire n_13127;
wire n_9389;
wire n_12598;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_10001;
wire n_13561;
wire n_7378;
wire n_9623;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_7877;
wire n_14336;
wire n_11351;
wire n_7787;
wire n_7836;
wire n_8515;
wire n_8725;
wire n_12626;
wire n_11094;
wire n_10960;
wire n_10712;
wire n_8007;
wire n_13911;
wire n_14313;
wire n_2387;
wire n_4318;
wire n_332;
wire n_13961;
wire n_13343;
wire n_12546;
wire n_8910;
wire n_5227;
wire n_14091;
wire n_830;
wire n_10100;
wire n_5902;
wire n_987;
wire n_2510;
wire n_9164;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_11366;
wire n_2793;
wire n_5282;
wire n_9387;
wire n_8301;
wire n_7871;
wire n_6764;
wire n_14512;
wire n_541;
wire n_499;
wire n_13539;
wire n_10162;
wire n_2639;
wire n_9840;
wire n_7016;
wire n_4738;
wire n_12100;
wire n_2603;
wire n_8892;
wire n_11399;
wire n_9637;
wire n_5386;
wire n_1167;
wire n_12676;
wire n_4554;
wire n_7571;
wire n_8252;
wire n_4526;
wire n_4105;
wire n_10535;
wire n_10674;
wire n_13584;
wire n_6215;
wire n_969;
wire n_3663;
wire n_9491;
wire n_1663;
wire n_7563;
wire n_6955;
wire n_10774;
wire n_10337;
wire n_5952;
wire n_7180;
wire n_13107;
wire n_10407;
wire n_14655;
wire n_10577;
wire n_2086;
wire n_14481;
wire n_13778;
wire n_1926;
wire n_8972;
wire n_14531;
wire n_8494;
wire n_12999;
wire n_14709;
wire n_10264;
wire n_6569;
wire n_1630;
wire n_7919;
wire n_13740;
wire n_9992;
wire n_14606;
wire n_14089;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_8278;
wire n_443;
wire n_3431;
wire n_11549;
wire n_8180;
wire n_14437;
wire n_12362;
wire n_3355;
wire n_7031;
wire n_13913;
wire n_1738;
wire n_13367;
wire n_5716;
wire n_10313;
wire n_10843;
wire n_12983;
wire n_14003;
wire n_8941;
wire n_10771;
wire n_8891;
wire n_406;
wire n_3897;
wire n_7103;
wire n_12360;
wire n_139;
wire n_13570;
wire n_6605;
wire n_10724;
wire n_1735;
wire n_391;
wire n_5888;
wire n_9266;
wire n_4005;
wire n_14409;
wire n_8270;
wire n_8231;
wire n_4181;
wire n_2543;
wire n_2597;
wire n_1077;
wire n_2321;
wire n_11983;
wire n_6832;
wire n_12313;
wire n_12604;
wire n_5980;
wire n_8683;
wire n_956;
wire n_9391;
wire n_765;
wire n_4092;
wire n_12558;
wire n_10445;
wire n_4875;
wire n_7771;
wire n_8903;
wire n_4255;
wire n_13284;
wire n_2758;
wire n_385;
wire n_6544;
wire n_8810;
wire n_12596;
wire n_6469;
wire n_12840;
wire n_11119;
wire n_1271;
wire n_12696;
wire n_5036;
wire n_6332;
wire n_10863;
wire n_10958;
wire n_2186;
wire n_11215;
wire n_13730;
wire n_5790;
wire n_399;
wire n_7130;
wire n_10174;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_13960;
wire n_8932;
wire n_6310;
wire n_8264;
wire n_12435;
wire n_2471;
wire n_9695;
wire n_7134;
wire n_3042;
wire n_8288;
wire n_13411;
wire n_1067;
wire n_11954;
wire n_14629;
wire n_14778;
wire n_1323;
wire n_11526;
wire n_13438;
wire n_14010;
wire n_11591;
wire n_10403;
wire n_1937;
wire n_11972;
wire n_4142;
wire n_5118;
wire n_9834;
wire n_900;
wire n_5485;
wire n_9901;
wire n_5525;
wire n_7102;
wire n_10015;
wire n_10076;
wire n_6259;
wire n_3004;
wire n_14432;
wire n_1551;
wire n_5271;
wire n_4849;
wire n_13410;
wire n_2039;
wire n_7133;
wire n_9800;
wire n_1285;
wire n_10745;
wire n_193;
wire n_733;
wire n_761;
wire n_3838;
wire n_6651;
wire n_6289;
wire n_9255;
wire n_8882;
wire n_14308;
wire n_12460;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_12733;
wire n_8388;
wire n_5445;
wire n_2734;
wire n_8067;
wire n_13600;
wire n_8385;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_8670;
wire n_4504;
wire n_10460;
wire n_14299;
wire n_14215;
wire n_3598;
wire n_4917;
wire n_7813;
wire n_7706;
wire n_8142;
wire n_13332;
wire n_14265;
wire n_13942;
wire n_2420;
wire n_7992;
wire n_9085;
wire n_7643;
wire n_11204;
wire n_153;
wire n_648;
wire n_6836;
wire n_12939;
wire n_3273;
wire n_9120;
wire n_2918;
wire n_6595;
wire n_10415;
wire n_11302;
wire n_835;
wire n_9899;
wire n_12374;
wire n_9136;
wire n_12261;
wire n_6186;
wire n_11561;
wire n_10227;
wire n_1865;
wire n_2641;
wire n_13490;
wire n_2463;
wire n_14198;
wire n_2580;
wire n_401;
wire n_7628;
wire n_1792;
wire n_13381;
wire n_5628;
wire n_504;
wire n_5245;
wire n_2062;
wire n_483;
wire n_4489;
wire n_9436;
wire n_14013;
wire n_11385;
wire n_822;
wire n_1459;
wire n_2153;
wire n_12065;
wire n_13204;
wire n_5329;
wire n_12275;
wire n_8224;
wire n_5472;
wire n_9042;
wire n_10884;
wire n_6035;
wire n_13375;
wire n_839;
wire n_1754;
wire n_7236;
wire n_9570;
wire n_4833;
wire n_3394;
wire n_9239;
wire n_6405;
wire n_8345;
wire n_11054;
wire n_11777;
wire n_9644;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_9343;
wire n_8614;
wire n_8242;
wire n_6786;
wire n_4564;
wire n_8299;
wire n_1848;
wire n_9131;
wire n_1172;
wire n_13286;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_9060;
wire n_9792;
wire n_3581;
wire n_8110;
wire n_5072;
wire n_8529;
wire n_3778;
wire n_14204;
wire n_13384;
wire n_11325;
wire n_10801;
wire n_6769;
wire n_10325;
wire n_13013;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_8951;
wire n_2260;
wire n_323;
wire n_1660;
wire n_1315;
wire n_11217;
wire n_4080;
wire n_2206;
wire n_997;
wire n_635;
wire n_13582;
wire n_12752;
wire n_10327;
wire n_8700;
wire n_6766;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_14157;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_11651;
wire n_6232;
wire n_2347;
wire n_13255;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_7802;
wire n_7519;
wire n_10505;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_12979;
wire n_14140;
wire n_2362;
wire n_7457;
wire n_14723;
wire n_11196;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_11672;
wire n_11557;
wire n_9982;
wire n_2422;
wire n_11552;
wire n_6416;
wire n_654;
wire n_13682;
wire n_2933;
wire n_8468;
wire n_9031;
wire n_12715;
wire n_12910;
wire n_7515;
wire n_3387;
wire n_7639;
wire n_11084;
wire n_12787;
wire n_8933;
wire n_6214;
wire n_3952;
wire n_9006;
wire n_8636;
wire n_10408;
wire n_11442;
wire n_9221;
wire n_13424;
wire n_4365;
wire n_3584;
wire n_14102;
wire n_4349;
wire n_3446;
wire n_10514;
wire n_1059;
wire n_7049;
wire n_7884;
wire n_6945;
wire n_8378;
wire n_6143;
wire n_14603;
wire n_2736;
wire n_6491;
wire n_10091;
wire n_7592;
wire n_7749;
wire n_11195;
wire n_3825;
wire n_4198;
wire n_10562;
wire n_7172;
wire n_539;
wire n_10586;
wire n_10893;
wire n_8283;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_7914;
wire n_1866;
wire n_8860;
wire n_2664;
wire n_12401;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_14104;
wire n_4390;
wire n_459;
wire n_10593;
wire n_13304;
wire n_1782;
wire n_11517;
wire n_7892;
wire n_1558;
wire n_4107;
wire n_12722;
wire n_13716;
wire n_2519;
wire n_9523;
wire n_10821;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_7325;
wire n_11918;
wire n_14561;
wire n_13460;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_723;
wire n_1393;
wire n_7674;
wire n_8686;
wire n_13590;
wire n_12712;
wire n_10961;
wire n_6175;
wire n_6445;
wire n_9829;
wire n_8563;
wire n_11077;
wire n_4571;
wire n_13914;
wire n_3137;
wire n_2544;
wire n_11579;
wire n_809;
wire n_10197;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_8493;
wire n_6198;
wire n_5172;
wire n_14119;
wire n_13670;
wire n_13148;
wire n_10950;
wire n_881;
wire n_1019;
wire n_1477;
wire n_9411;
wire n_6499;
wire n_1982;
wire n_12209;
wire n_7983;
wire n_641;
wire n_5311;
wire n_8765;
wire n_14168;
wire n_14494;
wire n_910;
wire n_13452;
wire n_290;
wire n_14506;
wire n_5164;
wire n_11640;
wire n_13688;
wire n_4964;
wire n_10180;
wire n_9153;
wire n_4700;
wire n_6842;
wire n_4002;
wire n_217;
wire n_10079;
wire n_7361;
wire n_1114;
wire n_11656;
wire n_1742;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_201;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_11845;
wire n_1199;
wire n_11679;
wire n_14007;
wire n_13671;
wire n_1273;
wire n_2982;
wire n_8653;
wire n_5495;
wire n_6281;
wire n_13005;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_13313;
wire n_5547;
wire n_4693;
wire n_10361;
wire n_14154;
wire n_11635;
wire n_8601;
wire n_1043;
wire n_9675;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_255;
wire n_2869;
wire n_8333;
wire n_9097;
wire n_9571;
wire n_12323;
wire n_12835;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_10075;
wire n_11572;
wire n_9789;
wire n_2674;
wire n_13387;
wire n_13068;
wire n_5820;
wire n_11529;
wire n_9925;
wire n_1737;
wire n_7309;
wire n_7119;
wire n_1613;
wire n_14426;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_7696;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_13173;
wire n_10012;
wire n_3902;
wire n_14351;
wire n_196;
wire n_12873;
wire n_12830;
wire n_12015;
wire n_12348;
wire n_12767;
wire n_3244;
wire n_10939;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_10008;
wire n_11384;
wire n_14382;
wire n_9511;
wire n_9795;
wire n_3196;
wire n_231;
wire n_11134;
wire n_8708;
wire n_10503;
wire n_5964;
wire n_2673;
wire n_10111;
wire n_10982;
wire n_10798;
wire n_11630;
wire n_4678;
wire n_664;
wire n_1591;
wire n_12867;
wire n_13479;
wire n_13710;
wire n_5301;
wire n_13203;
wire n_13263;
wire n_14700;
wire n_5126;
wire n_13211;
wire n_8659;
wire n_8759;
wire n_6732;
wire n_2548;
wire n_3488;
wire n_9622;
wire n_2381;
wire n_12198;
wire n_9761;
wire n_14707;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_544;
wire n_7646;
wire n_14249;
wire n_9954;
wire n_14530;
wire n_3779;
wire n_599;
wire n_13848;
wire n_12617;
wire n_6982;
wire n_537;
wire n_1063;
wire n_7291;
wire n_10669;
wire n_8790;
wire n_991;
wire n_2275;
wire n_13052;
wire n_7668;
wire n_7435;
wire n_4606;
wire n_8832;
wire n_13282;
wire n_8305;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_8453;
wire n_6560;
wire n_6634;
wire n_14275;
wire n_5348;
wire n_583;
wire n_12666;
wire n_9847;
wire n_13818;
wire n_1000;
wire n_313;
wire n_4868;
wire n_7017;
wire n_13846;
wire n_378;
wire n_12845;
wire n_11617;
wire n_4072;
wire n_7848;
wire n_2792;
wire n_13312;
wire n_4465;
wire n_9640;
wire n_8127;
wire n_13565;
wire n_2596;
wire n_5217;
wire n_8337;
wire n_9115;
wire n_3986;
wire n_7861;
wire n_3725;
wire n_12047;
wire n_5558;
wire n_10190;
wire n_12411;
wire n_9534;
wire n_472;
wire n_4026;
wire n_13788;
wire n_4245;
wire n_11422;
wire n_5520;
wire n_2524;
wire n_7889;
wire n_13295;
wire n_208;
wire n_3894;
wire n_1702;
wire n_12594;
wire n_10542;
wire n_14349;
wire n_5909;
wire n_4852;
wire n_275;
wire n_7554;
wire n_3202;
wire n_11289;
wire n_8508;
wire n_4290;
wire n_4945;
wire n_11376;
wire n_5750;
wire n_7648;
wire n_8968;
wire n_147;
wire n_1232;
wire n_1211;
wire n_996;
wire n_10752;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_11157;
wire n_2318;
wire n_14718;
wire n_866;
wire n_10868;
wire n_11013;
wire n_2819;
wire n_1722;
wire n_9594;
wire n_11017;
wire n_2229;
wire n_7653;
wire n_11765;
wire n_6400;
wire n_12885;
wire n_1644;
wire n_11307;
wire n_7846;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_8347;
wire n_2255;
wire n_5554;
wire n_9503;
wire n_1252;
wire n_12811;
wire n_3045;
wire n_9919;
wire n_250;
wire n_13346;
wire n_773;
wire n_13331;
wire n_5135;
wire n_7551;
wire n_11793;
wire n_11574;
wire n_4599;
wire n_13307;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_10017;
wire n_13574;
wire n_718;
wire n_12073;
wire n_1434;
wire n_8093;
wire n_9385;
wire n_8899;
wire n_12913;
wire n_1905;
wire n_13027;
wire n_1569;
wire n_14563;
wire n_5448;
wire n_2573;
wire n_6480;
wire n_7737;
wire n_5837;
wire n_11836;
wire n_2336;
wire n_5412;
wire n_523;
wire n_1662;
wire n_8481;
wire n_14169;
wire n_3249;
wire n_3483;
wire n_6851;
wire n_6621;
wire n_4046;
wire n_11747;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_7606;
wire n_9963;
wire n_7420;
wire n_10572;
wire n_11193;
wire n_9885;
wire n_8115;
wire n_4869;
wire n_13939;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_11670;
wire n_1244;
wire n_1796;
wire n_14042;
wire n_484;
wire n_10642;
wire n_2719;
wire n_10115;
wire n_10517;
wire n_14429;
wire n_14098;
wire n_13289;
wire n_10247;
wire n_2876;
wire n_13851;
wire n_13852;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_12451;
wire n_12585;
wire n_12029;
wire n_12963;
wire n_13616;
wire n_6226;
wire n_14490;
wire n_9827;
wire n_1574;
wire n_12169;
wire n_14748;
wire n_3033;
wire n_12801;
wire n_893;
wire n_9182;
wire n_10620;
wire n_1582;
wire n_8182;
wire n_9426;
wire n_9293;
wire n_1981;
wire n_2824;
wire n_10065;
wire n_7973;
wire n_7545;
wire n_5327;
wire n_4417;
wire n_796;
wire n_11762;
wire n_14030;
wire n_14500;
wire n_531;
wire n_1374;
wire n_2089;
wire n_7896;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_9581;
wire n_8629;
wire n_12657;
wire n_5900;
wire n_8186;
wire n_7319;
wire n_1486;
wire n_11758;
wire n_3619;
wire n_6158;
wire n_13366;
wire n_9400;
wire n_4013;
wire n_10744;
wire n_3434;
wire n_9246;
wire n_4342;
wire n_691;
wire n_6819;
wire n_4903;
wire n_6122;
wire n_2131;
wire n_3853;
wire n_8233;
wire n_4382;
wire n_2509;
wire n_423;
wire n_4085;
wire n_6898;
wire n_14734;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_9445;
wire n_8282;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5432;
wire n_7516;
wire n_5851;
wire n_6928;
wire n_6317;
wire n_10609;
wire n_13860;
wire n_11958;
wire n_6707;
wire n_10009;
wire n_13847;
wire n_7244;
wire n_187;
wire n_11314;
wire n_1463;
wire n_4626;
wire n_12210;
wire n_10072;
wire n_12443;
wire n_12699;
wire n_7625;
wire n_8750;
wire n_10130;
wire n_4997;
wire n_8183;
wire n_13657;
wire n_5065;
wire n_9104;
wire n_13450;
wire n_6806;
wire n_924;
wire n_10956;
wire n_7991;
wire n_781;
wire n_8637;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_9542;
wire n_11490;
wire n_11515;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_8792;
wire n_6835;
wire n_7286;
wire n_2436;
wire n_3517;
wire n_13610;
wire n_6269;
wire n_7857;
wire n_13871;
wire n_7970;
wire n_9302;
wire n_1706;
wire n_2461;
wire n_10829;
wire n_8258;
wire n_3719;
wire n_7154;
wire n_11356;
wire n_524;
wire n_12781;
wire n_1214;
wire n_634;
wire n_10506;
wire n_3526;
wire n_3888;
wire n_9960;
wire n_12573;
wire n_13326;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_8416;
wire n_8390;
wire n_13881;
wire n_11678;
wire n_12744;
wire n_6088;
wire n_10236;
wire n_11374;
wire n_14519;
wire n_1181;
wire n_1999;
wire n_11176;
wire n_7194;
wire n_4841;
wire n_11402;
wire n_4683;
wire n_5173;
wire n_11162;
wire n_2873;
wire n_10002;
wire n_8696;
wire n_9185;
wire n_9601;
wire n_13137;
wire n_2084;
wire n_13226;
wire n_3330;
wire n_3514;
wire n_11771;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_7175;
wire n_13431;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_7163;
wire n_5855;
wire n_14402;
wire n_14507;
wire n_14020;
wire n_3797;
wire n_1836;
wire n_13552;
wire n_13164;
wire n_7027;
wire n_3416;
wire n_8552;
wire n_12006;
wire n_4600;
wire n_5861;
wire n_1453;
wire n_6964;
wire n_3943;
wire n_10855;
wire n_3145;
wire n_14389;
wire n_7964;
wire n_5749;
wire n_6320;
wire n_9403;
wire n_14558;
wire n_11322;
wire n_6316;
wire n_8619;
wire n_419;
wire n_11484;
wire n_7068;
wire n_9972;
wire n_11711;
wire n_13227;
wire n_2908;
wire n_8594;
wire n_9878;
wire n_14541;
wire n_10139;
wire n_14183;
wire n_270;
wire n_4106;
wire n_9541;
wire n_10941;
wire n_14689;
wire n_285;
wire n_2156;
wire n_12548;
wire n_1184;
wire n_202;
wire n_8162;
wire n_9735;
wire n_754;
wire n_9576;
wire n_14528;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_7327;
wire n_12727;
wire n_1277;
wire n_1746;
wire n_12240;
wire n_13045;
wire n_6610;
wire n_13620;
wire n_1062;
wire n_5998;
wire n_8318;
wire n_14742;
wire n_4702;
wire n_5102;
wire n_9974;
wire n_4954;
wire n_740;
wire n_10992;
wire n_167;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_8425;
wire n_6752;
wire n_13001;
wire n_6959;
wire n_9704;
wire n_6250;
wire n_13919;
wire n_11392;
wire n_12372;
wire n_3283;
wire n_11803;
wire n_259;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_11912;
wire n_13862;
wire n_13784;
wire n_7864;
wire n_11139;
wire n_3451;
wire n_10650;
wire n_8051;
wire n_4734;
wire n_11021;
wire n_6675;
wire n_7955;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_9039;
wire n_12914;
wire n_7384;
wire n_12844;
wire n_267;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_1988;
wire n_12952;
wire n_5678;
wire n_6561;
wire n_11379;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_13271;
wire n_7512;
wire n_1718;
wire n_7814;
wire n_12276;
wire n_12096;
wire n_8389;
wire n_4515;
wire n_10417;
wire n_2149;
wire n_2277;
wire n_200;
wire n_10029;
wire n_12150;
wire n_14271;
wire n_13595;
wire n_2539;
wire n_8620;
wire n_10125;
wire n_6850;
wire n_5555;
wire n_13757;
wire n_2078;
wire n_8886;
wire n_1145;
wire n_4809;
wire n_7152;
wire n_14770;
wire n_787;
wire n_4012;
wire n_10253;
wire n_11899;
wire n_1195;
wire n_13761;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_13136;
wire n_13190;
wire n_6823;
wire n_10693;
wire n_3606;
wire n_14461;
wire n_7062;
wire n_7090;
wire n_12449;
wire n_8202;
wire n_13633;
wire n_2232;
wire n_11966;
wire n_1847;
wire n_14205;
wire n_5815;
wire n_4320;
wire n_12118;
wire n_10599;
wire n_5084;
wire n_7223;
wire n_14266;
wire n_12770;
wire n_5251;
wire n_1314;
wire n_8755;
wire n_13174;
wire n_1512;
wire n_8668;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_10977;
wire n_13528;
wire n_2192;
wire n_6796;
wire n_8979;
wire n_5407;
wire n_2988;
wire n_12814;
wire n_11553;
wire n_4560;
wire n_14064;
wire n_14322;
wire n_13220;
wire n_12009;
wire n_14466;
wire n_13456;
wire n_13916;
wire n_7761;
wire n_10947;
wire n_8141;
wire n_10386;
wire n_3793;
wire n_3230;
wire n_859;
wire n_8199;
wire n_5042;
wire n_12826;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_10267;
wire n_6090;
wire n_693;
wire n_5368;
wire n_929;
wire n_10401;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_9908;
wire n_11127;
wire n_8004;
wire n_11926;
wire n_8383;
wire n_14763;
wire n_3607;
wire n_1637;
wire n_9688;
wire n_9864;
wire n_2427;
wire n_12144;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_7388;
wire n_1751;
wire n_7056;
wire n_10428;
wire n_14585;
wire n_10212;
wire n_7437;
wire n_11460;
wire n_6489;
wire n_11486;
wire n_9023;
wire n_5310;
wire n_2769;
wire n_8895;
wire n_438;
wire n_8680;
wire n_1548;
wire n_14208;
wire n_4987;
wire n_6714;
wire n_8394;
wire n_440;
wire n_7849;
wire n_10539;
wire n_14152;
wire n_7726;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_7417;
wire n_2739;
wire n_12937;
wire n_3962;
wire n_11148;
wire n_4988;
wire n_7446;
wire n_6038;
wire n_10728;
wire n_12312;
wire n_2902;
wire n_6030;
wire n_6620;
wire n_4360;
wire n_1544;
wire n_6245;
wire n_6791;
wire n_4540;
wire n_9220;
wire n_13929;
wire n_6821;
wire n_9317;
wire n_12580;
wire n_13965;
wire n_2094;
wire n_13796;
wire n_5588;
wire n_3854;
wire n_8198;
wire n_9993;
wire n_1354;
wire n_10879;
wire n_13474;
wire n_8665;
wire n_12393;
wire n_6583;
wire n_10545;
wire n_2349;
wire n_3652;
wire n_12201;
wire n_7859;
wire n_3449;
wire n_13240;
wire n_1021;
wire n_13187;
wire n_13594;
wire n_3089;
wire n_4854;
wire n_9561;
wire n_491;
wire n_10516;
wire n_14640;
wire n_9444;
wire n_1595;
wire n_10497;
wire n_1142;
wire n_8017;
wire n_11675;
wire n_5477;
wire n_260;
wire n_2727;
wire n_942;
wire n_10705;
wire n_7523;
wire n_12082;
wire n_13966;
wire n_11032;
wire n_5234;
wire n_14035;
wire n_12322;
wire n_1416;
wire n_6890;
wire n_9184;
wire n_10432;
wire n_11454;
wire n_7559;
wire n_14345;
wire n_9037;
wire n_7576;
wire n_6988;
wire n_10779;
wire n_8303;
wire n_11554;
wire n_1599;
wire n_5871;
wire n_11988;
wire n_13981;
wire n_4747;
wire n_14647;
wire n_8000;
wire n_11197;
wire n_14286;
wire n_3472;
wire n_14686;
wire n_2527;
wire n_6052;
wire n_7769;
wire n_11416;
wire n_9505;
wire n_9193;
wire n_14360;
wire n_7257;
wire n_3126;
wire n_12986;
wire n_2759;
wire n_6973;
wire n_10869;
wire n_8852;
wire n_5007;
wire n_8709;
wire n_4881;
wire n_10314;
wire n_2038;
wire n_10504;
wire n_6488;
wire n_4495;
wire n_3958;
wire n_10687;
wire n_13691;
wire n_4737;
wire n_1838;
wire n_9218;
wire n_9755;
wire n_4357;
wire n_11341;
wire n_7729;
wire n_2806;
wire n_4502;
wire n_11045;
wire n_287;
wire n_3191;
wire n_1716;
wire n_12373;
wire n_302;
wire n_7005;
wire n_12741;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_8782;
wire n_7081;
wire n_10882;
wire n_7742;
wire n_5253;
wire n_10293;
wire n_3588;
wire n_355;
wire n_6280;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_9506;
wire n_9162;
wire n_13629;
wire n_3095;
wire n_947;
wire n_7341;
wire n_5792;
wire n_13155;
wire n_14581;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_11569;
wire n_468;
wire n_13152;
wire n_10256;
wire n_182;
wire n_696;
wire n_1442;
wire n_4775;
wire n_6256;
wire n_482;
wire n_2620;
wire n_1833;
wire n_8716;
wire n_12412;
wire n_1691;
wire n_8250;
wire n_12677;
wire n_7264;
wire n_7842;
wire n_14315;
wire n_12181;
wire n_12833;
wire n_2549;
wire n_2499;
wire n_6648;
wire n_9415;
wire n_10298;
wire n_12115;
wire n_12631;
wire n_7492;
wire n_13194;
wire n_13546;
wire n_804;
wire n_6649;
wire n_8714;
wire n_1656;
wire n_8357;
wire n_12567;
wire n_1382;
wire n_3093;
wire n_12175;
wire n_2970;
wire n_6910;
wire n_9990;
wire n_3885;
wire n_955;
wire n_8466;
wire n_4264;
wire n_5954;
wire n_9015;
wire n_10326;
wire n_2166;
wire n_13446;
wire n_10235;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_514;
wire n_6431;
wire n_418;
wire n_8589;
wire n_12754;
wire n_3250;
wire n_4223;
wire n_14141;
wire n_12455;
wire n_3538;
wire n_13363;
wire n_3915;
wire n_11990;
wire n_8266;
wire n_3839;
wire n_8587;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_10725;
wire n_10274;
wire n_13728;
wire n_13601;
wire n_3875;
wire n_4029;
wire n_8876;
wire n_11541;
wire n_9214;
wire n_14780;
wire n_4206;
wire n_12340;
wire n_2415;
wire n_4099;
wire n_10799;
wire n_8922;
wire n_11680;
wire n_10090;
wire n_3120;
wire n_6512;
wire n_12686;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_9070;
wire n_8498;
wire n_4794;
wire n_9933;
wire n_4843;
wire n_12734;
wire n_669;
wire n_5580;
wire n_5215;
wire n_337;
wire n_437;
wire n_12331;
wire n_3937;
wire n_4763;
wire n_10874;
wire n_9339;
wire n_11596;
wire n_1418;
wire n_9991;
wire n_12880;
wire n_9486;
wire n_8457;
wire n_6243;
wire n_14113;
wire n_5795;
wire n_10763;
wire n_5715;
wire n_4170;
wire n_10266;
wire n_12184;
wire n_12425;
wire n_8267;
wire n_5561;
wire n_2462;
wire n_7051;
wire n_13918;
wire n_11180;
wire n_6773;
wire n_10290;
wire n_2155;
wire n_6231;
wire n_12472;
wire n_615;
wire n_13048;
wire n_12266;
wire n_7503;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_12432;
wire n_517;
wire n_8124;
wire n_3604;
wire n_8545;
wire n_5430;
wire n_8526;
wire n_6041;
wire n_824;
wire n_12300;
wire n_159;
wire n_13593;
wire n_8319;
wire n_7997;
wire n_12527;
wire n_5659;
wire n_11839;
wire n_9279;
wire n_6859;
wire n_7716;
wire n_4272;
wire n_10732;
wire n_5195;
wire n_12110;
wire n_13744;
wire n_3176;
wire n_9790;
wire n_144;
wire n_11404;
wire n_3792;
wire n_7950;
wire n_11548;
wire n_6323;
wire n_13515;
wire n_5720;
wire n_4267;
wire n_8581;
wire n_12122;
wire n_10873;
wire n_8214;
wire n_7793;
wire n_9053;
wire n_8516;
wire n_2083;
wire n_815;
wire n_12310;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_470;
wire n_11343;
wire n_3021;
wire n_8989;
wire n_13028;
wire n_7746;
wire n_477;
wire n_11362;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_11007;
wire n_3950;
wire n_7570;
wire n_9650;
wire n_9880;
wire n_11497;
wire n_2898;
wire n_1825;
wire n_10720;
wire n_6912;
wire n_3567;
wire n_14574;
wire n_7425;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_14014;
wire n_12827;
wire n_14078;
wire n_10220;
wire n_9217;
wire n_9499;
wire n_5783;
wire n_7829;
wire n_6837;
wire n_13467;
wire n_13245;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_10081;
wire n_12804;
wire n_3812;
wire n_3127;
wire n_9282;
wire n_1731;
wire n_799;
wire n_7894;
wire n_10145;
wire n_1147;
wire n_11347;
wire n_12892;
wire n_7957;
wire n_8262;
wire n_2378;
wire n_10167;
wire n_5530;
wire n_12656;
wire n_6718;
wire n_8289;
wire n_965;
wire n_13804;
wire n_5809;
wire n_10447;
wire n_12418;
wire n_934;
wire n_2213;
wire n_7531;
wire n_12448;
wire n_6410;
wire n_7121;
wire n_12219;
wire n_12729;
wire n_356;
wire n_13549;
wire n_13921;
wire n_6473;
wire n_8087;
wire n_4056;
wire n_10238;
wire n_13345;
wire n_4806;
wire n_11029;
wire n_7961;
wire n_1674;
wire n_9920;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_7687;
wire n_9948;
wire n_5299;
wire n_4462;
wire n_13216;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_11226;
wire n_2142;
wire n_8863;
wire n_9371;
wire n_4517;
wire n_2896;
wire n_8701;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_13036;
wire n_1042;
wire n_3170;
wire n_9237;
wire n_2311;
wire n_13398;
wire n_6857;
wire n_8705;
wire n_14148;
wire n_1455;
wire n_2287;
wire n_9815;
wire n_836;
wire n_3415;
wire n_10292;
wire n_12644;
wire n_6975;
wire n_10820;
wire n_7763;
wire n_13258;
wire n_3464;
wire n_6646;
wire n_3414;
wire n_6290;
wire n_205;
wire n_7703;
wire n_11760;
wire n_13827;
wire n_7928;
wire n_4234;
wire n_10395;
wire n_760;
wire n_1483;
wire n_12576;
wire n_10168;
wire n_14350;
wire n_1363;
wire n_8722;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_11664;
wire n_713;
wire n_3179;
wire n_598;
wire n_6622;
wire n_12187;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_7677;
wire n_5262;
wire n_7665;
wire n_13169;
wire n_14782;
wire n_3262;
wire n_10366;
wire n_5319;
wire n_10287;
wire n_14017;
wire n_927;
wire n_13940;
wire n_7469;
wire n_261;
wire n_3699;
wire n_10163;
wire n_6118;
wire n_706;
wire n_2120;
wire n_7125;
wire n_7856;
wire n_6028;
wire n_6663;
wire n_14145;
wire n_11006;
wire n_6532;
wire n_1419;
wire n_13406;
wire n_10431;
wire n_8622;
wire n_3816;
wire n_8099;
wire n_8729;
wire n_9479;
wire n_10876;
wire n_11485;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_9480;
wire n_12453;
wire n_12593;
wire n_4207;
wire n_11449;
wire n_8085;
wire n_2404;
wire n_2757;
wire n_2168;
wire n_4725;
wire n_9597;
wire n_10614;
wire n_10786;
wire n_13873;
wire n_13335;
wire n_14273;
wire n_348;
wire n_9173;
wire n_10352;
wire n_2312;
wire n_9641;
wire n_8947;
wire n_7203;
wire n_13714;
wire n_7797;
wire n_1826;
wire n_9983;
wire n_9267;
wire n_14565;
wire n_6556;
wire n_5943;
wire n_10039;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_13070;
wire n_6216;
wire n_13866;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_637;
wire n_7128;
wire n_9849;
wire n_11831;
wire n_5335;
wire n_1259;
wire n_11096;
wire n_11417;
wire n_8459;
wire n_2801;
wire n_7111;
wire n_1177;
wire n_4334;
wire n_8478;
wire n_5284;
wire n_12288;
wire n_8786;
wire n_9414;
wire n_4978;
wire n_11677;
wire n_13025;
wire n_14256;
wire n_5771;
wire n_3246;
wire n_9419;
wire n_3299;
wire n_8887;
wire n_980;
wire n_1618;
wire n_1869;
wire n_12091;
wire n_3623;
wire n_905;
wire n_2718;
wire n_11898;
wire n_4707;
wire n_14749;
wire n_2687;
wire n_8851;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_8540;
wire n_5516;
wire n_7284;
wire n_3615;
wire n_8276;
wire n_7057;
wire n_1802;
wire n_13457;
wire n_9823;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_9152;
wire n_8706;
wire n_3200;
wire n_6167;
wire n_12357;
wire n_3642;
wire n_145;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_11826;
wire n_7064;
wire n_12629;
wire n_8532;
wire n_9533;
wire n_10750;
wire n_5433;
wire n_3682;
wire n_11825;
wire n_5429;
wire n_7278;
wire n_12893;
wire n_9281;
wire n_9103;
wire n_9111;
wire n_6772;
wire n_7799;
wire n_7088;
wire n_9618;
wire n_10383;
wire n_5698;
wire n_10856;
wire n_5731;
wire n_14532;
wire n_14105;
wire n_10883;
wire n_12935;
wire n_8871;
wire n_4007;
wire n_1456;
wire n_9065;
wire n_8433;
wire n_10429;
wire n_14627;
wire n_14463;
wire n_1879;
wire n_14735;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_12732;
wire n_7048;
wire n_7979;
wire n_12569;
wire n_9674;
wire n_6617;
wire n_553;
wire n_7725;
wire n_13547;
wire n_814;
wire n_578;
wire n_10859;
wire n_5120;
wire n_3572;
wire n_8371;
wire n_2975;
wire n_2399;
wire n_8547;
wire n_11538;
wire n_10815;
wire n_1134;
wire n_11008;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_8467;
wire n_12980;
wire n_647;
wire n_11093;
wire n_11585;
wire n_2027;
wire n_2932;
wire n_8409;
wire n_6217;
wire n_600;
wire n_3118;
wire n_10303;
wire n_9157;
wire n_11616;
wire n_5560;
wire n_9170;
wire n_4441;
wire n_10424;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_502;
wire n_8640;
wire n_11001;
wire n_6777;
wire n_10196;
wire n_6742;
wire n_1467;
wire n_7447;
wire n_5209;
wire n_10684;
wire n_247;
wire n_13154;
wire n_6307;
wire n_5704;
wire n_14129;
wire n_4889;
wire n_2159;
wire n_4458;
wire n_8431;
wire n_14547;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_13280;
wire n_3618;
wire n_5916;
wire n_8415;
wire n_10184;
wire n_3705;
wire n_3022;
wire n_13904;
wire n_10421;
wire n_13944;
wire n_13359;
wire n_1709;
wire n_6479;
wire n_11472;
wire n_14376;
wire n_13855;
wire n_13073;
wire n_5099;
wire n_11063;
wire n_681;
wire n_3286;
wire n_5781;
wire n_11179;
wire n_5619;
wire n_2023;
wire n_14777;
wire n_9416;
wire n_11885;
wire n_3974;
wire n_9368;
wire n_7365;
wire n_3443;
wire n_8329;
wire n_13083;
wire n_14201;
wire n_2599;
wire n_3988;
wire n_7792;
wire n_8089;
wire n_9208;
wire n_11657;
wire n_13124;
wire n_9223;
wire n_6370;
wire n_5022;
wire n_2075;
wire n_13771;
wire n_1726;
wire n_10329;
wire n_10924;
wire n_13845;
wire n_11921;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_14224;
wire n_10285;
wire n_7275;
wire n_5353;
wire n_4771;
wire n_12099;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_1098;
wire n_9781;
wire n_3009;
wire n_13609;
wire n_13572;
wire n_13817;
wire n_8633;
wire n_12897;
wire n_777;
wire n_7095;
wire n_7390;
wire n_9392;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_9422;
wire n_920;
wire n_8541;
wire n_10084;
wire n_12924;
wire n_8762;
wire n_14162;
wire n_12619;
wire n_12541;
wire n_3951;
wire n_5518;
wire n_9970;
wire n_3035;
wire n_13428;
wire n_4261;
wire n_7037;
wire n_13104;
wire n_1132;
wire n_9338;
wire n_11647;
wire n_8125;
wire n_501;
wire n_1823;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_10077;
wire n_3942;
wire n_3023;
wire n_10964;
wire n_14367;
wire n_9492;
wire n_2254;
wire n_3290;
wire n_14566;
wire n_6693;
wire n_10759;
wire n_9226;
wire n_6712;
wire n_7530;
wire n_10129;
wire n_10101;
wire n_1402;
wire n_3957;
wire n_13844;
wire n_11757;
wire n_3418;
wire n_10566;
wire n_1607;
wire n_7471;
wire n_9328;
wire n_6465;
wire n_221;
wire n_8188;
wire n_10192;
wire n_5673;
wire n_14363;
wire n_861;
wire n_11846;
wire n_11519;
wire n_14571;
wire n_8615;
wire n_5814;
wire n_1666;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_8011;
wire n_12191;
wire n_10207;
wire n_2214;
wire n_11530;
wire n_6730;
wire n_13526;
wire n_13998;
wire n_6367;
wire n_2256;
wire n_8923;
wire n_11488;
wire n_281;
wire n_3326;
wire n_11389;
wire n_8624;
wire n_262;
wire n_8222;
wire n_11928;
wire n_12429;
wire n_12825;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_6515;
wire n_8206;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_9513;
wire n_11315;
wire n_3224;
wire n_9393;
wire n_13267;
wire n_1969;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_13506;
wire n_8065;
wire n_9914;
wire n_14398;
wire n_527;
wire n_2949;
wire n_7008;
wire n_12318;
wire n_12918;
wire n_14731;
wire n_7709;
wire n_6468;
wire n_4269;
wire n_1927;
wire n_7540;
wire n_10886;
wire n_12923;
wire n_13632;
wire n_14600;
wire n_10804;
wire n_7581;
wire n_12077;
wire n_343;
wire n_10362;
wire n_1222;
wire n_7139;
wire n_10437;
wire n_10384;
wire n_13834;
wire n_8935;
wire n_14213;
wire n_13444;
wire n_10885;
wire n_11962;
wire n_11002;
wire n_3803;
wire n_14331;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_13885;
wire n_12805;
wire n_1791;
wire n_7782;
wire n_7432;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_13067;
wire n_8155;
wire n_9334;
wire n_2449;
wire n_14059;
wire n_11648;
wire n_10093;
wire n_13924;
wire n_14289;
wire n_4428;
wire n_12808;
wire n_745;
wire n_6483;
wire n_1572;
wire n_7770;
wire n_12853;
wire n_9684;
wire n_12591;
wire n_8397;
wire n_8568;
wire n_4463;
wire n_10600;
wire n_10480;
wire n_11994;
wire n_5357;
wire n_8175;
wire n_7173;
wire n_3648;
wire n_10796;
wire n_9254;
wire n_6576;
wire n_6810;
wire n_10003;
wire n_1975;
wire n_5421;
wire n_9083;
wire n_11050;
wire n_11250;
wire n_1388;
wire n_1266;
wire n_11316;
wire n_14727;
wire n_14485;
wire n_12987;
wire n_4396;
wire n_13717;
wire n_1990;
wire n_6708;
wire n_12251;
wire n_10252;
wire n_12948;
wire n_8026;
wire n_6667;
wire n_9175;
wire n_9838;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_11428;
wire n_2474;
wire n_12467;
wire n_12756;
wire n_2623;
wire n_11463;
wire n_1075;
wire n_6040;
wire n_10495;
wire n_1890;
wire n_6847;
wire n_8974;
wire n_6305;
wire n_8836;
wire n_10812;
wire n_4034;
wire n_12678;
wire n_14211;
wire n_4228;
wire n_14641;
wire n_12700;
wire n_1227;
wire n_11674;
wire n_11097;
wire n_11069;
wire n_12602;
wire n_10894;
wire n_3166;
wire n_14155;
wire n_7251;
wire n_12194;
wire n_7356;
wire n_3649;
wire n_7412;
wire n_3065;
wire n_8168;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_11318;
wire n_7751;
wire n_12351;
wire n_7951;
wire n_12965;
wire n_657;
wire n_7060;
wire n_14184;
wire n_3924;
wire n_9336;
wire n_3997;
wire n_12367;
wire n_13603;
wire n_8873;
wire n_14111;
wire n_10311;
wire n_7591;
wire n_10702;
wire n_3564;
wire n_862;
wire n_7444;
wire n_2637;
wire n_6750;
wire n_10490;
wire n_5769;
wire n_7911;
wire n_3795;
wire n_7595;
wire n_4931;
wire n_2306;
wire n_7790;
wire n_11586;
wire n_2071;
wire n_7426;
wire n_11786;
wire n_430;
wire n_13571;
wire n_4400;
wire n_3953;
wire n_7502;
wire n_2414;
wire n_13492;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_10906;
wire n_1532;
wire n_6855;
wire n_10891;
wire n_10840;
wire n_8170;
wire n_14257;
wire n_1030;
wire n_5181;
wire n_6239;
wire n_10181;
wire n_3208;
wire n_13673;
wire n_12036;
wire n_9554;
wire n_14589;
wire n_5768;
wire n_1342;
wire n_11330;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_8120;
wire n_12263;
wire n_9116;
wire n_9830;
wire n_9315;
wire n_8825;
wire n_14416;
wire n_852;
wire n_9169;
wire n_2916;
wire n_7252;
wire n_11201;
wire n_1060;
wire n_5963;
wire n_9999;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_7532;
wire n_12703;
wire n_4192;
wire n_8003;
wire n_11979;
wire n_12253;
wire n_9215;
wire n_1748;
wire n_1301;
wire n_6789;
wire n_8395;
wire n_3400;
wire n_5972;
wire n_13986;
wire n_7065;
wire n_1466;
wire n_8083;
wire n_11888;
wire n_6177;
wire n_14596;
wire n_8057;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_9259;
wire n_5146;
wire n_7367;
wire n_10755;
wire n_14274;
wire n_11835;
wire n_11537;
wire n_8164;
wire n_10525;
wire n_11583;
wire n_12776;
wire n_14714;
wire n_7405;
wire n_7267;
wire n_4646;
wire n_4221;
wire n_12445;
wire n_1037;
wire n_3650;
wire n_8877;
wire n_1329;
wire n_6825;
wire n_7614;
wire n_1993;
wire n_1545;
wire n_6460;
wire n_4035;
wire n_9150;
wire n_6952;
wire n_9595;
wire n_1480;
wire n_3670;
wire n_11420;
wire n_8366;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_8476;
wire n_1605;
wire n_11527;
wire n_3060;
wire n_6218;
wire n_10435;
wire n_10342;
wire n_11048;
wire n_7685;
wire n_14584;
wire n_11933;
wire n_6486;
wire n_13826;
wire n_2984;
wire n_4009;
wire n_11900;
wire n_157;
wire n_12620;
wire n_7619;
wire n_11106;
wire n_2489;
wire n_12299;
wire n_13078;
wire n_5013;
wire n_4145;
wire n_10983;
wire n_11266;
wire n_6852;
wire n_11340;
wire n_11929;
wire n_624;
wire n_5577;
wire n_876;
wire n_12673;
wire n_13557;
wire n_9100;
wire n_7883;
wire n_13516;
wire n_5872;
wire n_10397;
wire n_6692;
wire n_13208;
wire n_9707;
wire n_5017;
wire n_8854;
wire n_736;
wire n_13523;
wire n_12834;
wire n_10202;
wire n_14549;
wire n_12821;
wire n_10677;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_7560;
wire n_1327;
wire n_10648;
wire n_1475;
wire n_2106;
wire n_9262;
wire n_5976;
wire n_4717;
wire n_9249;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_602;
wire n_11964;
wire n_12247;
wire n_13030;
wire n_854;
wire n_8256;
wire n_2091;
wire n_393;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_13065;
wire n_7270;
wire n_14751;
wire n_10273;
wire n_12927;
wire n_1658;
wire n_12324;
wire n_12817;
wire n_1072;
wire n_11255;
wire n_8621;
wire n_13753;
wire n_1305;
wire n_11751;
wire n_4750;
wire n_2348;
wire n_10978;
wire n_9806;
wire n_10834;
wire n_1873;
wire n_13430;
wire n_8577;
wire n_9019;
wire n_10097;
wire n_13880;
wire n_2667;
wire n_2725;
wire n_9361;
wire n_3746;
wire n_7731;
wire n_13050;
wire n_13175;
wire n_4537;
wire n_6626;
wire n_1046;
wire n_10890;
wire n_5838;
wire n_13732;
wire n_10816;
wire n_7034;
wire n_8654;
wire n_3694;
wire n_12887;
wire n_13133;
wire n_6854;
wire n_7940;
wire n_771;
wire n_6793;
wire n_14188;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_9814;
wire n_2307;
wire n_11930;
wire n_421;
wire n_3702;
wire n_5930;
wire n_11269;
wire n_10462;
wire n_12316;
wire n_12539;
wire n_13358;
wire n_8952;
wire n_13823;
wire n_12758;
wire n_1984;
wire n_12414;
wire n_3453;
wire n_9438;
wire n_1556;
wire n_7537;
wire n_12600;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_11985;
wire n_4427;
wire n_7458;
wire n_1824;
wire n_7740;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_819;
wire n_12949;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1324;
wire n_3543;
wire n_9856;
wire n_8421;
wire n_11205;
wire n_7179;
wire n_10832;
wire n_1776;
wire n_3448;
wire n_7433;
wire n_13499;
wire n_4279;
wire n_14057;
wire n_9327;
wire n_9313;
wire n_605;
wire n_3609;
wire n_2936;
wire n_4330;
wire n_13560;
wire n_6334;
wire n_6257;
wire n_10142;
wire n_4152;
wire n_6874;
wire n_14079;
wire n_14073;
wire n_10300;
wire n_8911;
wire n_5537;
wire n_9518;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_7658;
wire n_3017;
wire n_10335;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_10753;
wire n_14220;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_12783;
wire n_13658;
wire n_807;
wire n_5142;
wire n_12431;
wire n_10921;
wire n_10177;
wire n_8971;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_10567;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_7226;
wire n_11915;
wire n_7987;
wire n_9291;
wire n_1987;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_9009;
wire n_2368;
wire n_9882;
wire n_6377;
wire n_802;
wire n_10492;
wire n_14137;
wire n_12061;
wire n_5401;
wire n_4595;
wire n_960;
wire n_7272;
wire n_11873;
wire n_8215;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_12628;
wire n_790;
wire n_9722;
wire n_5551;
wire n_5416;
wire n_14175;
wire n_4404;
wire n_2377;
wire n_14644;
wire n_151;
wire n_7906;
wire n_2652;
wire n_11260;
wire n_5498;
wire n_5543;
wire n_12359;
wire n_4054;
wire n_9760;
wire n_6018;
wire n_7765;
wire n_14320;
wire n_1286;
wire n_6021;
wire n_11880;
wire n_11605;
wire n_13615;
wire n_4617;
wire n_14022;
wire n_12974;
wire n_13156;
wire n_1685;
wire n_10741;
wire n_2477;
wire n_4611;
wire n_10037;
wire n_8949;
wire n_2279;
wire n_3169;
wire n_12136;
wire n_2222;
wire n_5797;
wire n_9454;
wire n_10760;
wire n_6511;
wire n_13849;
wire n_12121;
wire n_7815;
wire n_1052;
wire n_12658;
wire n_11838;
wire n_13956;
wire n_4732;
wire n_14768;
wire n_10607;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_13702;
wire n_8983;
wire n_4969;
wire n_11089;
wire n_14314;
wire n_8121;
wire n_5252;
wire n_11629;
wire n_11259;
wire n_5777;
wire n_11100;
wire n_13119;
wire n_8942;
wire n_7785;
wire n_11608;
wire n_13756;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_12364;
wire n_14628;
wire n_13867;
wire n_566;
wire n_7728;
wire n_8280;
wire n_2607;
wire n_11632;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_169;
wire n_12156;
wire n_7181;
wire n_11443;
wire n_173;
wire n_2796;
wire n_858;
wire n_13409;
wire n_13832;
wire n_5393;
wire n_10658;
wire n_8328;
wire n_4817;
wire n_8861;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_8427;
wire n_11161;
wire n_2136;
wire n_11770;
wire n_433;
wire n_13509;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_14399;
wire n_2771;
wire n_6322;
wire n_7359;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_11466;
wire n_10489;
wire n_9826;
wire n_253;
wire n_928;
wire n_9937;
wire n_10347;
wire n_12632;
wire n_3769;
wire n_11810;
wire n_7825;
wire n_13168;
wire n_1565;
wire n_4437;
wire n_6419;
wire n_7916;
wire n_13581;
wire n_10952;
wire n_3055;
wire n_8194;
wire n_420;
wire n_10758;
wire n_4070;
wire n_5346;
wire n_7283;
wire n_9453;
wire n_748;
wire n_7903;
wire n_9900;
wire n_12033;
wire n_7089;
wire n_1045;
wire n_8217;
wire n_14534;
wire n_10518;
wire n_9331;
wire n_1881;
wire n_2635;
wire n_7604;
wire n_7647;
wire n_2999;
wire n_988;
wire n_11789;
wire n_12465;
wire n_13447;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_330;
wire n_14164;
wire n_14771;
wire n_5868;
wire n_6417;
wire n_328;
wire n_368;
wire n_8521;
wire n_8285;
wire n_10808;
wire n_1958;
wire n_12358;
wire n_7145;
wire n_4867;
wire n_3667;
wire n_12446;
wire n_9178;
wire n_7803;
wire n_9689;
wire n_13999;
wire n_2713;
wire n_1422;
wire n_8448;
wire n_14526;
wire n_1965;
wire n_644;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_11690;
wire n_12684;
wire n_5986;
wire n_6979;
wire n_9355;
wire n_12851;
wire n_13725;
wire n_9489;
wire n_13319;
wire n_12307;
wire n_6932;
wire n_10971;
wire n_2934;
wire n_7258;
wire n_13019;
wire n_5104;
wire n_12341;
wire n_13807;
wire n_6961;
wire n_576;
wire n_8732;
wire n_511;
wire n_13297;
wire n_7622;
wire n_14610;
wire n_11968;
wire n_9359;
wire n_429;
wire n_13395;
wire n_7839;
wire n_11854;
wire n_6792;
wire n_7720;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_8136;
wire n_10404;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_1049;
wire n_11797;
wire n_8420;
wire n_13672;
wire n_141;
wire n_4430;
wire n_8386;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_7440;
wire n_10802;
wire n_1356;
wire n_9568;
wire n_6831;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_14302;
wire n_2666;
wire n_5578;
wire n_12654;
wire n_312;
wire n_728;
wire n_4409;
wire n_4191;
wire n_12921;
wire n_11991;
wire n_2401;
wire n_7809;
wire n_3255;
wire n_10340;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_14170;
wire n_935;
wire n_7072;
wire n_10681;
wire n_14303;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_11618;
wire n_911;
wire n_623;
wire n_3509;
wire n_11502;
wire n_10452;
wire n_10221;
wire n_8746;
wire n_10051;
wire n_1403;
wire n_5395;
wire n_453;
wire n_3006;
wire n_4531;
wire n_12498;
wire n_3770;
wire n_6458;
wire n_11465;
wire n_12768;
wire n_9401;
wire n_8857;
wire n_543;
wire n_11335;
wire n_6986;
wire n_9495;
wire n_3456;
wire n_12625;
wire n_13221;
wire n_10987;
wire n_4532;
wire n_236;
wire n_601;
wire n_10551;
wire n_7564;
wire n_12063;
wire n_628;
wire n_10396;
wire n_10646;
wire n_13471;
wire n_13021;
wire n_10955;
wire n_5863;
wire n_8185;
wire n_11382;
wire n_6633;
wire n_8313;
wire n_13062;
wire n_3790;
wire n_14298;
wire n_7775;
wire n_907;
wire n_9234;
wire n_7118;
wire n_13706;
wire n_7960;
wire n_6152;
wire n_9431;
wire n_5734;
wire n_10308;
wire n_10023;
wire n_8281;
wire n_12347;
wire n_847;
wire n_747;
wire n_12543;
wire n_1135;
wire n_2566;
wire n_12958;
wire n_11254;
wire n_5095;
wire n_3101;
wire n_10538;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_12532;
wire n_7069;
wire n_11388;
wire n_5199;
wire n_13347;
wire n_6546;
wire n_14051;
wire n_4257;
wire n_4282;
wire n_11043;
wire n_7636;
wire n_4341;
wire n_10199;
wire n_1694;
wire n_6925;
wire n_10673;
wire n_7186;
wire n_593;
wire n_10467;
wire n_8766;
wire n_13976;
wire n_1695;
wire n_4027;
wire n_12334;
wire n_4650;
wire n_4309;
wire n_5480;
wire n_12876;
wire n_609;
wire n_6428;
wire n_6924;
wire n_3077;
wire n_4944;
wire n_8066;
wire n_11252;
wire n_9340;
wire n_12774;
wire n_12544;
wire n_13793;
wire n_9380;
wire n_7666;
wire n_12353;
wire n_6425;
wire n_12653;
wire n_11824;
wire n_10581;
wire n_14594;
wire n_3478;
wire n_14369;
wire n_3062;
wire n_1774;
wire n_9976;
wire n_4994;
wire n_10818;
wire n_10226;
wire n_7967;
wire n_5977;
wire n_519;
wire n_14515;
wire n_8314;
wire n_384;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_1994;
wire n_11724;
wire n_3978;
wire n_12052;
wire n_11507;
wire n_3836;
wire n_11086;
wire n_10647;
wire n_13184;
wire n_9064;
wire n_3409;
wire n_4381;
wire n_8239;
wire n_9092;
wire n_14721;
wire n_3583;
wire n_11533;
wire n_4316;
wire n_7301;
wire n_11905;
wire n_14160;
wire n_4860;
wire n_4469;
wire n_9746;
wire n_12994;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_8497;
wire n_10637;
wire n_1157;
wire n_7262;
wire n_234;
wire n_5959;
wire n_13856;
wire n_8210;
wire n_10769;
wire n_3563;
wire n_8056;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_12215;
wire n_10519;
wire n_3689;
wire n_13218;
wire n_7584;
wire n_7748;
wire n_1789;
wire n_9066;
wire n_763;
wire n_14637;
wire n_6301;
wire n_2174;
wire n_13298;
wire n_540;
wire n_5668;
wire n_12535;
wire n_3442;
wire n_3972;
wire n_14248;
wire n_2315;
wire n_4209;
wire n_12582;
wire n_1687;
wire n_4703;
wire n_6282;
wire n_4934;
wire n_7686;
wire n_11800;
wire n_9870;
wire n_14391;
wire n_9817;
wire n_2638;
wire n_12505;
wire n_13396;
wire n_2046;
wire n_13988;
wire n_14648;
wire n_7059;
wire n_6985;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_13132;
wire n_395;
wire n_6737;
wire n_1587;
wire n_10723;
wire n_12875;
wire n_213;
wire n_2340;
wire n_9857;
wire n_13794;
wire n_4804;
wire n_8404;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_9455;
wire n_10056;
wire n_6459;
wire n_1427;
wire n_7670;
wire n_13400;
wire n_2977;
wire n_3991;
wire n_13813;
wire n_14307;
wire n_4936;
wire n_8505;
wire n_10653;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_585;
wire n_9916;
wire n_1617;
wire n_10157;
wire n_2600;
wire n_8606;
wire n_13542;
wire n_7443;
wire n_10701;
wire n_10470;
wire n_10923;
wire n_12828;
wire n_3436;
wire n_5973;
wire n_7484;
wire n_1962;
wire n_12402;
wire n_14387;
wire n_3806;
wire n_9440;
wire n_4759;
wire n_10038;
wire n_9059;
wire n_11691;
wire n_9812;
wire n_14666;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_6753;
wire n_9690;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_13879;
wire n_11594;
wire n_9912;
wire n_11687;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_9002;
wire n_11513;
wire n_3402;
wire n_9620;
wire n_1621;
wire n_10619;
wire n_13522;
wire n_6448;
wire n_9229;
wire n_12524;
wire n_14535;
wire n_5186;
wire n_14196;
wire n_7930;
wire n_7487;
wire n_4585;
wire n_1785;
wire n_13403;
wire n_10454;
wire n_11655;
wire n_3406;
wire n_13241;
wire n_580;
wire n_3664;
wire n_4218;
wire n_9464;
wire n_11386;
wire n_434;
wire n_4687;
wire n_7077;
wire n_14060;
wire n_10656;
wire n_394;
wire n_10871;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_8518;
wire n_11111;
wire n_4720;
wire n_2889;
wire n_13270;
wire n_11938;
wire n_6268;
wire n_12670;
wire n_6043;
wire n_9497;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_14543;
wire n_7663;
wire n_3470;
wire n_243;
wire n_8741;
wire n_8350;
wire n_10444;
wire n_11833;
wire n_5221;
wire n_7024;
wire n_1407;
wire n_11866;
wire n_8148;
wire n_8408;
wire n_6145;
wire n_12308;
wire n_2865;
wire n_10846;
wire n_12659;
wire n_13934;
wire n_13024;
wire n_5925;
wire n_6529;
wire n_973;
wire n_5591;
wire n_4762;
wire n_13223;
wire n_3844;
wire n_3259;
wire n_8236;
wire n_14202;
wire n_11192;
wire n_11229;
wire n_7214;
wire n_11244;
wire n_8806;
wire n_14352;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_8295;
wire n_1176;
wire n_9587;
wire n_3677;
wire n_1054;
wire n_13888;
wire n_7977;
wire n_14719;
wire n_5387;
wire n_13529;
wire n_12452;
wire n_3292;
wire n_6311;
wire n_11848;
wire n_8167;
wire n_8377;
wire n_13530;
wire n_3989;
wire n_7652;
wire n_13591;
wire n_10558;
wire n_9783;
wire n_4644;
wire n_8956;
wire n_4752;
wire n_8673;
wire n_4746;
wire n_7566;
wire n_14631;
wire n_1057;
wire n_4131;
wire n_11876;
wire n_12667;
wire n_5449;
wire n_8760;
wire n_4215;
wire n_978;
wire n_12707;
wire n_2488;
wire n_1509;
wire n_828;
wire n_6134;
wire n_322;
wire n_4158;
wire n_10466;
wire n_6812;
wire n_3079;
wire n_10044;
wire n_10546;
wire n_12878;
wire n_5190;
wire n_6733;
wire n_11666;
wire n_3269;
wire n_558;
wire n_5325;
wire n_13354;
wire n_10527;
wire n_4231;
wire n_8960;
wire n_8957;
wire n_9008;
wire n_10143;
wire n_12361;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_10233;
wire n_653;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_8207;
wire n_6938;
wire n_2197;
wire n_12709;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_10461;
wire n_5344;
wire n_2550;
wire n_556;
wire n_170;
wire n_1536;
wire n_3177;
wire n_6160;
wire n_10186;
wire n_4667;
wire n_5813;
wire n_10113;
wire n_12721;
wire n_6235;
wire n_1471;
wire n_13023;
wire n_6212;
wire n_3440;
wire n_9381;
wire n_9194;
wire n_6816;
wire n_8904;
wire n_3658;
wire n_12264;
wire n_14683;
wire n_7374;
wire n_12464;
wire n_13268;
wire n_12753;
wire n_3404;
wire n_2291;
wire n_13887;
wire n_3346;
wire n_2816;
wire n_12968;
wire n_1620;
wire n_2542;
wire n_10120;
wire n_5892;
wire n_9549;
wire n_7678;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_11248;
wire n_788;
wire n_13660;
wire n_7110;
wire n_5714;
wire n_12111;
wire n_2169;
wire n_6953;
wire n_9652;
wire n_7975;
wire n_9957;
wire n_13481;
wire n_12609;
wire n_13143;
wire n_12482;
wire n_8451;
wire n_6089;
wire n_591;
wire n_10591;
wire n_11780;
wire n_12966;
wire n_5634;
wire n_5133;
wire n_14607;
wire n_7553;
wire n_8527;
wire n_5305;
wire n_5990;
wire n_2175;
wire n_1625;
wire n_7732;
wire n_5689;
wire n_7086;
wire n_7891;
wire n_13383;
wire n_13419;
wire n_9089;
wire n_4578;
wire n_318;
wire n_8840;
wire n_11424;
wire n_11467;
wire n_5644;
wire n_9137;
wire n_9390;
wire n_3644;
wire n_11995;
wire n_12178;
wire n_8038;
wire n_8190;
wire n_9439;
wire n_11701;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_6138;
wire n_528;
wire n_9080;
wire n_14773;
wire n_13351;
wire n_1922;
wire n_9296;
wire n_12997;
wire n_940;
wire n_10625;
wire n_13544;
wire n_1537;
wire n_4877;
wire n_14173;
wire n_9312;
wire n_10662;
wire n_2065;
wire n_12818;
wire n_9151;
wire n_8179;
wire n_7038;
wire n_7994;
wire n_4470;
wire n_4187;
wire n_9883;
wire n_13420;
wire n_14576;
wire n_8287;
wire n_10697;
wire n_1904;
wire n_8111;
wire n_8341;
wire n_13527;
wire n_8830;
wire n_13206;
wire n_13235;
wire n_4998;
wire n_10200;
wire n_14436;
wire n_5576;
wire n_13399;
wire n_2395;
wire n_2868;
wire n_10935;
wire n_7345;
wire n_9324;
wire n_13317;
wire n_9631;
wire n_10547;
wire n_8308;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_13622;
wire n_5918;
wire n_631;
wire n_8021;
wire n_11092;
wire n_5852;
wire n_1170;
wire n_10933;
wire n_2724;
wire n_9736;
wire n_8965;
wire n_2258;
wire n_7041;
wire n_9365;
wire n_10632;
wire n_6717;
wire n_14651;
wire n_7593;
wire n_8265;
wire n_13564;
wire n_898;
wire n_11166;
wire n_6881;
wire n_10085;
wire n_3328;
wire n_2012;
wire n_9600;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_9816;
wire n_5343;
wire n_6672;
wire n_9869;
wire n_7757;
wire n_1093;
wire n_8251;
wire n_9402;
wire n_7866;
wire n_6518;
wire n_7334;
wire n_13276;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_8773;
wire n_12195;
wire n_14383;
wire n_14400;
wire n_5947;
wire n_6242;
wire n_14143;
wire n_336;
wire n_6601;
wire n_8570;
wire n_12536;
wire n_10645;
wire n_2268;
wire n_3469;
wire n_10041;
wire n_12168;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_10096;
wire n_668;
wire n_12533;
wire n_8579;
wire n_2111;
wire n_3743;
wire n_8079;
wire n_5542;
wire n_9615;
wire n_11869;
wire n_14106;
wire n_2948;
wire n_5015;
wire n_13792;
wire n_3099;
wire n_12560;
wire n_5527;
wire n_2897;
wire n_9759;
wire n_9711;
wire n_4812;
wire n_8973;
wire n_8506;
wire n_13171;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_13764;
wire n_8291;
wire n_3155;
wire n_14725;
wire n_4300;
wire n_2024;
wire n_11264;
wire n_10336;
wire n_9820;
wire n_1770;
wire n_701;
wire n_1003;
wire n_7758;
wire n_8635;
wire n_12477;
wire n_8320;
wire n_9703;
wire n_4472;
wire n_12516;
wire n_9819;
wire n_9118;
wire n_11060;
wire n_2699;
wire n_9321;
wire n_12523;
wire n_11493;
wire n_11562;
wire n_13698;
wire n_5819;
wire n_3901;
wire n_291;
wire n_5180;
wire n_1640;
wire n_8375;
wire n_10703;
wire n_11575;
wire n_2973;
wire n_10449;
wire n_10892;
wire n_13462;
wire n_10280;
wire n_9428;
wire n_8612;
wire n_10198;
wire n_8778;
wire n_11065;
wire n_5893;
wire n_9292;
wire n_11452;
wire n_2710;
wire n_7705;
wire n_6092;
wire n_12486;
wire n_6462;
wire n_2505;
wire n_11345;
wire n_4519;
wire n_9018;
wire n_13741;
wire n_5025;
wire n_2397;
wire n_8872;
wire n_12743;
wire n_240;
wire n_369;
wire n_10371;
wire n_7333;
wire n_3878;
wire n_12246;
wire n_4197;
wire n_12297;
wire n_13440;
wire n_6669;
wire n_8006;
wire n_11495;
wire n_9565;
wire n_2721;
wire n_13325;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_8491;
wire n_8218;
wire n_1212;
wire n_13089;
wire n_13578;
wire n_7337;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_7439;
wire n_12610;
wire n_4371;
wire n_5726;
wire n_14006;
wire n_14757;
wire n_10483;
wire n_188;
wire n_12771;
wire n_1902;
wire n_7744;
wire n_2784;
wire n_10346;
wire n_7210;
wire n_3898;
wire n_5828;
wire n_11864;
wire n_694;
wire n_6228;
wire n_10805;
wire n_14107;
wire n_6702;
wire n_7358;
wire n_8240;
wire n_10059;
wire n_9961;
wire n_4749;
wire n_12763;
wire n_7707;
wire n_5924;
wire n_1845;
wire n_7733;
wire n_13496;
wire n_14074;
wire n_921;
wire n_14536;
wire n_5545;
wire n_8458;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_8853;
wire n_9603;
wire n_11293;
wire n_5083;
wire n_7684;
wire n_10700;
wire n_11984;
wire n_3253;
wire n_11961;
wire n_8306;
wire n_2088;
wire n_11981;
wire n_1275;
wire n_14599;
wire n_6997;
wire n_9692;
wire n_4238;
wire n_6371;
wire n_13222;
wire n_904;
wire n_11559;
wire n_7673;
wire n_2005;
wire n_1696;
wire n_14642;
wire n_12172;
wire n_11942;
wire n_11207;
wire n_11686;
wire n_12280;
wire n_12883;
wire n_8013;
wire n_7187;
wire n_2108;
wire n_14476;
wire n_3824;
wire n_8342;
wire n_10502;
wire n_12064;
wire n_12480;
wire n_2246;
wire n_7313;
wire n_10974;
wire n_5899;
wire n_11239;
wire n_14221;
wire n_10250;
wire n_10511;
wire n_9012;
wire n_11482;
wire n_3846;
wire n_12682;
wire n_10831;
wire n_5122;
wire n_11992;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_12621;
wire n_4479;
wire n_13754;
wire n_10613;
wire n_6641;
wire n_3845;
wire n_12283;
wire n_6463;
wire n_10172;
wire n_3203;
wire n_10351;
wire n_383;
wire n_13285;
wire n_4986;
wire n_10333;
wire n_1316;
wire n_4668;
wire n_950;
wire n_9868;
wire n_711;
wire n_6264;
wire n_5782;
wire n_8119;
wire n_9264;
wire n_630;
wire n_4168;
wire n_1369;
wire n_8582;
wire n_7036;
wire n_11479;
wire n_4298;
wire n_10594;
wire n_11814;
wire n_7370;
wire n_7931;
wire n_4743;
wire n_13181;
wire n_11622;
wire n_8445;
wire n_12225;
wire n_1781;
wire n_9720;
wire n_4250;
wire n_13004;
wire n_11067;
wire n_3143;
wire n_8044;
wire n_13413;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_8363;
wire n_8464;
wire n_8921;
wire n_12208;
wire n_14072;
wire n_13608;
wire n_12126;
wire n_13397;
wire n_235;
wire n_2188;
wire n_11083;
wire n_14282;
wire n_10010;
wire n_10588;
wire n_11907;
wire n_2430;
wire n_2504;
wire n_12396;
wire n_12984;
wire n_5637;
wire n_4211;
wire n_11952;
wire n_3094;
wire n_741;
wire n_9646;
wire n_6084;
wire n_7480;
wire n_13997;
wire n_12158;
wire n_8843;
wire n_371;
wire n_13513;
wire n_5185;
wire n_8405;
wire n_13232;
wire n_2964;
wire n_13296;
wire n_13816;
wire n_14713;
wire n_8376;
wire n_308;
wire n_13859;
wire n_5032;
wire n_11506;
wire n_6990;
wire n_865;
wire n_5034;
wire n_3312;
wire n_7071;
wire n_1041;
wire n_2451;
wire n_10797;
wire n_8694;
wire n_2913;
wire n_8848;
wire n_6288;
wire n_993;
wire n_13989;
wire n_1862;
wire n_14573;
wire n_3752;
wire n_8752;
wire n_10643;
wire n_3672;
wire n_922;
wire n_1004;
wire n_8625;
wire n_8894;
wire n_7380;
wire n_14058;
wire n_2839;
wire n_8813;
wire n_3237;
wire n_7708;
wire n_12690;
wire n_12813;
wire n_11524;
wire n_10905;
wire n_9842;
wire n_11859;
wire n_4128;
wire n_11228;
wire n_12725;
wire n_4036;
wire n_9671;
wire n_5269;
wire n_8430;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_10784;
wire n_11035;
wire n_4807;
wire n_11023;
wire n_8770;
wire n_6277;
wire n_8426;
wire n_14009;
wire n_5115;
wire n_12474;
wire n_7376;
wire n_11174;
wire n_8411;
wire n_13759;
wire n_902;
wire n_8817;
wire n_8461;
wire n_10438;
wire n_1723;
wire n_3918;
wire n_10234;
wire n_10946;
wire n_11582;
wire n_9230;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_11705;
wire n_4391;
wire n_11796;
wire n_596;
wire n_12484;
wire n_9893;
wire n_6409;
wire n_4095;
wire n_8391;
wire n_8507;
wire n_1310;
wire n_12021;
wire n_5927;
wire n_9188;
wire n_8691;
wire n_11003;
wire n_4485;
wire n_9032;
wire n_7657;
wire n_6388;
wire n_10275;
wire n_574;
wire n_3593;
wire n_6839;
wire n_14284;
wire n_5163;
wire n_9614;
wire n_8967;
wire n_12990;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_9628;
wire n_1896;
wire n_9231;
wire n_10854;
wire n_6864;
wire n_14309;
wire n_13652;
wire n_1516;
wire n_13207;
wire n_4890;
wire n_10204;
wire n_8856;
wire n_8084;
wire n_2485;
wire n_12778;
wire n_12685;
wire n_6679;
wire n_12862;
wire n_11528;
wire n_10734;
wire n_13442;
wire n_10201;
wire n_8631;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_8219;
wire n_9730;
wire n_5507;
wire n_10608;
wire n_195;
wire n_4573;
wire n_1328;
wire n_10746;
wire n_4943;
wire n_2875;
wire n_10676;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_14423;
wire n_12177;
wire n_13128;
wire n_7504;
wire n_14086;
wire n_4042;
wire n_7099;
wire n_7586;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_12672;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_8428;
wire n_7052;
wire n_9172;
wire n_12141;
wire n_14665;
wire n_1634;
wire n_14342;
wire n_1203;
wire n_9926;
wire n_1699;
wire n_14634;
wire n_6738;
wire n_12665;
wire n_13719;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_11615;
wire n_11079;
wire n_8338;
wire n_14772;
wire n_1631;
wire n_7602;
wire n_9180;
wire n_9017;
wire n_12024;
wire n_156;
wire n_12795;
wire n_9269;
wire n_6566;
wire n_9026;
wire n_13453;
wire n_1794;
wire n_9462;
wire n_10900;
wire n_5696;
wire n_7998;
wire n_13370;
wire n_8666;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_204;
wire n_11438;
wire n_11700;
wire n_7557;
wire n_3772;
wire n_12940;
wire n_7408;
wire n_12555;
wire n_14539;
wire n_2891;
wire n_496;
wire n_4335;
wire n_7026;
wire n_3128;
wire n_10052;
wire n_13656;
wire n_11668;
wire n_6146;
wire n_13667;
wire n_5677;
wire n_13641;
wire n_4277;
wire n_12487;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_7394;
wire n_11387;
wire n_9515;
wire n_10560;
wire n_9502;
wire n_13103;
wire n_263;
wire n_4516;
wire n_5235;
wire n_360;
wire n_13183;
wire n_13720;
wire n_1129;
wire n_13971;
wire n_11099;
wire n_7627;
wire n_6436;
wire n_12305;
wire n_1464;
wire n_7719;
wire n_2798;
wire n_10773;
wire n_7450;
wire n_165;
wire n_9316;
wire n_3217;
wire n_11996;
wire n_8938;
wire n_6081;
wire n_13436;
wire n_14479;
wire n_10455;
wire n_1249;
wire n_14410;
wire n_329;
wire n_7852;
wire n_5724;
wire n_3821;
wire n_340;
wire n_12526;
wire n_3201;
wire n_12622;
wire n_7462;
wire n_12456;
wire n_7780;
wire n_3503;
wire n_10391;
wire n_8523;
wire n_12857;
wire n_5979;
wire n_10476;
wire n_10559;
wire n_10630;
wire n_13797;
wire n_6027;
wire n_13321;
wire n_1870;
wire n_10911;
wire n_11547;
wire n_10121;
wire n_11064;
wire n_12439;
wire n_4467;
wire n_177;
wire n_13809;
wire n_364;
wire n_258;
wire n_7582;
wire n_10540;
wire n_5521;
wire n_431;
wire n_2654;
wire n_3935;
wire n_7421;
wire n_13575;
wire n_1861;
wire n_11104;
wire n_9873;
wire n_1228;
wire n_2319;
wire n_10473;
wire n_12287;
wire n_10828;
wire n_12182;
wire n_13390;
wire n_8924;
wire n_2965;
wire n_12366;
wire n_7555;
wire n_4955;
wire n_11112;
wire n_10114;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_447;
wire n_2689;
wire n_6110;
wire n_12552;
wire n_14123;
wire n_1762;
wire n_10269;
wire n_14258;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_8380;
wire n_13371;
wire n_12777;
wire n_9978;
wire n_5241;
wire n_12492;
wire n_10418;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_13231;
wire n_5331;
wire n_7478;
wire n_3308;
wire n_6326;
wire n_841;
wire n_3204;
wire n_10672;
wire n_7451;
wire n_9494;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_14601;
wire n_11850;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_12437;
wire n_2345;
wire n_1730;
wire n_6612;
wire n_10922;
wire n_5258;

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_23),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_24),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_19),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_10),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_105),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_32),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_34),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_44),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_96),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_109),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_128),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_12),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_90),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_98),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_2),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_57),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_11),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_93),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_68),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_49),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_70),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_13),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_9),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_87),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_99),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_58),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_47),
.Y(n_171)
);

BUFx2_ASAP7_75t_R g172 ( 
.A(n_104),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_84),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_26),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_88),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_82),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_1),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_131),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_29),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_27),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_51),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_3),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_43),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_92),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_40),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_1),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_83),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_106),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_74),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_117),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_78),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_33),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_81),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_133),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_59),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_30),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_55),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_62),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_38),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_53),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_60),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_64),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_89),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_52),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_16),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_95),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_6),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_10),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_91),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_85),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_56),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_119),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_35),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_129),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_126),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_54),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_102),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_76),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_135),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_127),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_112),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_6),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_21),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_37),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_22),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_2),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_116),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_100),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_20),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_0),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_14),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_110),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_77),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_25),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_65),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_122),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_28),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_48),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_86),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_103),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_50),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_31),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_97),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_121),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_4),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_8),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_67),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_120),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_3),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_72),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_79),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_111),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_9),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_36),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_46),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_113),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_71),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_18),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_41),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_132),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_17),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_39),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_15),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_118),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_8),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_4),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_75),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_255),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_268),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_141),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_187),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_137),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_181),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_183),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_177),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_194),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_213),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_243),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_155),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_227),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_228),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_167),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_182),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_201),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_180),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_187),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_211),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_187),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_221),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_221),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_136),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_186),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_209),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_138),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_232),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_142),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_247),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_157),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_248),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_223),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_161),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_251),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_267),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_139),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_266),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_162),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_143),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_164),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_171),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_278),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_303),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_274),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_277),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_280),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_202),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_270),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_173),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_276),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_281),
.B(n_144),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_145),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_271),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_279),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_311),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_295),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_296),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_298),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_300),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_146),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_275),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_272),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_305),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_294),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_287),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_297),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_308),
.B(n_188),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_292),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_293),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_288),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_304),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_301),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_286),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_290),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_273),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_273),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_273),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_289),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_289),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_291),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_352),
.Y(n_362)
);

BUFx8_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_329),
.Y(n_364)
);

AND2x6_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_187),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_314),
.A2(n_172),
.B1(n_160),
.B2(n_154),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_344),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_322),
.B(n_151),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_192),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_343),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_358),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_316),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_346),
.B(n_291),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_318),
.Y(n_375)
);

INVx5_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_355),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_355),
.Y(n_378)
);

OA21x2_ASAP7_75t_L g379 ( 
.A1(n_359),
.A2(n_230),
.B(n_253),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_345),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_339),
.B(n_196),
.Y(n_383)
);

OA21x2_ASAP7_75t_L g384 ( 
.A1(n_350),
.A2(n_240),
.B(n_236),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_199),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_315),
.B(n_0),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_320),
.B(n_291),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_330),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_204),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_349),
.B(n_214),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_324),
.B(n_291),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_342),
.B(n_216),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_353),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_331),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_325),
.Y(n_399)
);

AND2x2_ASAP7_75t_SL g400 ( 
.A(n_321),
.B(n_140),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_332),
.B(n_217),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_333),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_335),
.A2(n_250),
.B(n_235),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_341),
.B(n_147),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_336),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_336),
.Y(n_407)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_317),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_348),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_347),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_323),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_327),
.B(n_231),
.Y(n_412)
);

INVx5_ASAP7_75t_L g413 ( 
.A(n_315),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_313),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_352),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_346),
.A2(n_262),
.B1(n_261),
.B2(n_256),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_322),
.B(n_148),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_358),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_358),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_322),
.B(n_149),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_334),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_358),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_339),
.B(n_249),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_322),
.A2(n_254),
.B(n_258),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_334),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_346),
.A2(n_197),
.B1(n_265),
.B2(n_264),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_334),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_352),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_339),
.B(n_150),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_314),
.A2(n_224),
.B1(n_205),
.B2(n_260),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_330),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_334),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_346),
.A2(n_269),
.B1(n_263),
.B2(n_259),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_316),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_322),
.B(n_191),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_358),
.Y(n_438)
);

OA21x2_ASAP7_75t_L g439 ( 
.A1(n_359),
.A2(n_184),
.B(n_159),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_330),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_330),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_330),
.B(n_252),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_352),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_323),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_354),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_352),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_334),
.Y(n_448)
);

AOI22x1_ASAP7_75t_SL g449 ( 
.A1(n_314),
.A2(n_189),
.B1(n_241),
.B2(n_239),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_357),
.B(n_245),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_346),
.A2(n_190),
.B1(n_246),
.B2(n_244),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_359),
.A2(n_179),
.B(n_242),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_334),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_339),
.B(n_178),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_344),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_344),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_322),
.B(n_185),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_334),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_334),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_314),
.A2(n_176),
.B1(n_238),
.B2(n_237),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_324),
.B(n_175),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_334),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_316),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_352),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_334),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_322),
.A2(n_174),
.B1(n_234),
.B2(n_233),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_352),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_322),
.B(n_170),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_339),
.B(n_169),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_334),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_352),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_357),
.B(n_192),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_352),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_357),
.B(n_192),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_316),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_357),
.B(n_192),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_334),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_322),
.A2(n_168),
.B1(n_229),
.B2(n_226),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_352),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_330),
.B(n_166),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_352),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_358),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_346),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_322),
.B(n_165),
.Y(n_484)
);

OA21x2_ASAP7_75t_L g485 ( 
.A1(n_359),
.A2(n_193),
.B(n_225),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_344),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_336),
.Y(n_487)
);

BUFx8_ASAP7_75t_L g488 ( 
.A(n_314),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_373),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_484),
.B(n_163),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_472),
.B(n_5),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_446),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_375),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_380),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_483),
.B(n_5),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_381),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_397),
.B(n_207),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_368),
.B(n_158),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_362),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_388),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_445),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_417),
.B(n_222),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_361),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_377),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_404),
.B(n_156),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_377),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_411),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_371),
.Y(n_509)
);

NAND2x1p5_ASAP7_75t_L g510 ( 
.A(n_408),
.B(n_195),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_421),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_442),
.B(n_220),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_401),
.A2(n_153),
.B1(n_219),
.B2(n_218),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_426),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_429),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_371),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_448),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_453),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_418),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_413),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_458),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_433),
.Y(n_523)
);

INVx6_ASAP7_75t_L g524 ( 
.A(n_406),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_418),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_459),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_400),
.B(n_152),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_462),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_465),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_470),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_367),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_477),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_413),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_364),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_390),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_415),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_424),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_430),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_443),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_390),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_447),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_464),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_398),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_398),
.Y(n_545)
);

OA21x2_ASAP7_75t_L g546 ( 
.A1(n_425),
.A2(n_206),
.B(n_215),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_412),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_419),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_413),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_392),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_467),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_422),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_420),
.B(n_212),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_471),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_473),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_479),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_481),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_436),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_463),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_475),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_386),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_422),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_438),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_372),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_378),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_376),
.Y(n_567)
);

OA21x2_ASAP7_75t_L g568 ( 
.A1(n_403),
.A2(n_210),
.B(n_200),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_389),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_444),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_374),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_395),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_394),
.B(n_7),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_384),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_444),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_472),
.B(n_198),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_384),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_482),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_474),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_474),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_476),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_476),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_376),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_437),
.B(n_257),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_376),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_423),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_366),
.B(n_42),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_482),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_379),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_379),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_457),
.B(n_257),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_439),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_439),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_399),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_370),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_370),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_367),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_387),
.A2(n_257),
.B1(n_203),
.B2(n_195),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_408),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_468),
.B(n_257),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_402),
.B(n_203),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_452),
.Y(n_602)
);

OAI22xp33_ASAP7_75t_SL g603 ( 
.A1(n_416),
.A2(n_203),
.B1(n_195),
.B2(n_66),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_396),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_440),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_485),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_396),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_487),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_450),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_450),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_385),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_485),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_427),
.B(n_203),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_408),
.B(n_195),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_480),
.B(n_45),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_365),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_455),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_428),
.B(n_61),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_385),
.Y(n_619)
);

AND2x2_ASAP7_75t_SL g620 ( 
.A(n_441),
.B(n_455),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_383),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_393),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_393),
.Y(n_623)
);

OA21x2_ASAP7_75t_L g624 ( 
.A1(n_461),
.A2(n_69),
.B(n_94),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_365),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_456),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_365),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_369),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_369),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_456),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_369),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_431),
.B(n_125),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_454),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_469),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_391),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_405),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_435),
.B(n_115),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_451),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_432),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_407),
.Y(n_640)
);

INVx6_ASAP7_75t_L g641 ( 
.A(n_363),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_414),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_486),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_466),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_478),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_460),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_449),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_L g648 ( 
.A(n_409),
.B(n_123),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_486),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_488),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_410),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_387),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_373),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_373),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_373),
.Y(n_655)
);

CKINVDCx8_ASAP7_75t_R g656 ( 
.A(n_406),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_411),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_373),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_411),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_373),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_373),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_377),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_411),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_446),
.Y(n_664)
);

CKINVDCx6p67_ASAP7_75t_R g665 ( 
.A(n_406),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_373),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_373),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_373),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_442),
.B(n_480),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_SL g670 ( 
.A(n_428),
.B(n_441),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_445),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_377),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_412),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_483),
.B(n_330),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_442),
.B(n_480),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_373),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_373),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_484),
.B(n_483),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_445),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_373),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_373),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_377),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_373),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_373),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_377),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_373),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_362),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_411),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_483),
.B(n_330),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_362),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_362),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_373),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_362),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_445),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_371),
.Y(n_695)
);

AND2x6_ASAP7_75t_L g696 ( 
.A(n_472),
.B(n_474),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_373),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_446),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_373),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_373),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_373),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_362),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_373),
.Y(n_703)
);

XOR2xp5_ASAP7_75t_L g704 ( 
.A(n_445),
.B(n_314),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_484),
.B(n_483),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_373),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_362),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_373),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_373),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_373),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_446),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_446),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_446),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_373),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_362),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_362),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_362),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_377),
.Y(n_718)
);

CKINVDCx16_ASAP7_75t_R g719 ( 
.A(n_406),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_373),
.Y(n_720)
);

NOR2x1_ASAP7_75t_L g721 ( 
.A(n_428),
.B(n_441),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_446),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_373),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_446),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_362),
.Y(n_725)
);

OA21x2_ASAP7_75t_L g726 ( 
.A1(n_425),
.A2(n_403),
.B(n_378),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_373),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_SL g728 ( 
.A1(n_387),
.A2(n_303),
.B1(n_445),
.B2(n_314),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_484),
.B(n_483),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_362),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_472),
.B(n_474),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_362),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_373),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_483),
.B(n_330),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_377),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_362),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_362),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_445),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_362),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_377),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_373),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_442),
.B(n_480),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_373),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_377),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_483),
.B(n_401),
.C(n_331),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_SL g746 ( 
.A1(n_387),
.A2(n_303),
.B1(n_445),
.B2(n_314),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_373),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_373),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_483),
.B(n_330),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_373),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_362),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_373),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_373),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_445),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_362),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_373),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_362),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_484),
.B(n_483),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_362),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_377),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_373),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_483),
.A2(n_401),
.B1(n_484),
.B2(n_480),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_362),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_362),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_373),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_373),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_362),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_373),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_373),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_446),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_362),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_484),
.B(n_483),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_411),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_484),
.B(n_483),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_373),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_373),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_446),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_472),
.B(n_474),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_472),
.B(n_474),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_362),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_373),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_362),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_445),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_362),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_377),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_362),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_445),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_446),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_362),
.Y(n_789)
);

NOR2x1p5_ASAP7_75t_L g790 ( 
.A(n_665),
.B(n_523),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_762),
.B(n_678),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_489),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_524),
.Y(n_793)
);

INVx5_ASAP7_75t_L g794 ( 
.A(n_696),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_499),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_538),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_524),
.B(n_641),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_539),
.Y(n_798)
);

OR2x6_ASAP7_75t_L g799 ( 
.A(n_641),
.B(n_536),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_505),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_505),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_547),
.B(n_673),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_505),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_502),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_749),
.B(n_729),
.C(n_705),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_492),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_639),
.A2(n_646),
.B1(n_778),
.B2(n_731),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_493),
.Y(n_808)
);

BUFx4f_ASAP7_75t_L g809 ( 
.A(n_536),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_758),
.B(n_772),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_SL g811 ( 
.A1(n_527),
.A2(n_607),
.B1(n_604),
.B2(n_611),
.Y(n_811)
);

BUFx6f_ASAP7_75t_SL g812 ( 
.A(n_620),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_494),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_507),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_774),
.B(n_638),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_696),
.B(n_586),
.Y(n_816)
);

OAI22xp33_ASAP7_75t_L g817 ( 
.A1(n_745),
.A2(n_633),
.B1(n_634),
.B2(n_605),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_548),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_496),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_674),
.B(n_689),
.Y(n_820)
);

BUFx10_ASAP7_75t_L g821 ( 
.A(n_618),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_734),
.B(n_509),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_L g823 ( 
.A(n_497),
.B(n_513),
.C(n_550),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_500),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_597),
.B(n_532),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_507),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_696),
.B(n_506),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_509),
.B(n_517),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_687),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_690),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_679),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_691),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_507),
.Y(n_833)
);

BUFx8_ASAP7_75t_SL g834 ( 
.A(n_679),
.Y(n_834)
);

AO22x2_ASAP7_75t_L g835 ( 
.A1(n_704),
.A2(n_587),
.B1(n_491),
.B2(n_731),
.Y(n_835)
);

OR2x6_ASAP7_75t_L g836 ( 
.A(n_541),
.B(n_544),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_669),
.A2(n_675),
.B1(n_742),
.B2(n_491),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_573),
.B(n_571),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_501),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_693),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_653),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_654),
.B(n_655),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_495),
.A2(n_778),
.B1(n_779),
.B2(n_645),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_509),
.B(n_517),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_658),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_660),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_661),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_694),
.Y(n_848)
);

NOR2x1p5_ASAP7_75t_L g849 ( 
.A(n_650),
.B(n_608),
.Y(n_849)
);

NAND3xp33_ASAP7_75t_L g850 ( 
.A(n_644),
.B(n_642),
.C(n_490),
.Y(n_850)
);

AND2x6_ASAP7_75t_L g851 ( 
.A(n_779),
.B(n_618),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_694),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_598),
.A2(n_576),
.B1(n_619),
.B2(n_580),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_671),
.B(n_754),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_597),
.B(n_649),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_702),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_666),
.Y(n_857)
);

INVxp33_ASAP7_75t_L g858 ( 
.A(n_704),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_579),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_667),
.Y(n_860)
);

AND3x1_ASAP7_75t_L g861 ( 
.A(n_647),
.B(n_659),
.C(n_657),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_548),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_649),
.B(n_576),
.Y(n_863)
);

INVxp33_ASAP7_75t_SL g864 ( 
.A(n_663),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_738),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_517),
.B(n_588),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_581),
.A2(n_582),
.B1(n_596),
.B2(n_595),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_662),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_492),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_707),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_668),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_588),
.B(n_562),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_609),
.A2(n_610),
.B1(n_623),
.B2(n_622),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_715),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_662),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_716),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_537),
.A2(n_557),
.B1(n_556),
.B2(n_555),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_676),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_662),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_717),
.Y(n_880)
);

AND2x6_ASAP7_75t_L g881 ( 
.A(n_616),
.B(n_588),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_632),
.A2(n_601),
.B1(n_695),
.B2(n_525),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_677),
.Y(n_883)
);

INVxp67_ASAP7_75t_SL g884 ( 
.A(n_664),
.Y(n_884)
);

BUFx4f_ASAP7_75t_L g885 ( 
.A(n_541),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_680),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_562),
.B(n_563),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_725),
.Y(n_888)
);

INVxp33_ASAP7_75t_L g889 ( 
.A(n_728),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_672),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_730),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_563),
.B(n_599),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_672),
.Y(n_893)
);

AND3x2_ASAP7_75t_L g894 ( 
.A(n_738),
.B(n_787),
.C(n_783),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_681),
.B(n_683),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_684),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_783),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_672),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_686),
.B(n_692),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_697),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_711),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_787),
.B(n_652),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_699),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_700),
.B(n_701),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_732),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_703),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_736),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_599),
.B(n_525),
.Y(n_908)
);

OR2x6_ASAP7_75t_L g909 ( 
.A(n_544),
.B(n_545),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_711),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_621),
.B(n_508),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_575),
.B(n_695),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_706),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_682),
.Y(n_914)
);

OR2x6_ASAP7_75t_L g915 ( 
.A(n_545),
.B(n_713),
.Y(n_915)
);

INVx5_ASAP7_75t_L g916 ( 
.A(n_575),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_614),
.B(n_670),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_708),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_709),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_614),
.B(n_498),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_737),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_739),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_710),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_714),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_617),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_720),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_682),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_719),
.B(n_508),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_751),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_723),
.Y(n_930)
);

NAND2xp33_ASAP7_75t_L g931 ( 
.A(n_721),
.B(n_503),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_755),
.Y(n_932)
);

OAI22xp33_ASAP7_75t_L g933 ( 
.A1(n_636),
.A2(n_640),
.B1(n_656),
.B2(n_776),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_630),
.B(n_643),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_757),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_727),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_688),
.B(n_773),
.Y(n_937)
);

INVx5_ASAP7_75t_L g938 ( 
.A(n_713),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_626),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_626),
.B(n_520),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_540),
.A2(n_542),
.B1(n_543),
.B2(n_551),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_759),
.Y(n_942)
);

AO22x2_ASAP7_75t_L g943 ( 
.A1(n_587),
.A2(n_746),
.B1(n_635),
.B2(n_651),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_733),
.B(n_741),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_743),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_747),
.B(n_748),
.Y(n_946)
);

INVxp67_ASAP7_75t_SL g947 ( 
.A(n_698),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_682),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_770),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_750),
.B(n_752),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_712),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_685),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_685),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_763),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_722),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_764),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_770),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_753),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_685),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_724),
.B(n_777),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_767),
.Y(n_961)
);

OAI22xp33_ASAP7_75t_L g962 ( 
.A1(n_756),
.A2(n_775),
.B1(n_765),
.B2(n_769),
.Y(n_962)
);

BUFx10_ASAP7_75t_L g963 ( 
.A(n_777),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_761),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_766),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_718),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_771),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_718),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_788),
.B(n_531),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_768),
.B(n_781),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_504),
.B(n_511),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_788),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_780),
.Y(n_973)
);

OR2x6_ASAP7_75t_L g974 ( 
.A(n_552),
.B(n_566),
.Y(n_974)
);

CKINVDCx16_ASAP7_75t_R g975 ( 
.A(n_521),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_782),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_570),
.B(n_578),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_558),
.B(n_559),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_718),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_534),
.Y(n_980)
);

NOR3xp33_ASAP7_75t_L g981 ( 
.A(n_560),
.B(n_512),
.C(n_553),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_514),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_515),
.B(n_528),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_516),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_784),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_SL g986 ( 
.A(n_549),
.B(n_603),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_510),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_518),
.B(n_519),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_522),
.B(n_526),
.Y(n_989)
);

BUFx10_ASAP7_75t_L g990 ( 
.A(n_594),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_529),
.B(n_530),
.Y(n_991)
);

AND2x6_ASAP7_75t_L g992 ( 
.A(n_616),
.B(n_628),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_533),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_535),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_735),
.Y(n_995)
);

AND3x2_ASAP7_75t_L g996 ( 
.A(n_554),
.B(n_789),
.C(n_786),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_569),
.B(n_572),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_735),
.B(n_785),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_565),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_561),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_564),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_583),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_613),
.B(n_785),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_735),
.B(n_785),
.Y(n_1004)
);

OAI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_637),
.A2(n_615),
.B1(n_760),
.B2(n_744),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_740),
.Y(n_1006)
);

AND2x2_ASAP7_75t_SL g1007 ( 
.A(n_648),
.B(n_616),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_740),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_585),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_740),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_567),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_744),
.B(n_760),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_744),
.Y(n_1013)
);

OR2x6_ASAP7_75t_L g1014 ( 
.A(n_760),
.B(n_625),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_624),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_726),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_726),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_574),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_593),
.Y(n_1019)
);

NAND2xp33_ASAP7_75t_L g1020 ( 
.A(n_584),
.B(n_600),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_591),
.B(n_631),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_577),
.B(n_589),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_592),
.Y(n_1023)
);

NAND3xp33_ASAP7_75t_L g1024 ( 
.A(n_602),
.B(n_606),
.C(n_612),
.Y(n_1024)
);

NAND2xp33_ASAP7_75t_L g1025 ( 
.A(n_627),
.B(n_629),
.Y(n_1025)
);

NAND3xp33_ASAP7_75t_L g1026 ( 
.A(n_568),
.B(n_546),
.C(n_624),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_590),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_568),
.B(n_546),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_489),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_499),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_499),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_505),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_762),
.B(n_390),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_678),
.B(n_705),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_547),
.B(n_673),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_SL g1036 ( 
.A(n_523),
.B(n_433),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_548),
.Y(n_1037)
);

INVxp33_ASAP7_75t_L g1038 ( 
.A(n_704),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_499),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_489),
.Y(n_1040)
);

NAND2xp33_ASAP7_75t_L g1041 ( 
.A(n_762),
.B(n_390),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_678),
.B(n_705),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_502),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_499),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_547),
.B(n_673),
.Y(n_1045)
);

NAND3xp33_ASAP7_75t_L g1046 ( 
.A(n_547),
.B(n_673),
.C(n_749),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_547),
.B(n_673),
.Y(n_1047)
);

BUFx10_ASAP7_75t_L g1048 ( 
.A(n_523),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_499),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_548),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_678),
.B(n_705),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_499),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_R g1053 ( 
.A(n_523),
.B(n_433),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_704),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_489),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_678),
.B(n_705),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_489),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_762),
.A2(n_547),
.B1(n_673),
.B2(n_678),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_499),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_499),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_547),
.B(n_673),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_523),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_489),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_762),
.B(n_390),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_505),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_489),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_505),
.Y(n_1067)
);

OAI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_762),
.A2(n_547),
.B1(n_673),
.B2(n_678),
.Y(n_1068)
);

AND3x4_ASAP7_75t_L g1069 ( 
.A(n_721),
.B(n_647),
.C(n_396),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_762),
.B(n_390),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_678),
.B(n_705),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_548),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_762),
.A2(n_547),
.B1(n_673),
.B2(n_678),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_762),
.B(n_390),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_762),
.B(n_390),
.Y(n_1075)
);

AND3x2_ASAP7_75t_L g1076 ( 
.A(n_679),
.B(n_455),
.C(n_367),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_524),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_489),
.Y(n_1078)
);

INVx4_ASAP7_75t_L g1079 ( 
.A(n_548),
.Y(n_1079)
);

NAND2xp33_ASAP7_75t_L g1080 ( 
.A(n_762),
.B(n_390),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_499),
.Y(n_1081)
);

OR2x6_ASAP7_75t_L g1082 ( 
.A(n_524),
.B(n_641),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_704),
.B(n_671),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_678),
.B(n_705),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_505),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_505),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_547),
.B(n_673),
.Y(n_1087)
);

BUFx4f_ASAP7_75t_L g1088 ( 
.A(n_665),
.Y(n_1088)
);

OR2x2_ASAP7_75t_L g1089 ( 
.A(n_704),
.B(n_671),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_499),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_547),
.B(n_673),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_762),
.B(n_390),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_499),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_505),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_499),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_762),
.B(n_390),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_547),
.B(n_673),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_505),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_505),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_489),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_762),
.A2(n_547),
.B1(n_673),
.B2(n_678),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_548),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_489),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_502),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_548),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_489),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_489),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_489),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_489),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_489),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_499),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_499),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_762),
.B(n_390),
.Y(n_1113)
);

NAND2xp33_ASAP7_75t_L g1114 ( 
.A(n_762),
.B(n_390),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_524),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_505),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_678),
.B(n_705),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_678),
.B(n_705),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_547),
.B(n_673),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_499),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_SL g1121 ( 
.A(n_523),
.B(n_433),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_505),
.Y(n_1122)
);

INVx4_ASAP7_75t_L g1123 ( 
.A(n_548),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_499),
.Y(n_1124)
);

BUFx8_ASAP7_75t_SL g1125 ( 
.A(n_502),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_678),
.B(n_705),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_489),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_502),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_489),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_499),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_505),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_489),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_499),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_678),
.B(n_705),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_505),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_489),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_524),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_489),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_547),
.B(n_673),
.C(n_749),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_L g1140 ( 
.A(n_547),
.B(n_673),
.C(n_749),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_548),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_548),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_547),
.B(n_673),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_489),
.Y(n_1144)
);

BUFx10_ASAP7_75t_L g1145 ( 
.A(n_523),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_505),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_547),
.B(n_673),
.Y(n_1147)
);

OAI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_762),
.A2(n_547),
.B1(n_673),
.B2(n_678),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_502),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_547),
.B(n_673),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_499),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_SL g1152 ( 
.A(n_620),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_704),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_547),
.B(n_673),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_762),
.B(n_390),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_762),
.A2(n_547),
.B1(n_673),
.B2(n_678),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_731),
.B(n_778),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_499),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_499),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_523),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_505),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_489),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_762),
.B(n_390),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_704),
.B(n_671),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_489),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_505),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_499),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_547),
.B(n_673),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_696),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_639),
.A2(n_400),
.B1(n_646),
.B2(n_731),
.Y(n_1170)
);

INVx4_ASAP7_75t_L g1171 ( 
.A(n_548),
.Y(n_1171)
);

AND2x6_ASAP7_75t_L g1172 ( 
.A(n_491),
.B(n_731),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_502),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_489),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_704),
.B(n_671),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_505),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_762),
.B(n_390),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_505),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_524),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_762),
.A2(n_547),
.B1(n_673),
.B2(n_678),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_524),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_489),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_489),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_489),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_678),
.B(n_705),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_502),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_505),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_547),
.B(n_673),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_678),
.B(n_705),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_499),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_489),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_489),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_489),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_505),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_505),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_489),
.Y(n_1196)
);

NAND2xp33_ASAP7_75t_SL g1197 ( 
.A(n_599),
.B(n_428),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_505),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_762),
.B(n_390),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_678),
.B(n_705),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_489),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_704),
.B(n_671),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_489),
.Y(n_1203)
);

INVx4_ASAP7_75t_L g1204 ( 
.A(n_548),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_499),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_499),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_489),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_489),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_678),
.B(n_705),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_547),
.B(n_673),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_489),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_489),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_499),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_524),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_489),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_489),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_489),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_499),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1001),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1068),
.B(n_1148),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_991),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_813),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_991),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_813),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1051),
.B(n_1056),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_819),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_794),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_795),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1071),
.B(n_1084),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1117),
.B(n_1118),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_796),
.Y(n_1232)
);

NOR2xp67_ASAP7_75t_L g1233 ( 
.A(n_916),
.B(n_1062),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1126),
.B(n_1134),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1125),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1185),
.B(n_1189),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1200),
.A2(n_1209),
.B1(n_1058),
.B2(n_1101),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_815),
.B(n_791),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_794),
.B(n_1169),
.Y(n_1239)
);

INVxp33_ASAP7_75t_L g1240 ( 
.A(n_825),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1046),
.B(n_1139),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_810),
.B(n_1073),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1140),
.B(n_1156),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_805),
.B(n_802),
.Y(n_1244)
);

NAND3xp33_ASAP7_75t_L g1245 ( 
.A(n_1035),
.B(n_1061),
.C(n_1047),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_934),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_798),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1180),
.B(n_1036),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1121),
.B(n_1091),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_819),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_1160),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1045),
.B(n_1087),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1132),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1119),
.B(n_1147),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1132),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1154),
.B(n_1168),
.Y(n_1256)
);

OAI21xp33_ASAP7_75t_L g1257 ( 
.A1(n_1097),
.A2(n_1150),
.B(n_1143),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1188),
.B(n_1210),
.Y(n_1258)
);

NAND2xp33_ASAP7_75t_L g1259 ( 
.A(n_851),
.B(n_981),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_823),
.A2(n_850),
.B(n_827),
.C(n_838),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1170),
.B(n_855),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_925),
.Y(n_1262)
);

NAND2xp33_ASAP7_75t_L g1263 ( 
.A(n_851),
.B(n_1197),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1136),
.B(n_1138),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_809),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_820),
.B(n_864),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1136),
.B(n_1138),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1144),
.B(n_1162),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_SL g1269 ( 
.A(n_797),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_809),
.Y(n_1270)
);

NOR2xp67_ASAP7_75t_SL g1271 ( 
.A(n_928),
.B(n_916),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1144),
.B(n_1162),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_L g1273 ( 
.A(n_1041),
.B(n_1114),
.C(n_1080),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1165),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1165),
.Y(n_1275)
);

NOR3xp33_ASAP7_75t_L g1276 ( 
.A(n_817),
.B(n_1064),
.C(n_1033),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_885),
.B(n_916),
.Y(n_1277)
);

NOR2xp67_ASAP7_75t_L g1278 ( 
.A(n_938),
.B(n_793),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_829),
.Y(n_1279)
);

NAND3xp33_ASAP7_75t_L g1280 ( 
.A(n_986),
.B(n_1053),
.C(n_937),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1174),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1174),
.B(n_997),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_851),
.B(n_1172),
.Y(n_1283)
);

AND2x2_ASAP7_75t_SL g1284 ( 
.A(n_853),
.B(n_1088),
.Y(n_1284)
);

OR2x6_ASAP7_75t_L g1285 ( 
.A(n_797),
.B(n_1082),
.Y(n_1285)
);

INVx8_ASAP7_75t_L g1286 ( 
.A(n_1082),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_885),
.B(n_912),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_792),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_938),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_808),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_830),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_851),
.A2(n_854),
.B1(n_1172),
.B2(n_1069),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1172),
.B(n_842),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1172),
.B(n_895),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_899),
.B(n_904),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1070),
.B(n_1074),
.Y(n_1296)
);

NOR2x1p5_ASAP7_75t_L g1297 ( 
.A(n_1104),
.B(n_1128),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_R g1298 ( 
.A(n_1088),
.B(n_1048),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_SL g1299 ( 
.A(n_812),
.B(n_1152),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_834),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_944),
.B(n_946),
.Y(n_1301)
);

INVxp33_ASAP7_75t_L g1302 ( 
.A(n_1083),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_SL g1303 ( 
.A(n_1048),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_832),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1075),
.B(n_1092),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_912),
.B(n_951),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_807),
.B(n_837),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_SL g1308 ( 
.A(n_1145),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_840),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_950),
.A2(n_971),
.B1(n_983),
.B2(n_970),
.Y(n_1310)
);

AO221x1_ASAP7_75t_L g1311 ( 
.A1(n_835),
.A2(n_943),
.B1(n_933),
.B2(n_1005),
.C(n_962),
.Y(n_1311)
);

INVxp33_ASAP7_75t_L g1312 ( 
.A(n_1089),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_856),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_799),
.B(n_915),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_870),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1096),
.B(n_1113),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_821),
.B(n_938),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_821),
.B(n_794),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_824),
.Y(n_1319)
);

NAND3xp33_ASAP7_75t_L g1320 ( 
.A(n_882),
.B(n_1163),
.C(n_1155),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_988),
.B(n_989),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_865),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_839),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_841),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_845),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_874),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_846),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1157),
.B(n_847),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_963),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_SL g1330 ( 
.A(n_1145),
.Y(n_1330)
);

NAND2xp33_ASAP7_75t_L g1331 ( 
.A(n_881),
.B(n_1169),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1169),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_911),
.B(n_863),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1157),
.B(n_857),
.Y(n_1334)
);

NOR2x1p5_ASAP7_75t_L g1335 ( 
.A(n_1149),
.B(n_1173),
.Y(n_1335)
);

NOR2xp67_ASAP7_75t_L g1336 ( 
.A(n_1077),
.B(n_1115),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_881),
.Y(n_1337)
);

INVxp67_ASAP7_75t_SL g1338 ( 
.A(n_1186),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_876),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_880),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_843),
.B(n_960),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1177),
.B(n_1199),
.C(n_920),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1164),
.B(n_1175),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_818),
.B(n_862),
.Y(n_1344)
);

NOR3xp33_ASAP7_75t_L g1345 ( 
.A(n_822),
.B(n_848),
.C(n_831),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_860),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_888),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_818),
.B(n_862),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_871),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_878),
.B(n_883),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_886),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_896),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_900),
.B(n_903),
.Y(n_1353)
);

OR2x2_ASAP7_75t_SL g1354 ( 
.A(n_1054),
.B(n_1153),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1037),
.B(n_1050),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_906),
.B(n_913),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_918),
.B(n_919),
.Y(n_1357)
);

INVxp33_ASAP7_75t_L g1358 ( 
.A(n_1202),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_891),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1037),
.B(n_1050),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1072),
.B(n_1079),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_L g1362 ( 
.A(n_931),
.B(n_978),
.C(n_917),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_923),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_924),
.B(n_926),
.Y(n_1364)
);

NAND2xp33_ASAP7_75t_L g1365 ( 
.A(n_881),
.B(n_801),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_858),
.B(n_1038),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_963),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_930),
.B(n_936),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_945),
.Y(n_1369)
);

NAND2xp33_ASAP7_75t_L g1370 ( 
.A(n_881),
.B(n_801),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_958),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_SL g1372 ( 
.A(n_799),
.Y(n_1372)
);

INVxp33_ASAP7_75t_L g1373 ( 
.A(n_804),
.Y(n_1373)
);

AO221x1_ASAP7_75t_L g1374 ( 
.A1(n_835),
.A2(n_943),
.B1(n_939),
.B2(n_801),
.C(n_803),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_905),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_964),
.B(n_965),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_902),
.B(n_852),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_982),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1072),
.B(n_1079),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_803),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_984),
.Y(n_1381)
);

AOI221xp5_ASAP7_75t_L g1382 ( 
.A1(n_861),
.A2(n_1193),
.B1(n_1192),
.B2(n_1191),
.C(n_1207),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_993),
.B(n_994),
.Y(n_1383)
);

NOR2xp67_ASAP7_75t_L g1384 ( 
.A(n_1137),
.B(n_1179),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_907),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1029),
.B(n_1040),
.Y(n_1386)
);

OR2x6_ASAP7_75t_L g1387 ( 
.A(n_915),
.B(n_836),
.Y(n_1387)
);

NAND2xp33_ASAP7_75t_L g1388 ( 
.A(n_803),
.B(n_879),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1055),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1057),
.B(n_1063),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1066),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1078),
.B(n_1100),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1102),
.B(n_1105),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_897),
.B(n_811),
.Y(n_1394)
);

BUFx4_ASAP7_75t_L g1395 ( 
.A(n_812),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1103),
.B(n_1106),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1107),
.B(n_1108),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_921),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1109),
.B(n_1110),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_889),
.B(n_836),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_922),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1127),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_816),
.B(n_1043),
.Y(n_1403)
);

NOR2xp67_ASAP7_75t_L g1404 ( 
.A(n_1181),
.B(n_1214),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1129),
.B(n_1182),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1102),
.B(n_1105),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_909),
.B(n_969),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_SL g1408 ( 
.A(n_806),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1152),
.B(n_1123),
.Y(n_1409)
);

INVxp67_ASAP7_75t_SL g1410 ( 
.A(n_940),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1183),
.B(n_1184),
.Y(n_1411)
);

OR2x6_ASAP7_75t_L g1412 ( 
.A(n_909),
.B(n_949),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1196),
.B(n_1201),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1203),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1208),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_949),
.B(n_884),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1211),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_929),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_932),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1123),
.B(n_1141),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1212),
.B(n_1215),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1141),
.B(n_1142),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1142),
.B(n_1171),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_879),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_SL g1425 ( 
.A(n_869),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1216),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_955),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1217),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1000),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_859),
.B(n_947),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_901),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_867),
.B(n_873),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_935),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1003),
.A2(n_1007),
.B(n_1002),
.C(n_1009),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_974),
.B(n_910),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_942),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_SL g1437 ( 
.A(n_1171),
.B(n_1204),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1204),
.B(n_975),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1011),
.B(n_877),
.C(n_941),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_954),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_996),
.B(n_956),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_957),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_879),
.B(n_898),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_961),
.B(n_967),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_898),
.B(n_914),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_973),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_972),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_976),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_980),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_985),
.B(n_1030),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1031),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1039),
.B(n_1044),
.Y(n_1452)
);

NAND2xp33_ASAP7_75t_SL g1453 ( 
.A(n_790),
.B(n_908),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1049),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1052),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1059),
.B(n_1060),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1081),
.B(n_1090),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_974),
.Y(n_1458)
);

NOR2xp67_ASAP7_75t_SL g1459 ( 
.A(n_898),
.B(n_914),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_849),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_887),
.B(n_1093),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_872),
.B(n_1012),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_914),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1095),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1111),
.B(n_1112),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1120),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1124),
.B(n_1130),
.Y(n_1467)
);

NAND2xp33_ASAP7_75t_L g1468 ( 
.A(n_952),
.B(n_966),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1133),
.B(n_1151),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1027),
.B(n_1018),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_952),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1158),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_894),
.Y(n_1473)
);

NOR3xp33_ASAP7_75t_L g1474 ( 
.A(n_977),
.B(n_866),
.C(n_844),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_952),
.B(n_966),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1159),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_966),
.B(n_995),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1023),
.B(n_1019),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_995),
.B(n_1032),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1167),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_828),
.B(n_1076),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_995),
.B(n_1122),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1022),
.B(n_999),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1190),
.B(n_1218),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1205),
.B(n_1213),
.Y(n_1485)
);

AOI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_892),
.A2(n_1013),
.B1(n_1206),
.B2(n_826),
.C(n_833),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_800),
.B(n_814),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1032),
.Y(n_1488)
);

NOR2xp67_ASAP7_75t_L g1489 ( 
.A(n_800),
.B(n_814),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1006),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_998),
.B(n_1004),
.C(n_1195),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1008),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1010),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1032),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_826),
.B(n_833),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_868),
.A2(n_875),
.B1(n_890),
.B2(n_893),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_868),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_875),
.B(n_890),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_893),
.B(n_927),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1094),
.B(n_1198),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1094),
.B(n_1198),
.Y(n_1501)
);

INVxp33_ASAP7_75t_L g1502 ( 
.A(n_1094),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_927),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_948),
.B(n_953),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_990),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_L g1506 ( 
.A(n_1098),
.B(n_1198),
.C(n_1195),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1098),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_948),
.B(n_953),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1098),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_959),
.B(n_968),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_959),
.B(n_968),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_979),
.B(n_1085),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_979),
.B(n_1085),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1116),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1065),
.B(n_1086),
.Y(n_1515)
);

INVxp33_ASAP7_75t_L g1516 ( 
.A(n_1116),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1065),
.B(n_1086),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1116),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1067),
.B(n_1176),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1067),
.Y(n_1520)
);

OR2x6_ASAP7_75t_L g1521 ( 
.A(n_1014),
.B(n_987),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1099),
.B(n_1166),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_990),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1099),
.B(n_1187),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1131),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1131),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1014),
.B(n_1187),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1122),
.B(n_1195),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1135),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1135),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1161),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1161),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1166),
.B(n_1178),
.Y(n_1533)
);

NOR3xp33_ASAP7_75t_L g1534 ( 
.A(n_1176),
.B(n_1178),
.C(n_1021),
.Y(n_1534)
);

NAND3xp33_ASAP7_75t_L g1535 ( 
.A(n_1122),
.B(n_1194),
.C(n_1146),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1146),
.B(n_1194),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1146),
.B(n_1194),
.Y(n_1537)
);

NAND2xp33_ASAP7_75t_L g1538 ( 
.A(n_992),
.B(n_1016),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1017),
.B(n_1015),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_992),
.B(n_1024),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_992),
.B(n_1025),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_992),
.B(n_1015),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1026),
.B(n_1028),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_SL g1544 ( 
.A(n_1020),
.Y(n_1544)
);

NOR3xp33_ASAP7_75t_L g1545 ( 
.A(n_805),
.B(n_749),
.C(n_745),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_813),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_809),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1001),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1001),
.Y(n_1550)
);

AO221x1_ASAP7_75t_L g1551 ( 
.A1(n_1068),
.A2(n_673),
.B1(n_547),
.B2(n_1148),
.C(n_835),
.Y(n_1551)
);

NOR3xp33_ASAP7_75t_L g1552 ( 
.A(n_805),
.B(n_749),
.C(n_745),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_794),
.B(n_1169),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1001),
.Y(n_1554)
);

AND2x6_ASAP7_75t_L g1555 ( 
.A(n_1157),
.B(n_491),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1045),
.B(n_547),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1125),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1001),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_794),
.B(n_1169),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_813),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1068),
.B(n_390),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_794),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1001),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1034),
.B(n_547),
.Y(n_1564)
);

NOR2xp67_ASAP7_75t_L g1565 ( 
.A(n_916),
.B(n_428),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_813),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1068),
.B(n_390),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1045),
.B(n_547),
.Y(n_1569)
);

INVxp33_ASAP7_75t_L g1570 ( 
.A(n_825),
.Y(n_1570)
);

NOR2xp67_ASAP7_75t_L g1571 ( 
.A(n_916),
.B(n_428),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1068),
.B(n_390),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1034),
.B(n_547),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_794),
.B(n_1169),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_813),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1001),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1001),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1034),
.B(n_547),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_813),
.Y(n_1583)
);

NAND2xp33_ASAP7_75t_L g1584 ( 
.A(n_1034),
.B(n_390),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_825),
.Y(n_1586)
);

NAND2xp33_ASAP7_75t_L g1587 ( 
.A(n_1034),
.B(n_390),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1001),
.Y(n_1588)
);

NOR3xp33_ASAP7_75t_L g1589 ( 
.A(n_805),
.B(n_749),
.C(n_745),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_813),
.Y(n_1591)
);

OR2x6_ASAP7_75t_L g1592 ( 
.A(n_797),
.B(n_1082),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_813),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_813),
.Y(n_1594)
);

NAND2xp33_ASAP7_75t_L g1595 ( 
.A(n_1034),
.B(n_390),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1001),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1034),
.B(n_547),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_813),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_813),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_R g1603 ( 
.A(n_1053),
.B(n_523),
.Y(n_1603)
);

NOR2xp67_ASAP7_75t_L g1604 ( 
.A(n_916),
.B(n_428),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_R g1605 ( 
.A(n_1053),
.B(n_523),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_794),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_813),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_813),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_813),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1001),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1034),
.B(n_547),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_825),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_889),
.A2(n_1170),
.B1(n_639),
.B2(n_400),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_794),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_813),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1617)
);

NOR3xp33_ASAP7_75t_L g1618 ( 
.A(n_805),
.B(n_749),
.C(n_745),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_813),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1068),
.B(n_390),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_794),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1034),
.B(n_547),
.Y(n_1623)
);

NAND3xp33_ASAP7_75t_L g1624 ( 
.A(n_805),
.B(n_673),
.C(n_547),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1034),
.B(n_547),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1001),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_813),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1034),
.B(n_547),
.Y(n_1631)
);

NOR2xp67_ASAP7_75t_L g1632 ( 
.A(n_916),
.B(n_428),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_889),
.A2(n_1170),
.B1(n_639),
.B2(n_400),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1125),
.Y(n_1635)
);

AND2x2_ASAP7_75t_SL g1636 ( 
.A(n_1170),
.B(n_491),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1068),
.B(n_390),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1034),
.B(n_547),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_813),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1045),
.B(n_547),
.Y(n_1640)
);

INVx2_ASAP7_75t_SL g1641 ( 
.A(n_809),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_825),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1034),
.B(n_671),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_809),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1650)
);

INVxp33_ASAP7_75t_L g1651 ( 
.A(n_825),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1068),
.B(n_390),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1001),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_825),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_813),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_813),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1068),
.B(n_390),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1034),
.B(n_547),
.Y(n_1660)
);

AO21x2_ASAP7_75t_L g1661 ( 
.A1(n_1028),
.A2(n_1026),
.B(n_1024),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1001),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1663)
);

INVxp67_ASAP7_75t_L g1664 ( 
.A(n_825),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_813),
.Y(n_1665)
);

INVxp67_ASAP7_75t_SL g1666 ( 
.A(n_825),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1045),
.B(n_547),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_794),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_813),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1068),
.B(n_390),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1068),
.B(n_390),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1068),
.B(n_390),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1001),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_813),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_813),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1034),
.B(n_547),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1001),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_813),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_SL g1679 ( 
.A(n_797),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_SL g1680 ( 
.A(n_797),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1034),
.B(n_547),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_813),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_805),
.B(n_673),
.C(n_547),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1068),
.B(n_390),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_813),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_SL g1689 ( 
.A(n_1068),
.B(n_390),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_813),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_813),
.Y(n_1691)
);

NAND3xp33_ASAP7_75t_L g1692 ( 
.A(n_805),
.B(n_673),
.C(n_547),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1001),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1001),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1045),
.B(n_547),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_813),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1001),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_825),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_813),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_809),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1034),
.B(n_547),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1034),
.B(n_547),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1034),
.B(n_547),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1706)
);

BUFx6f_ASAP7_75t_L g1707 ( 
.A(n_794),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1068),
.B(n_390),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_825),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1068),
.B(n_390),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_813),
.Y(n_1711)
);

XOR2x2_ASAP7_75t_L g1712 ( 
.A(n_1054),
.B(n_728),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1001),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1001),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1001),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_809),
.Y(n_1716)
);

INVx4_ASAP7_75t_L g1717 ( 
.A(n_794),
.Y(n_1717)
);

OR2x6_ASAP7_75t_L g1718 ( 
.A(n_797),
.B(n_1082),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1068),
.B(n_390),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_825),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1053),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1068),
.B(n_390),
.Y(n_1724)
);

AO221x1_ASAP7_75t_L g1725 ( 
.A1(n_1068),
.A2(n_673),
.B1(n_547),
.B2(n_1148),
.C(n_835),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_794),
.B(n_1169),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1068),
.B(n_390),
.Y(n_1728)
);

INVxp33_ASAP7_75t_L g1729 ( 
.A(n_825),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1068),
.B(n_390),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_813),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1001),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1045),
.B(n_547),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1735)
);

INVxp33_ASAP7_75t_L g1736 ( 
.A(n_825),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1001),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1034),
.B(n_547),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_813),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1034),
.B(n_547),
.Y(n_1740)
);

NOR3xp33_ASAP7_75t_L g1741 ( 
.A(n_805),
.B(n_749),
.C(n_745),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_809),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1001),
.Y(n_1744)
);

NOR2xp67_ASAP7_75t_L g1745 ( 
.A(n_916),
.B(n_428),
.Y(n_1745)
);

INVxp67_ASAP7_75t_L g1746 ( 
.A(n_825),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_825),
.Y(n_1747)
);

INVx8_ASAP7_75t_L g1748 ( 
.A(n_797),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1068),
.B(n_390),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1068),
.B(n_390),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1001),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1753)
);

INVx2_ASAP7_75t_SL g1754 ( 
.A(n_809),
.Y(n_1754)
);

NOR2xp67_ASAP7_75t_L g1755 ( 
.A(n_916),
.B(n_428),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_825),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1001),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1034),
.B(n_547),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1125),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_813),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1764)
);

INVx1_ASAP7_75t_SL g1765 ( 
.A(n_825),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1034),
.B(n_547),
.Y(n_1766)
);

NOR3xp33_ASAP7_75t_L g1767 ( 
.A(n_805),
.B(n_749),
.C(n_745),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1034),
.B(n_547),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1001),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_809),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1068),
.B(n_390),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_813),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1001),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_813),
.Y(n_1775)
);

A2O1A1Ixp33_ASAP7_75t_L g1776 ( 
.A1(n_1034),
.A2(n_762),
.B(n_1051),
.C(n_1042),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1034),
.B(n_547),
.Y(n_1777)
);

NOR3xp33_ASAP7_75t_L g1778 ( 
.A(n_805),
.B(n_749),
.C(n_745),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1068),
.B(n_390),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_825),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1782)
);

INVxp67_ASAP7_75t_SL g1783 ( 
.A(n_825),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1001),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_825),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_813),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1034),
.B(n_547),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_813),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1034),
.B(n_547),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1001),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_813),
.Y(n_1793)
);

A2O1A1Ixp33_ASAP7_75t_L g1794 ( 
.A1(n_1034),
.A2(n_762),
.B(n_1051),
.C(n_1042),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1034),
.B(n_547),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1797)
);

INVx8_ASAP7_75t_L g1798 ( 
.A(n_797),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1034),
.B(n_547),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1045),
.B(n_547),
.Y(n_1801)
);

NAND3xp33_ASAP7_75t_L g1802 ( 
.A(n_805),
.B(n_673),
.C(n_547),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1034),
.B(n_547),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_SL g1804 ( 
.A(n_1036),
.B(n_433),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1001),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1068),
.B(n_390),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_794),
.Y(n_1808)
);

NOR3xp33_ASAP7_75t_L g1809 ( 
.A(n_805),
.B(n_749),
.C(n_745),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_813),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_L g1812 ( 
.A(n_805),
.B(n_673),
.C(n_547),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1813)
);

INVxp33_ASAP7_75t_L g1814 ( 
.A(n_825),
.Y(n_1814)
);

NOR3xp33_ASAP7_75t_L g1815 ( 
.A(n_805),
.B(n_749),
.C(n_745),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1068),
.B(n_390),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_794),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_813),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1068),
.B(n_390),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_809),
.Y(n_1822)
);

NOR3xp33_ASAP7_75t_L g1823 ( 
.A(n_805),
.B(n_749),
.C(n_745),
.Y(n_1823)
);

AOI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_802),
.A2(n_673),
.B1(n_547),
.B2(n_433),
.Y(n_1824)
);

INVxp33_ASAP7_75t_L g1825 ( 
.A(n_825),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1034),
.B(n_547),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1001),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1068),
.B(n_390),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1045),
.B(n_547),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1034),
.B(n_547),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1838)
);

AO221x1_ASAP7_75t_L g1839 ( 
.A1(n_1068),
.A2(n_673),
.B1(n_547),
.B2(n_1148),
.C(n_835),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_813),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_813),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1034),
.B(n_547),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1068),
.B(n_390),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1045),
.B(n_547),
.Y(n_1847)
);

INVxp33_ASAP7_75t_L g1848 ( 
.A(n_825),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1001),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_794),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_813),
.Y(n_1853)
);

BUFx6f_ASAP7_75t_L g1854 ( 
.A(n_794),
.Y(n_1854)
);

NAND2xp33_ASAP7_75t_L g1855 ( 
.A(n_1034),
.B(n_390),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1034),
.B(n_547),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_813),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1377),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1220),
.A2(n_1575),
.B1(n_1582),
.B2(n_1564),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1226),
.B(n_1856),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1599),
.B(n_1611),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1661),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1623),
.B(n_1625),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1843),
.B(n_1631),
.Y(n_1864)
);

INVxp67_ASAP7_75t_L g1865 ( 
.A(n_1343),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1661),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1638),
.B(n_1660),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1776),
.B(n_1794),
.Y(n_1868)
);

NOR2xp67_ASAP7_75t_L g1869 ( 
.A(n_1273),
.B(n_1362),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1478),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1676),
.B(n_1682),
.Y(n_1871)
);

INVx2_ASAP7_75t_SL g1872 ( 
.A(n_1286),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1478),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1470),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1703),
.B(n_1704),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1470),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1705),
.B(n_1738),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1224),
.B(n_1230),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1264),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1740),
.B(n_1760),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1264),
.Y(n_1881)
);

OAI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1310),
.A2(n_1237),
.B(n_1260),
.Y(n_1882)
);

AO22x1_ASAP7_75t_L g1883 ( 
.A1(n_1276),
.A2(n_1296),
.B1(n_1316),
.B2(n_1305),
.Y(n_1883)
);

INVx2_ASAP7_75t_SL g1884 ( 
.A(n_1286),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1254),
.B(n_1256),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1766),
.A2(n_1768),
.B1(n_1788),
.B2(n_1777),
.Y(n_1886)
);

INVx2_ASAP7_75t_SL g1887 ( 
.A(n_1286),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1267),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1254),
.B(n_1256),
.Y(n_1889)
);

AO22x1_ASAP7_75t_L g1890 ( 
.A1(n_1394),
.A2(n_1310),
.B1(n_1555),
.B2(n_1307),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1267),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1790),
.B(n_1795),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1666),
.B(n_1783),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1800),
.B(n_1803),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1245),
.B(n_1248),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1830),
.B(n_1836),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1224),
.B(n_1230),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1824),
.B(n_1244),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1311),
.A2(n_1614),
.B1(n_1634),
.B2(n_1636),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1613),
.B(n_1617),
.Y(n_1900)
);

INVx2_ASAP7_75t_SL g1901 ( 
.A(n_1748),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1246),
.B(n_1243),
.Y(n_1902)
);

NOR2xp67_ASAP7_75t_L g1903 ( 
.A(n_1717),
.B(n_1337),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1543),
.Y(n_1904)
);

CKINVDCx11_ASAP7_75t_R g1905 ( 
.A(n_1635),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1622),
.B(n_1627),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1231),
.B(n_1234),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1853),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1629),
.B(n_1630),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1231),
.A2(n_1758),
.B(n_1597),
.Y(n_1910)
);

AO221x1_ASAP7_75t_L g1911 ( 
.A1(n_1551),
.A2(n_1725),
.B1(n_1839),
.B2(n_1337),
.C(n_1280),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1633),
.B(n_1646),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_L g1913 ( 
.A(n_1234),
.B(n_1236),
.Y(n_1913)
);

AND2x2_ASAP7_75t_SL g1914 ( 
.A(n_1538),
.B(n_1331),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1857),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1648),
.B(n_1656),
.Y(n_1916)
);

AND2x2_ASAP7_75t_SL g1917 ( 
.A(n_1284),
.B(n_1337),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1657),
.B(n_1663),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1603),
.Y(n_1919)
);

INVx4_ASAP7_75t_L g1920 ( 
.A(n_1555),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1804),
.B(n_1236),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1743),
.B(n_1752),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1268),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1792),
.B(n_1796),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1268),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1272),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1797),
.B(n_1799),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1549),
.B(n_1567),
.Y(n_1928)
);

BUFx3_ASAP7_75t_L g1929 ( 
.A(n_1748),
.Y(n_1929)
);

INVx2_ASAP7_75t_SL g1930 ( 
.A(n_1748),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1272),
.B(n_1721),
.Y(n_1931)
);

AOI22xp33_ASAP7_75t_L g1932 ( 
.A1(n_1374),
.A2(n_1261),
.B1(n_1712),
.B2(n_1432),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1549),
.B(n_1567),
.Y(n_1933)
);

AOI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1257),
.A2(n_1252),
.B1(n_1574),
.B2(n_1572),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1826),
.B(n_1827),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1283),
.B(n_1239),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1572),
.B(n_1574),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1828),
.B(n_1829),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1222),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1577),
.B(n_1578),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1831),
.B(n_1833),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1577),
.B(n_1578),
.Y(n_1942)
);

BUFx2_ASAP7_75t_L g1943 ( 
.A(n_1642),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1302),
.A2(n_1358),
.B1(n_1312),
.B2(n_1341),
.Y(n_1944)
);

AND2x6_ASAP7_75t_L g1945 ( 
.A(n_1283),
.B(n_1541),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1585),
.B(n_1590),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1225),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1585),
.B(n_1590),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1597),
.B(n_1598),
.Y(n_1949)
);

BUFx6f_ASAP7_75t_L g1950 ( 
.A(n_1228),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1227),
.Y(n_1951)
);

A2O1A1Ixp33_ASAP7_75t_L g1952 ( 
.A1(n_1598),
.A2(n_1643),
.B(n_1644),
.C(n_1600),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1250),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1600),
.B(n_1643),
.Y(n_1954)
);

BUFx3_ASAP7_75t_L g1955 ( 
.A(n_1798),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1644),
.B(n_1649),
.Y(n_1956)
);

CKINVDCx20_ASAP7_75t_R g1957 ( 
.A(n_1251),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1253),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1255),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1649),
.B(n_1650),
.Y(n_1960)
);

A2O1A1Ixp33_ASAP7_75t_L g1961 ( 
.A1(n_1650),
.A2(n_1684),
.B(n_1688),
.C(n_1681),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1681),
.B(n_1684),
.Y(n_1962)
);

AOI22xp33_ASAP7_75t_L g1963 ( 
.A1(n_1439),
.A2(n_1240),
.B1(n_1651),
.B2(n_1570),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1274),
.Y(n_1964)
);

AOI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1688),
.A2(n_1699),
.B1(n_1706),
.B2(n_1693),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1654),
.Y(n_1966)
);

CKINVDCx11_ASAP7_75t_R g1967 ( 
.A(n_1235),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1693),
.B(n_1699),
.Y(n_1968)
);

BUFx5_ASAP7_75t_L g1969 ( 
.A(n_1555),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1706),
.B(n_1720),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1720),
.B(n_1723),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1275),
.Y(n_1972)
);

INVx3_ASAP7_75t_L g1973 ( 
.A(n_1553),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1723),
.B(n_1726),
.Y(n_1974)
);

BUFx3_ASAP7_75t_L g1975 ( 
.A(n_1798),
.Y(n_1975)
);

BUFx8_ASAP7_75t_L g1976 ( 
.A(n_1269),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1281),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1726),
.B(n_1734),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_SL g1979 ( 
.A1(n_1555),
.A2(n_1410),
.B1(n_1299),
.B2(n_1765),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1546),
.Y(n_1980)
);

AOI22xp33_ASAP7_75t_SL g1981 ( 
.A1(n_1555),
.A2(n_1785),
.B1(n_1320),
.B2(n_1242),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1553),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1734),
.B(n_1735),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1560),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1566),
.Y(n_1985)
);

AND2x2_ASAP7_75t_SL g1986 ( 
.A(n_1365),
.B(n_1370),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1735),
.B(n_1753),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1753),
.B(n_1756),
.Y(n_1988)
);

AOI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1729),
.A2(n_1736),
.B1(n_1825),
.B2(n_1814),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1756),
.B(n_1758),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1761),
.B(n_1764),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1761),
.B(n_1764),
.Y(n_1992)
);

INVx2_ASAP7_75t_SL g1993 ( 
.A(n_1798),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1579),
.Y(n_1994)
);

NOR3xp33_ASAP7_75t_L g1995 ( 
.A(n_1561),
.B(n_1573),
.C(n_1568),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1583),
.Y(n_1996)
);

INVx2_ASAP7_75t_SL g1997 ( 
.A(n_1285),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1769),
.B(n_1779),
.Y(n_1998)
);

INVx2_ASAP7_75t_SL g1999 ( 
.A(n_1285),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1769),
.B(n_1779),
.Y(n_2000)
);

NOR2xp67_ASAP7_75t_L g2001 ( 
.A(n_1717),
.B(n_1562),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1591),
.Y(n_2002)
);

AOI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1782),
.A2(n_1806),
.B1(n_1810),
.B2(n_1787),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1593),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1782),
.B(n_1787),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1806),
.B(n_1810),
.Y(n_2006)
);

OR2x6_ASAP7_75t_SL g2007 ( 
.A(n_1722),
.B(n_1242),
.Y(n_2007)
);

AOI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_1813),
.A2(n_1818),
.B1(n_1837),
.B2(n_1817),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1594),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1813),
.B(n_1817),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1818),
.B(n_1837),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1601),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1602),
.Y(n_2013)
);

BUFx3_ASAP7_75t_L g2014 ( 
.A(n_1285),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1607),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1838),
.A2(n_1845),
.B1(n_1846),
.B2(n_1842),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1608),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1838),
.B(n_1842),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1609),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1845),
.B(n_1846),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1849),
.B(n_1851),
.Y(n_2021)
);

INVx2_ASAP7_75t_SL g2022 ( 
.A(n_1592),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1616),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1619),
.Y(n_2024)
);

O2A1O1Ixp33_ASAP7_75t_L g2025 ( 
.A1(n_1620),
.A2(n_1652),
.B(n_1659),
.C(n_1637),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1628),
.Y(n_2026)
);

OAI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1849),
.A2(n_1851),
.B1(n_1292),
.B2(n_1645),
.Y(n_2027)
);

AOI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1848),
.A2(n_1400),
.B1(n_1366),
.B2(n_1700),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1556),
.B(n_1569),
.Y(n_2029)
);

BUFx3_ASAP7_75t_L g2030 ( 
.A(n_1592),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1640),
.B(n_1667),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1696),
.B(n_1733),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1801),
.B(n_1835),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1639),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1847),
.B(n_1295),
.Y(n_2035)
);

NOR3xp33_ASAP7_75t_L g2036 ( 
.A(n_1670),
.B(n_1672),
.C(n_1671),
.Y(n_2036)
);

OAI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1238),
.A2(n_1434),
.B(n_1686),
.Y(n_2037)
);

O2A1O1Ixp33_ASAP7_75t_L g2038 ( 
.A1(n_1689),
.A2(n_1710),
.B(n_1719),
.C(n_1708),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1295),
.B(n_1301),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1655),
.Y(n_2040)
);

INVx2_ASAP7_75t_SL g2041 ( 
.A(n_1592),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1545),
.B(n_1552),
.Y(n_2042)
);

AOI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1724),
.A2(n_1730),
.B1(n_1749),
.B2(n_1728),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1301),
.B(n_1321),
.Y(n_2044)
);

OAI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1282),
.A2(n_1364),
.B1(n_1383),
.B2(n_1368),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1658),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_1219),
.A2(n_1550),
.B1(n_1554),
.B2(n_1548),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1238),
.B(n_1282),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1589),
.B(n_1618),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1586),
.B(n_1612),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1665),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_1249),
.B(n_1750),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1669),
.Y(n_2053)
);

NAND3xp33_ASAP7_75t_L g2054 ( 
.A(n_1741),
.B(n_1778),
.C(n_1767),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_1772),
.B(n_1780),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_L g2056 ( 
.A(n_1807),
.B(n_1816),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1674),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1675),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1809),
.B(n_1815),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1664),
.B(n_1709),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1746),
.B(n_1747),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1678),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1821),
.B(n_1834),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1757),
.B(n_1781),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1258),
.B(n_1221),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1223),
.B(n_1328),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1683),
.Y(n_2067)
);

O2A1O1Ixp33_ASAP7_75t_L g2068 ( 
.A1(n_1844),
.A2(n_1241),
.B(n_1823),
.C(n_1587),
.Y(n_2068)
);

AOI22xp5_ASAP7_75t_L g2069 ( 
.A1(n_1624),
.A2(n_1692),
.B1(n_1802),
.B2(n_1685),
.Y(n_2069)
);

INVx1_ASAP7_75t_SL g2070 ( 
.A(n_1407),
.Y(n_2070)
);

BUFx3_ASAP7_75t_L g2071 ( 
.A(n_1718),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1334),
.B(n_1364),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1687),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1690),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_1373),
.B(n_1812),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1293),
.B(n_1294),
.Y(n_2076)
);

INVxp67_ASAP7_75t_L g2077 ( 
.A(n_1447),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1368),
.B(n_1383),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1386),
.B(n_1390),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_SL g2080 ( 
.A(n_1293),
.B(n_1294),
.Y(n_2080)
);

CKINVDCx20_ASAP7_75t_R g2081 ( 
.A(n_1605),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_1228),
.Y(n_2082)
);

INVxp67_ASAP7_75t_L g2083 ( 
.A(n_1266),
.Y(n_2083)
);

NOR2xp33_ASAP7_75t_L g2084 ( 
.A(n_1322),
.B(n_1333),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_SL g2085 ( 
.A(n_1382),
.B(n_1430),
.Y(n_2085)
);

NOR2xp67_ASAP7_75t_L g2086 ( 
.A(n_1562),
.B(n_1606),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1691),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1697),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_1542),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_L g2090 ( 
.A(n_1262),
.B(n_1449),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1386),
.B(n_1390),
.Y(n_2091)
);

INVx3_ASAP7_75t_L g2092 ( 
.A(n_1239),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1392),
.B(n_1399),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_1403),
.B(n_1228),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_SL g2095 ( 
.A(n_1332),
.B(n_1615),
.Y(n_2095)
);

INVx2_ASAP7_75t_SL g2096 ( 
.A(n_1718),
.Y(n_2096)
);

OAI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_1392),
.A2(n_1405),
.B1(n_1399),
.B2(n_1701),
.Y(n_2097)
);

AOI22xp33_ASAP7_75t_L g2098 ( 
.A1(n_1558),
.A2(n_1580),
.B1(n_1581),
.B2(n_1563),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1405),
.B(n_1711),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_1588),
.A2(n_1610),
.B1(n_1626),
.B2(n_1596),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_1584),
.A2(n_1595),
.B1(n_1855),
.B2(n_1259),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1731),
.B(n_1739),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1332),
.B(n_1615),
.Y(n_2103)
);

OR2x2_ASAP7_75t_L g2104 ( 
.A(n_1483),
.B(n_1763),
.Y(n_2104)
);

INVx2_ASAP7_75t_SL g2105 ( 
.A(n_1718),
.Y(n_2105)
);

NOR2x1p5_ASAP7_75t_L g2106 ( 
.A(n_1557),
.B(n_1762),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1773),
.B(n_1775),
.Y(n_2107)
);

AOI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_1653),
.A2(n_1673),
.B1(n_1677),
.B2(n_1662),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1786),
.B(n_1789),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1793),
.B(n_1811),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1820),
.Y(n_2111)
);

NOR3xp33_ASAP7_75t_L g2112 ( 
.A(n_1453),
.B(n_1338),
.C(n_1342),
.Y(n_2112)
);

BUFx6f_ASAP7_75t_L g2113 ( 
.A(n_1332),
.Y(n_2113)
);

AOI22xp33_ASAP7_75t_L g2114 ( 
.A1(n_1694),
.A2(n_1698),
.B1(n_1713),
.B2(n_1695),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1840),
.B(n_1841),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_1615),
.B(n_1621),
.Y(n_2116)
);

NAND2xp33_ASAP7_75t_L g2117 ( 
.A(n_1298),
.B(n_1621),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_SL g2118 ( 
.A(n_1269),
.B(n_1679),
.Y(n_2118)
);

INVx4_ASAP7_75t_L g2119 ( 
.A(n_1559),
.Y(n_2119)
);

NOR2xp33_ASAP7_75t_L g2120 ( 
.A(n_1287),
.B(n_1427),
.Y(n_2120)
);

NOR2xp67_ASAP7_75t_L g2121 ( 
.A(n_1606),
.B(n_1808),
.Y(n_2121)
);

O2A1O1Ixp33_ASAP7_75t_L g2122 ( 
.A1(n_1263),
.A2(n_1350),
.B(n_1356),
.C(n_1353),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1357),
.B(n_1376),
.Y(n_2123)
);

AOI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_1679),
.A2(n_1680),
.B1(n_1345),
.B2(n_1297),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_1288),
.B(n_1290),
.Y(n_2125)
);

OAI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_1396),
.A2(n_1411),
.B1(n_1413),
.B2(n_1397),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1542),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_1539),
.A2(n_1541),
.B(n_1421),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1429),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1483),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_L g2131 ( 
.A(n_1416),
.B(n_1442),
.Y(n_2131)
);

NOR2xp67_ASAP7_75t_L g2132 ( 
.A(n_1808),
.B(n_1506),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_1335),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_SL g2134 ( 
.A(n_1621),
.B(n_1668),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1319),
.B(n_1323),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1540),
.Y(n_2136)
);

NOR2xp67_ASAP7_75t_L g2137 ( 
.A(n_1535),
.B(n_1559),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1324),
.B(n_1325),
.Y(n_2138)
);

INVx3_ASAP7_75t_L g2139 ( 
.A(n_1576),
.Y(n_2139)
);

AOI22xp33_ASAP7_75t_L g2140 ( 
.A1(n_1714),
.A2(n_1732),
.B1(n_1737),
.B2(n_1715),
.Y(n_2140)
);

AOI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_1680),
.A2(n_1372),
.B1(n_1437),
.B2(n_1271),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1327),
.B(n_1346),
.Y(n_2142)
);

OAI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_1314),
.A2(n_1387),
.B1(n_1412),
.B2(n_1505),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_SL g2144 ( 
.A(n_1668),
.B(n_1707),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1349),
.B(n_1351),
.Y(n_2145)
);

BUFx6f_ASAP7_75t_L g2146 ( 
.A(n_1668),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1352),
.B(n_1363),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_SL g2148 ( 
.A(n_1707),
.B(n_1819),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_1744),
.A2(n_1759),
.B1(n_1770),
.B2(n_1751),
.Y(n_2149)
);

AOI22xp33_ASAP7_75t_L g2150 ( 
.A1(n_1774),
.A2(n_1791),
.B1(n_1805),
.B2(n_1784),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1369),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_1576),
.Y(n_2152)
);

INVx2_ASAP7_75t_SL g2153 ( 
.A(n_1727),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1832),
.Y(n_2154)
);

A2O1A1Ixp33_ASAP7_75t_L g2155 ( 
.A1(n_1462),
.A2(n_1474),
.B(n_1378),
.C(n_1381),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_SL g2156 ( 
.A(n_1707),
.B(n_1819),
.Y(n_2156)
);

O2A1O1Ixp33_ASAP7_75t_L g2157 ( 
.A1(n_1329),
.A2(n_1367),
.B(n_1277),
.C(n_1523),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_1819),
.B(n_1852),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1850),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1371),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_1442),
.B(n_1502),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_SL g2162 ( 
.A(n_1852),
.B(n_1854),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_1516),
.B(n_1438),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_1389),
.B(n_1391),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1402),
.B(n_1414),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1415),
.Y(n_2166)
);

INVx3_ASAP7_75t_L g2167 ( 
.A(n_1727),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1417),
.B(n_1426),
.Y(n_2168)
);

INVx2_ASAP7_75t_SL g2169 ( 
.A(n_1289),
.Y(n_2169)
);

OAI22xp33_ASAP7_75t_L g2170 ( 
.A1(n_1314),
.A2(n_1387),
.B1(n_1412),
.B2(n_1458),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1428),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_1527),
.B(n_1852),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1527),
.B(n_1387),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_1306),
.B(n_1460),
.Y(n_2174)
);

OAI22xp5_ASAP7_75t_SL g2175 ( 
.A1(n_1354),
.A2(n_1314),
.B1(n_1300),
.B2(n_1412),
.Y(n_2175)
);

OR2x6_ASAP7_75t_L g2176 ( 
.A(n_1854),
.B(n_1441),
.Y(n_2176)
);

AOI22xp33_ASAP7_75t_L g2177 ( 
.A1(n_1229),
.A2(n_1232),
.B1(n_1480),
.B2(n_1247),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1854),
.B(n_1380),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1435),
.B(n_1431),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_L g2180 ( 
.A(n_1380),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_1265),
.B(n_1270),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1547),
.B(n_1641),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1484),
.Y(n_2183)
);

BUFx6f_ASAP7_75t_SL g2184 ( 
.A(n_1521),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1647),
.B(n_1702),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1380),
.B(n_1463),
.Y(n_2186)
);

INVxp67_ASAP7_75t_L g2187 ( 
.A(n_1372),
.Y(n_2187)
);

OAI221xp5_ASAP7_75t_L g2188 ( 
.A1(n_1716),
.A2(n_1822),
.B1(n_1771),
.B2(n_1754),
.C(n_1742),
.Y(n_2188)
);

NOR2xp33_ASAP7_75t_L g2189 ( 
.A(n_1420),
.B(n_1423),
.Y(n_2189)
);

AOI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_1388),
.A2(n_1468),
.B(n_1487),
.Y(n_2190)
);

INVx3_ASAP7_75t_L g2191 ( 
.A(n_1463),
.Y(n_2191)
);

AOI22xp5_ASAP7_75t_L g2192 ( 
.A1(n_1481),
.A2(n_1409),
.B1(n_1425),
.B2(n_1408),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1233),
.B(n_1521),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1303),
.Y(n_2194)
);

A2O1A1Ixp33_ASAP7_75t_SL g2195 ( 
.A1(n_1499),
.A2(n_1512),
.B(n_1533),
.C(n_1522),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_SL g2196 ( 
.A(n_1463),
.B(n_1471),
.Y(n_2196)
);

INVxp67_ASAP7_75t_L g2197 ( 
.A(n_1408),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1484),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_1492),
.B(n_1493),
.Y(n_2199)
);

OAI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_1565),
.A2(n_1755),
.B1(n_1745),
.B2(n_1632),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_1471),
.B(n_1488),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1521),
.B(n_1433),
.Y(n_2202)
);

AOI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_1425),
.A2(n_1534),
.B1(n_1544),
.B2(n_1317),
.Y(n_2203)
);

INVx4_ASAP7_75t_L g2204 ( 
.A(n_1471),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1440),
.B(n_1454),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_1488),
.B(n_1494),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1464),
.B(n_1466),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_1490),
.B(n_1424),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_1488),
.B(n_1494),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1476),
.B(n_1278),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1571),
.B(n_1604),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1485),
.Y(n_2212)
);

NOR2xp33_ASAP7_75t_L g2213 ( 
.A(n_1497),
.B(n_1503),
.Y(n_2213)
);

INVxp67_ASAP7_75t_L g2214 ( 
.A(n_1461),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1485),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1444),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_1424),
.B(n_1509),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1450),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_1494),
.B(n_1507),
.Y(n_2219)
);

NOR2xp67_ASAP7_75t_L g2220 ( 
.A(n_1491),
.B(n_1509),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1452),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1279),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1291),
.B(n_1304),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_1309),
.B(n_1313),
.Y(n_2224)
);

BUFx4_ASAP7_75t_L g2225 ( 
.A(n_1395),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1315),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_SL g2227 ( 
.A(n_1507),
.B(n_1514),
.Y(n_2227)
);

OR2x6_ASAP7_75t_L g2228 ( 
.A(n_1318),
.B(n_1487),
.Y(n_2228)
);

AND2x4_ASAP7_75t_L g2229 ( 
.A(n_1489),
.B(n_1507),
.Y(n_2229)
);

AOI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_1326),
.A2(n_1436),
.B1(n_1446),
.B2(n_1419),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1456),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_1520),
.B(n_1526),
.Y(n_2232)
);

AOI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_1544),
.A2(n_1303),
.B1(n_1308),
.B2(n_1330),
.Y(n_2233)
);

OR2x6_ASAP7_75t_L g2234 ( 
.A(n_1495),
.B(n_1498),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1339),
.B(n_1340),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1457),
.Y(n_2236)
);

OR2x2_ASAP7_75t_SL g2237 ( 
.A(n_1495),
.B(n_1524),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_1308),
.Y(n_2238)
);

NOR2xp33_ASAP7_75t_L g2239 ( 
.A(n_1518),
.B(n_1525),
.Y(n_2239)
);

OAI221xp5_ASAP7_75t_L g2240 ( 
.A1(n_1336),
.A2(n_1404),
.B1(n_1384),
.B2(n_1473),
.C(n_1496),
.Y(n_2240)
);

BUFx3_ASAP7_75t_L g2241 ( 
.A(n_1514),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_SL g2242 ( 
.A(n_1330),
.B(n_1459),
.Y(n_2242)
);

A2O1A1Ixp33_ASAP7_75t_L g2243 ( 
.A1(n_1486),
.A2(n_1508),
.B(n_1513),
.C(n_1504),
.Y(n_2243)
);

AND2x6_ASAP7_75t_L g2244 ( 
.A(n_1514),
.B(n_1536),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_1347),
.B(n_1401),
.Y(n_2245)
);

BUFx6f_ASAP7_75t_SL g2246 ( 
.A(n_1529),
.Y(n_2246)
);

INVxp67_ASAP7_75t_SL g2247 ( 
.A(n_1537),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1344),
.Y(n_2248)
);

OAI21xp33_ASAP7_75t_L g2249 ( 
.A1(n_1498),
.A2(n_1519),
.B(n_1511),
.Y(n_2249)
);

NOR2x1p5_ASAP7_75t_L g2250 ( 
.A(n_1510),
.B(n_1519),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1465),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_1510),
.B(n_1511),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_1530),
.B(n_1532),
.Y(n_2253)
);

AO22x1_ASAP7_75t_L g2254 ( 
.A1(n_1531),
.A2(n_1515),
.B1(n_1524),
.B2(n_1517),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_SL g2255 ( 
.A(n_1515),
.B(n_1517),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1467),
.Y(n_2256)
);

AOI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_1348),
.A2(n_1355),
.B1(n_1422),
.B2(n_1360),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_1359),
.B(n_1451),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_1375),
.B(n_1455),
.Y(n_2259)
);

AND2x2_ASAP7_75t_SL g2260 ( 
.A(n_1385),
.B(n_1472),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_1443),
.B(n_1528),
.Y(n_2261)
);

INVx1_ASAP7_75t_SL g2262 ( 
.A(n_1445),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1469),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_1475),
.B(n_1501),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1398),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_1418),
.B(n_1448),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_1361),
.B(n_1379),
.Y(n_2267)
);

NAND3xp33_ASAP7_75t_L g2268 ( 
.A(n_1477),
.B(n_1479),
.C(n_1482),
.Y(n_2268)
);

INVx8_ASAP7_75t_L g2269 ( 
.A(n_1500),
.Y(n_2269)
);

INVx2_ASAP7_75t_SL g2270 ( 
.A(n_1393),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1406),
.B(n_1226),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1478),
.Y(n_2272)
);

INVx3_ASAP7_75t_L g2273 ( 
.A(n_1337),
.Y(n_2273)
);

NAND3xp33_ASAP7_75t_L g2274 ( 
.A(n_1220),
.B(n_1244),
.C(n_762),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1478),
.Y(n_2278)
);

AOI22xp5_ASAP7_75t_L g2279 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1661),
.Y(n_2283)
);

OAI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_1220),
.A2(n_1237),
.B1(n_1226),
.B2(n_1776),
.Y(n_2284)
);

NAND2x1p5_ASAP7_75t_L g2285 ( 
.A(n_1337),
.B(n_794),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1478),
.Y(n_2286)
);

BUFx6f_ASAP7_75t_L g2287 ( 
.A(n_1337),
.Y(n_2287)
);

INVx3_ASAP7_75t_L g2288 ( 
.A(n_1337),
.Y(n_2288)
);

OAI22xp33_ASAP7_75t_L g2289 ( 
.A1(n_1254),
.A2(n_762),
.B1(n_547),
.B2(n_673),
.Y(n_2289)
);

NOR2x1p5_ASAP7_75t_L g2290 ( 
.A(n_1280),
.B(n_1283),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1661),
.Y(n_2292)
);

INVxp67_ASAP7_75t_SL g2293 ( 
.A(n_1430),
.Y(n_2293)
);

AOI22xp33_ASAP7_75t_L g2294 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2294)
);

INVx2_ASAP7_75t_SL g2295 ( 
.A(n_1286),
.Y(n_2295)
);

INVx3_ASAP7_75t_L g2296 ( 
.A(n_1337),
.Y(n_2296)
);

AOI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_SL g2299 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2299)
);

INVx2_ASAP7_75t_SL g2300 ( 
.A(n_1286),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2303)
);

AOI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_1310),
.A2(n_1794),
.B(n_1776),
.Y(n_2304)
);

AOI22xp33_ASAP7_75t_L g2305 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2305)
);

A2O1A1Ixp33_ASAP7_75t_SL g2306 ( 
.A1(n_1545),
.A2(n_1589),
.B(n_1618),
.C(n_1552),
.Y(n_2306)
);

NOR2xp33_ASAP7_75t_L g2307 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2308)
);

BUFx2_ASAP7_75t_L g2309 ( 
.A(n_1666),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1478),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2312)
);

BUFx6f_ASAP7_75t_L g2313 ( 
.A(n_1337),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2314)
);

BUFx3_ASAP7_75t_L g2315 ( 
.A(n_1286),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_SL g2316 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2316)
);

AOI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2317)
);

AOI22xp5_ASAP7_75t_L g2318 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2319)
);

OAI22xp33_ASAP7_75t_L g2320 ( 
.A1(n_1254),
.A2(n_762),
.B1(n_547),
.B2(n_673),
.Y(n_2320)
);

INVx2_ASAP7_75t_SL g2321 ( 
.A(n_1286),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2322)
);

A2O1A1Ixp33_ASAP7_75t_L g2323 ( 
.A1(n_1226),
.A2(n_762),
.B(n_1220),
.C(n_1776),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_1603),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_1661),
.Y(n_2325)
);

NOR2xp67_ASAP7_75t_L g2326 ( 
.A(n_1273),
.B(n_1362),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_SL g2328 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2329)
);

NOR3xp33_ASAP7_75t_SL g2330 ( 
.A(n_1300),
.B(n_1053),
.C(n_440),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1478),
.Y(n_2332)
);

AO22x1_ASAP7_75t_L g2333 ( 
.A1(n_1276),
.A2(n_433),
.B1(n_440),
.B2(n_1296),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_1661),
.Y(n_2334)
);

A2O1A1Ixp33_ASAP7_75t_SL g2335 ( 
.A1(n_1545),
.A2(n_1589),
.B(n_1618),
.C(n_1552),
.Y(n_2335)
);

AND2x6_ASAP7_75t_SL g2336 ( 
.A(n_1244),
.B(n_797),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_L g2338 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2338)
);

AOI21x1_ASAP7_75t_L g2339 ( 
.A1(n_1543),
.A2(n_1028),
.B(n_1026),
.Y(n_2339)
);

AOI22xp33_ASAP7_75t_L g2340 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2340)
);

AND2x6_ASAP7_75t_L g2341 ( 
.A(n_1337),
.B(n_1283),
.Y(n_2341)
);

INVxp67_ASAP7_75t_L g2342 ( 
.A(n_1377),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_1661),
.Y(n_2343)
);

AOI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2344)
);

NAND2xp33_ASAP7_75t_SL g2345 ( 
.A(n_1603),
.B(n_1605),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_1661),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_1661),
.Y(n_2347)
);

AND2x4_ASAP7_75t_SL g2348 ( 
.A(n_1337),
.B(n_1239),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_1478),
.Y(n_2352)
);

BUFx6f_ASAP7_75t_L g2353 ( 
.A(n_1337),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2354)
);

BUFx3_ASAP7_75t_L g2355 ( 
.A(n_1286),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1478),
.Y(n_2356)
);

OAI22xp5_ASAP7_75t_L g2357 ( 
.A1(n_1220),
.A2(n_1237),
.B1(n_1226),
.B2(n_1776),
.Y(n_2357)
);

O2A1O1Ixp5_ASAP7_75t_L g2358 ( 
.A1(n_1220),
.A2(n_1568),
.B(n_1573),
.C(n_1561),
.Y(n_2358)
);

OAI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_1220),
.A2(n_1237),
.B1(n_1226),
.B2(n_1776),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_1661),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2361)
);

AND2x4_ASAP7_75t_L g2362 ( 
.A(n_1273),
.B(n_1283),
.Y(n_2362)
);

AOI22xp33_ASAP7_75t_L g2363 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2363)
);

INVx2_ASAP7_75t_SL g2364 ( 
.A(n_1286),
.Y(n_2364)
);

NAND3xp33_ASAP7_75t_L g2365 ( 
.A(n_1220),
.B(n_1244),
.C(n_762),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_1478),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2369)
);

BUFx5_ASAP7_75t_L g2370 ( 
.A(n_1555),
.Y(n_2370)
);

AOI22xp33_ASAP7_75t_L g2371 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_1478),
.Y(n_2372)
);

INVx2_ASAP7_75t_SL g2373 ( 
.A(n_1286),
.Y(n_2373)
);

INVx8_ASAP7_75t_L g2374 ( 
.A(n_1555),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_1478),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2376)
);

INVx2_ASAP7_75t_SL g2377 ( 
.A(n_1286),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_1478),
.Y(n_2379)
);

AOI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_1478),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2385)
);

AND2x4_ASAP7_75t_L g2386 ( 
.A(n_1273),
.B(n_1283),
.Y(n_2386)
);

OR2x6_ASAP7_75t_L g2387 ( 
.A(n_1337),
.B(n_1310),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_1661),
.Y(n_2388)
);

OR2x2_ASAP7_75t_L g2389 ( 
.A(n_1310),
.B(n_1220),
.Y(n_2389)
);

NAND3xp33_ASAP7_75t_L g2390 ( 
.A(n_1220),
.B(n_1244),
.C(n_762),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2392)
);

AOI22xp5_ASAP7_75t_L g2393 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2394)
);

INVx8_ASAP7_75t_L g2395 ( 
.A(n_1555),
.Y(n_2395)
);

OAI22xp33_ASAP7_75t_L g2396 ( 
.A1(n_1254),
.A2(n_762),
.B1(n_547),
.B2(n_673),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1478),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2398)
);

AOI22xp5_ASAP7_75t_L g2399 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_1478),
.Y(n_2400)
);

NOR2xp33_ASAP7_75t_L g2401 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1478),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_1478),
.Y(n_2404)
);

NOR2xp33_ASAP7_75t_L g2405 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2407)
);

OR2x2_ASAP7_75t_L g2408 ( 
.A(n_1310),
.B(n_1220),
.Y(n_2408)
);

NOR2xp33_ASAP7_75t_L g2409 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_1661),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2411)
);

AOI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_1478),
.Y(n_2414)
);

INVx2_ASAP7_75t_SL g2415 ( 
.A(n_1286),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2416)
);

NOR2xp33_ASAP7_75t_L g2417 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2419)
);

HB1xp67_ASAP7_75t_L g2420 ( 
.A(n_1642),
.Y(n_2420)
);

INVx3_ASAP7_75t_L g2421 ( 
.A(n_1337),
.Y(n_2421)
);

INVx2_ASAP7_75t_SL g2422 ( 
.A(n_1286),
.Y(n_2422)
);

CKINVDCx20_ASAP7_75t_R g2423 ( 
.A(n_1635),
.Y(n_2423)
);

INVx2_ASAP7_75t_SL g2424 ( 
.A(n_1286),
.Y(n_2424)
);

INVxp67_ASAP7_75t_L g2425 ( 
.A(n_1377),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_1478),
.Y(n_2427)
);

BUFx3_ASAP7_75t_L g2428 ( 
.A(n_1286),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_1661),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2432)
);

OR2x6_ASAP7_75t_L g2433 ( 
.A(n_1337),
.B(n_1310),
.Y(n_2433)
);

NAND2x1p5_ASAP7_75t_L g2434 ( 
.A(n_1337),
.B(n_794),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_1478),
.Y(n_2436)
);

OAI22xp5_ASAP7_75t_SL g2437 ( 
.A1(n_1244),
.A2(n_1245),
.B1(n_1256),
.B2(n_1254),
.Y(n_2437)
);

O2A1O1Ixp5_ASAP7_75t_L g2438 ( 
.A1(n_1220),
.A2(n_1568),
.B(n_1573),
.C(n_1561),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_1661),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_SL g2441 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2441)
);

AOI22xp5_ASAP7_75t_L g2442 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_1478),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_1661),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_SL g2449 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_1478),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2451)
);

OR2x2_ASAP7_75t_L g2452 ( 
.A(n_1310),
.B(n_1220),
.Y(n_2452)
);

AOI22xp5_ASAP7_75t_L g2453 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_1478),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_1661),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_SL g2457 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_1478),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2460)
);

NAND3xp33_ASAP7_75t_SL g2461 ( 
.A(n_1220),
.B(n_762),
.C(n_440),
.Y(n_2461)
);

INVx1_ASAP7_75t_SL g2462 ( 
.A(n_1721),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_L g2466 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_L g2467 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_SL g2469 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2469)
);

NOR2xp33_ASAP7_75t_L g2470 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2470)
);

AND2x6_ASAP7_75t_SL g2471 ( 
.A(n_1244),
.B(n_797),
.Y(n_2471)
);

HB1xp67_ASAP7_75t_L g2472 ( 
.A(n_1642),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_1661),
.Y(n_2473)
);

BUFx6f_ASAP7_75t_L g2474 ( 
.A(n_1337),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_1478),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_L g2478 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2481)
);

AOI22xp5_ASAP7_75t_L g2482 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_1661),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2484)
);

AOI22xp33_ASAP7_75t_L g2485 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2486)
);

INVx2_ASAP7_75t_SL g2487 ( 
.A(n_1286),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_1661),
.Y(n_2488)
);

NOR3xp33_ASAP7_75t_L g2489 ( 
.A(n_1220),
.B(n_749),
.C(n_805),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_1478),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_1661),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2494)
);

INVxp67_ASAP7_75t_L g2495 ( 
.A(n_1377),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_SL g2496 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2496)
);

AND2x6_ASAP7_75t_SL g2497 ( 
.A(n_1244),
.B(n_797),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_1661),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_1478),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_1661),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_SL g2506 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_1478),
.Y(n_2507)
);

OR2x6_ASAP7_75t_L g2508 ( 
.A(n_1337),
.B(n_1310),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_SL g2510 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2510)
);

AND2x6_ASAP7_75t_SL g2511 ( 
.A(n_1244),
.B(n_797),
.Y(n_2511)
);

AND2x2_ASAP7_75t_SL g2512 ( 
.A(n_1636),
.B(n_1538),
.Y(n_2512)
);

INVxp67_ASAP7_75t_SL g2513 ( 
.A(n_1430),
.Y(n_2513)
);

AND2x6_ASAP7_75t_L g2514 ( 
.A(n_1337),
.B(n_1283),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_1478),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_SL g2517 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2517)
);

AOI22xp33_ASAP7_75t_L g2518 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2518)
);

AOI22xp33_ASAP7_75t_L g2519 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2519)
);

BUFx3_ASAP7_75t_L g2520 ( 
.A(n_1286),
.Y(n_2520)
);

OR2x2_ASAP7_75t_L g2521 ( 
.A(n_1310),
.B(n_1220),
.Y(n_2521)
);

INVx3_ASAP7_75t_L g2522 ( 
.A(n_1337),
.Y(n_2522)
);

INVx2_ASAP7_75t_SL g2523 ( 
.A(n_1286),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_1478),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2525)
);

AOI22xp33_ASAP7_75t_L g2526 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_1478),
.Y(n_2527)
);

BUFx3_ASAP7_75t_L g2528 ( 
.A(n_1286),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_1478),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_SL g2531 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2532)
);

O2A1O1Ixp5_ASAP7_75t_L g2533 ( 
.A1(n_1220),
.A2(n_1568),
.B(n_1573),
.C(n_1561),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2534)
);

O2A1O1Ixp33_ASAP7_75t_L g2535 ( 
.A1(n_1220),
.A2(n_705),
.B(n_729),
.C(n_678),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_1478),
.Y(n_2536)
);

AOI22xp33_ASAP7_75t_L g2537 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2537)
);

OAI22xp5_ASAP7_75t_L g2538 ( 
.A1(n_1220),
.A2(n_1237),
.B1(n_1226),
.B2(n_1776),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_L g2539 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2539)
);

OR2x2_ASAP7_75t_L g2540 ( 
.A(n_1310),
.B(n_1220),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_1661),
.Y(n_2542)
);

NAND2xp33_ASAP7_75t_L g2543 ( 
.A(n_1224),
.B(n_433),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_SL g2545 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_1478),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_1478),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_1478),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_1661),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_1478),
.Y(n_2552)
);

INVx1_ASAP7_75t_SL g2553 ( 
.A(n_1721),
.Y(n_2553)
);

NAND2x1_ASAP7_75t_L g2554 ( 
.A(n_1542),
.B(n_1273),
.Y(n_2554)
);

BUFx6f_ASAP7_75t_L g2555 ( 
.A(n_1337),
.Y(n_2555)
);

O2A1O1Ixp33_ASAP7_75t_L g2556 ( 
.A1(n_1220),
.A2(n_705),
.B(n_729),
.C(n_678),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2557)
);

BUFx6f_ASAP7_75t_L g2558 ( 
.A(n_1337),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2559)
);

NAND2xp33_ASAP7_75t_L g2560 ( 
.A(n_1224),
.B(n_433),
.Y(n_2560)
);

INVx1_ASAP7_75t_SL g2561 ( 
.A(n_1721),
.Y(n_2561)
);

NOR2x2_ASAP7_75t_L g2562 ( 
.A(n_1285),
.B(n_797),
.Y(n_2562)
);

INVx2_ASAP7_75t_SL g2563 ( 
.A(n_1286),
.Y(n_2563)
);

NOR2x1p5_ASAP7_75t_L g2564 ( 
.A(n_1280),
.B(n_1283),
.Y(n_2564)
);

AOI22xp33_ASAP7_75t_L g2565 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_1478),
.Y(n_2567)
);

AOI22xp5_ASAP7_75t_L g2568 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_L g2569 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2569)
);

O2A1O1Ixp5_ASAP7_75t_L g2570 ( 
.A1(n_1220),
.A2(n_1568),
.B(n_1573),
.C(n_1561),
.Y(n_2570)
);

OR2x2_ASAP7_75t_L g2571 ( 
.A(n_1310),
.B(n_1220),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_1478),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_1478),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_1478),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_1661),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_1478),
.Y(n_2577)
);

O2A1O1Ixp5_ASAP7_75t_L g2578 ( 
.A1(n_1220),
.A2(n_1568),
.B(n_1573),
.C(n_1561),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_SL g2579 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2579)
);

BUFx3_ASAP7_75t_L g2580 ( 
.A(n_1286),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_1603),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_1478),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2584)
);

AOI21xp5_ASAP7_75t_L g2585 ( 
.A1(n_1310),
.A2(n_1794),
.B(n_1776),
.Y(n_2585)
);

NOR2xp33_ASAP7_75t_L g2586 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_SL g2587 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2587)
);

A2O1A1Ixp33_ASAP7_75t_L g2588 ( 
.A1(n_1226),
.A2(n_762),
.B(n_1220),
.C(n_1776),
.Y(n_2588)
);

INVx2_ASAP7_75t_SL g2589 ( 
.A(n_1286),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_1478),
.Y(n_2592)
);

AOI22xp33_ASAP7_75t_SL g2593 ( 
.A1(n_1636),
.A2(n_943),
.B1(n_835),
.B2(n_1311),
.Y(n_2593)
);

INVx8_ASAP7_75t_L g2594 ( 
.A(n_1555),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_SL g2595 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_1478),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_1661),
.Y(n_2597)
);

AOI22xp33_ASAP7_75t_L g2598 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2598)
);

AND2x4_ASAP7_75t_L g2599 ( 
.A(n_1273),
.B(n_1283),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2600)
);

INVx2_ASAP7_75t_SL g2601 ( 
.A(n_1286),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_SL g2602 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_1478),
.Y(n_2603)
);

NOR2xp33_ASAP7_75t_L g2604 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_1661),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_1661),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_1661),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_1478),
.Y(n_2611)
);

AOI22xp33_ASAP7_75t_L g2612 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2612)
);

AOI22xp5_ASAP7_75t_L g2613 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2613)
);

AOI22xp33_ASAP7_75t_L g2614 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2615)
);

AOI22xp33_ASAP7_75t_L g2616 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2616)
);

NOR2xp67_ASAP7_75t_SL g2617 ( 
.A(n_1220),
.B(n_1337),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_1603),
.Y(n_2619)
);

OR2x2_ASAP7_75t_L g2620 ( 
.A(n_1310),
.B(n_1220),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2622)
);

INVx2_ASAP7_75t_SL g2623 ( 
.A(n_1286),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_1478),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_1661),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_1661),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_L g2629 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2630)
);

AOI22xp5_ASAP7_75t_L g2631 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2631)
);

AO22x1_ASAP7_75t_L g2632 ( 
.A1(n_1276),
.A2(n_433),
.B1(n_440),
.B2(n_1296),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_1478),
.Y(n_2633)
);

INVx2_ASAP7_75t_SL g2634 ( 
.A(n_1286),
.Y(n_2634)
);

OAI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_1220),
.A2(n_1237),
.B1(n_1226),
.B2(n_1776),
.Y(n_2635)
);

AOI22xp5_ASAP7_75t_L g2636 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2636)
);

NOR2xp33_ASAP7_75t_L g2637 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2638)
);

NOR2xp33_ASAP7_75t_L g2639 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2641)
);

INVx2_ASAP7_75t_SL g2642 ( 
.A(n_1286),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_SL g2643 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_SL g2644 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_SL g2645 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2645)
);

INVx3_ASAP7_75t_L g2646 ( 
.A(n_1337),
.Y(n_2646)
);

NOR2xp33_ASAP7_75t_L g2647 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2647)
);

AOI22xp33_ASAP7_75t_L g2648 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2648)
);

AOI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2649)
);

HB1xp67_ASAP7_75t_L g2650 ( 
.A(n_1642),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_SL g2652 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2652)
);

OAI21xp5_ASAP7_75t_L g2653 ( 
.A1(n_1220),
.A2(n_1794),
.B(n_1776),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_L g2655 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_1661),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2657)
);

AOI22xp33_ASAP7_75t_L g2658 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2658)
);

AOI22xp5_ASAP7_75t_L g2659 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2659)
);

INVxp67_ASAP7_75t_L g2660 ( 
.A(n_1377),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_1661),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2662)
);

A2O1A1Ixp33_ASAP7_75t_SL g2663 ( 
.A1(n_1545),
.A2(n_1589),
.B(n_1618),
.C(n_1552),
.Y(n_2663)
);

INVx1_ASAP7_75t_SL g2664 ( 
.A(n_1721),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_SL g2665 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2665)
);

AOI22xp5_ASAP7_75t_L g2666 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2666)
);

AND2x2_ASAP7_75t_L g2667 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2668)
);

O2A1O1Ixp33_ASAP7_75t_L g2669 ( 
.A1(n_1220),
.A2(n_705),
.B(n_729),
.C(n_678),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_SL g2670 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2670)
);

INVx2_ASAP7_75t_SL g2671 ( 
.A(n_1286),
.Y(n_2671)
);

NAND2x1p5_ASAP7_75t_L g2672 ( 
.A(n_1337),
.B(n_794),
.Y(n_2672)
);

AND2x6_ASAP7_75t_SL g2673 ( 
.A(n_1244),
.B(n_797),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2674)
);

OR2x6_ASAP7_75t_L g2675 ( 
.A(n_1337),
.B(n_1310),
.Y(n_2675)
);

NOR2xp33_ASAP7_75t_L g2676 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2676)
);

AOI22xp5_ASAP7_75t_L g2677 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2677)
);

AND2x4_ASAP7_75t_L g2678 ( 
.A(n_1273),
.B(n_1283),
.Y(n_2678)
);

AOI22xp33_ASAP7_75t_L g2679 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2679)
);

INVxp67_ASAP7_75t_L g2680 ( 
.A(n_1377),
.Y(n_2680)
);

NOR2xp33_ASAP7_75t_L g2681 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2681)
);

INVx3_ASAP7_75t_L g2682 ( 
.A(n_1337),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_1478),
.Y(n_2683)
);

AOI22xp5_ASAP7_75t_L g2684 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2684)
);

NOR2xp33_ASAP7_75t_L g2685 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2686)
);

BUFx4f_ASAP7_75t_L g2687 ( 
.A(n_1337),
.Y(n_2687)
);

BUFx6f_ASAP7_75t_L g2688 ( 
.A(n_1337),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_SL g2689 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_L g2691 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2691)
);

NOR2xp33_ASAP7_75t_L g2692 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_1478),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_1478),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2695)
);

NOR3xp33_ASAP7_75t_L g2696 ( 
.A(n_1220),
.B(n_749),
.C(n_805),
.Y(n_2696)
);

AND3x1_ASAP7_75t_L g2697 ( 
.A(n_1804),
.B(n_1121),
.C(n_1036),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2699)
);

BUFx3_ASAP7_75t_L g2700 ( 
.A(n_1286),
.Y(n_2700)
);

AND2x6_ASAP7_75t_SL g2701 ( 
.A(n_1244),
.B(n_797),
.Y(n_2701)
);

INVx2_ASAP7_75t_SL g2702 ( 
.A(n_1286),
.Y(n_2702)
);

AOI21xp5_ASAP7_75t_L g2703 ( 
.A1(n_1310),
.A2(n_1794),
.B(n_1776),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2704)
);

NOR3xp33_ASAP7_75t_SL g2705 ( 
.A(n_1300),
.B(n_1053),
.C(n_440),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_1478),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_1661),
.Y(n_2708)
);

INVx3_ASAP7_75t_L g2709 ( 
.A(n_1337),
.Y(n_2709)
);

INVxp67_ASAP7_75t_L g2710 ( 
.A(n_1377),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_1478),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_SL g2714 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2714)
);

INVx2_ASAP7_75t_SL g2715 ( 
.A(n_1286),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2716)
);

AOI22xp33_ASAP7_75t_L g2717 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_1661),
.Y(n_2719)
);

INVxp67_ASAP7_75t_L g2720 ( 
.A(n_1377),
.Y(n_2720)
);

BUFx6f_ASAP7_75t_L g2721 ( 
.A(n_1337),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2723)
);

NOR2xp33_ASAP7_75t_L g2724 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_1661),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_1478),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_1661),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_1478),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_SL g2729 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_1478),
.Y(n_2730)
);

AOI22xp5_ASAP7_75t_L g2731 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2731)
);

AOI22xp33_ASAP7_75t_L g2732 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2732)
);

OR2x6_ASAP7_75t_L g2733 ( 
.A(n_1337),
.B(n_1310),
.Y(n_2733)
);

O2A1O1Ixp5_ASAP7_75t_L g2734 ( 
.A1(n_1220),
.A2(n_1568),
.B(n_1573),
.C(n_1561),
.Y(n_2734)
);

NOR3xp33_ASAP7_75t_L g2735 ( 
.A(n_1220),
.B(n_749),
.C(n_805),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_1478),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2737)
);

OR2x2_ASAP7_75t_L g2738 ( 
.A(n_1310),
.B(n_1220),
.Y(n_2738)
);

A2O1A1Ixp33_ASAP7_75t_L g2739 ( 
.A1(n_1226),
.A2(n_762),
.B(n_1220),
.C(n_1776),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2740)
);

AOI22xp33_ASAP7_75t_L g2741 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2741)
);

AOI22xp33_ASAP7_75t_L g2742 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_1661),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_1478),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_SL g2746 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2746)
);

CKINVDCx5p33_ASAP7_75t_R g2747 ( 
.A(n_1603),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2748)
);

HB1xp67_ASAP7_75t_L g2749 ( 
.A(n_1642),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2751)
);

O2A1O1Ixp33_ASAP7_75t_L g2752 ( 
.A1(n_1220),
.A2(n_705),
.B(n_729),
.C(n_678),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_1478),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_1661),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2755)
);

AOI22xp5_ASAP7_75t_L g2756 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2756)
);

AND2x2_ASAP7_75t_SL g2757 ( 
.A(n_1636),
.B(n_1538),
.Y(n_2757)
);

AOI22xp5_ASAP7_75t_L g2758 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_1661),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_1661),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_1661),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_1661),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_L g2764 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_1661),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_SL g2770 ( 
.A(n_1237),
.B(n_1245),
.Y(n_2770)
);

BUFx5_ASAP7_75t_L g2771 ( 
.A(n_1555),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_1661),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_1478),
.Y(n_2773)
);

NAND2xp33_ASAP7_75t_L g2774 ( 
.A(n_1224),
.B(n_433),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2775)
);

AOI22xp33_ASAP7_75t_L g2776 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2776)
);

NOR2xp33_ASAP7_75t_L g2777 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2777)
);

OR2x2_ASAP7_75t_L g2778 ( 
.A(n_1310),
.B(n_1220),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2779)
);

AND2x4_ASAP7_75t_L g2780 ( 
.A(n_1273),
.B(n_1283),
.Y(n_2780)
);

BUFx3_ASAP7_75t_L g2781 ( 
.A(n_1286),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_1478),
.Y(n_2782)
);

INVx2_ASAP7_75t_SL g2783 ( 
.A(n_1286),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2784)
);

AOI22xp33_ASAP7_75t_L g2785 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_1776),
.B(n_1794),
.Y(n_2786)
);

AND2x4_ASAP7_75t_L g2787 ( 
.A(n_1273),
.B(n_1283),
.Y(n_2787)
);

NOR2xp33_ASAP7_75t_L g2788 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2788)
);

BUFx6f_ASAP7_75t_L g2789 ( 
.A(n_1337),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2790)
);

AOI22xp33_ASAP7_75t_L g2791 ( 
.A1(n_1311),
.A2(n_1634),
.B1(n_1614),
.B2(n_412),
.Y(n_2791)
);

OAI22xp33_ASAP7_75t_L g2792 ( 
.A1(n_1254),
.A2(n_762),
.B1(n_547),
.B2(n_673),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_1478),
.Y(n_2793)
);

AOI22xp5_ASAP7_75t_L g2794 ( 
.A1(n_1220),
.A2(n_1564),
.B1(n_1582),
.B2(n_1575),
.Y(n_2794)
);

BUFx3_ASAP7_75t_L g2795 ( 
.A(n_1286),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_1661),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_1226),
.B(n_1564),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_1478),
.Y(n_2800)
);

INVx8_ASAP7_75t_L g2801 ( 
.A(n_1555),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_L g2802 ( 
.A(n_1254),
.B(n_1256),
.Y(n_2802)
);

A2O1A1Ixp33_ASAP7_75t_L g2803 ( 
.A1(n_1226),
.A2(n_762),
.B(n_1220),
.C(n_1776),
.Y(n_2803)
);

NAND2x1p5_ASAP7_75t_L g2804 ( 
.A(n_1337),
.B(n_794),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_1661),
.Y(n_2805)
);

A2O1A1Ixp33_ASAP7_75t_L g2806 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_2806)
);

OAI21xp5_ASAP7_75t_L g2807 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_2807)
);

AOI21xp5_ASAP7_75t_L g2808 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_2808)
);

NOR2xp33_ASAP7_75t_L g2809 ( 
.A(n_1896),
.B(n_1886),
.Y(n_2809)
);

AOI21x1_ASAP7_75t_L g2810 ( 
.A1(n_2254),
.A2(n_1890),
.B(n_2554),
.Y(n_2810)
);

AOI21xp5_ASAP7_75t_L g2811 ( 
.A1(n_1882),
.A2(n_2357),
.B(n_2284),
.Y(n_2811)
);

CKINVDCx20_ASAP7_75t_R g2812 ( 
.A(n_1905),
.Y(n_2812)
);

CKINVDCx20_ASAP7_75t_R g2813 ( 
.A(n_2423),
.Y(n_2813)
);

AOI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_1882),
.A2(n_2538),
.B(n_2359),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2045),
.B(n_1879),
.Y(n_2815)
);

INVx3_ASAP7_75t_L g2816 ( 
.A(n_2554),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2136),
.Y(n_2817)
);

AOI21xp5_ASAP7_75t_L g2818 ( 
.A1(n_2538),
.A2(n_2635),
.B(n_1910),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2045),
.B(n_1879),
.Y(n_2819)
);

AOI21xp5_ASAP7_75t_L g2820 ( 
.A1(n_2635),
.A2(n_2588),
.B(n_2323),
.Y(n_2820)
);

AOI21xp5_ASAP7_75t_L g2821 ( 
.A1(n_2739),
.A2(n_2803),
.B(n_2653),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_1878),
.B(n_1897),
.Y(n_2822)
);

INVx3_ASAP7_75t_L g2823 ( 
.A(n_1945),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_1881),
.B(n_1888),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_1881),
.B(n_1888),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_1891),
.B(n_1923),
.Y(n_2826)
);

AOI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2653),
.A2(n_2097),
.B(n_2039),
.Y(n_2827)
);

NOR2xp33_ASAP7_75t_L g2828 ( 
.A(n_1886),
.B(n_1861),
.Y(n_2828)
);

AND2x2_ASAP7_75t_L g2829 ( 
.A(n_1878),
.B(n_1897),
.Y(n_2829)
);

AOI21xp5_ASAP7_75t_L g2830 ( 
.A1(n_2097),
.A2(n_1961),
.B(n_1952),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_1891),
.B(n_1923),
.Y(n_2831)
);

AND2x4_ASAP7_75t_L g2832 ( 
.A(n_2362),
.B(n_2386),
.Y(n_2832)
);

O2A1O1Ixp33_ASAP7_75t_L g2833 ( 
.A1(n_2282),
.A2(n_2302),
.B(n_2310),
.C(n_2299),
.Y(n_2833)
);

AOI21x1_ASAP7_75t_L g2834 ( 
.A1(n_2254),
.A2(n_1890),
.B(n_2339),
.Y(n_2834)
);

O2A1O1Ixp33_ASAP7_75t_L g2835 ( 
.A1(n_2312),
.A2(n_2316),
.B(n_2328),
.C(n_2314),
.Y(n_2835)
);

AOI21xp5_ASAP7_75t_L g2836 ( 
.A1(n_2389),
.A2(n_2452),
.B(n_2408),
.Y(n_2836)
);

AOI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2389),
.A2(n_2452),
.B(n_2408),
.Y(n_2837)
);

AOI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2521),
.A2(n_2571),
.B(n_2540),
.Y(n_2838)
);

OAI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2274),
.A2(n_2390),
.B(n_2365),
.Y(n_2839)
);

AOI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_2521),
.A2(n_2571),
.B(n_2540),
.Y(n_2840)
);

AOI21xp5_ASAP7_75t_L g2841 ( 
.A1(n_2620),
.A2(n_2778),
.B(n_2738),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_1925),
.B(n_1926),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2797),
.Y(n_2843)
);

OR2x2_ASAP7_75t_L g2844 ( 
.A(n_1893),
.B(n_2309),
.Y(n_2844)
);

AOI21xp5_ASAP7_75t_L g2845 ( 
.A1(n_2620),
.A2(n_2778),
.B(n_2738),
.Y(n_2845)
);

AOI21xp5_ASAP7_75t_L g2846 ( 
.A1(n_2126),
.A2(n_2383),
.B(n_2337),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_1990),
.B(n_2011),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_1925),
.B(n_1926),
.Y(n_2848)
);

AOI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_2126),
.A2(n_2398),
.B(n_2384),
.Y(n_2849)
);

BUFx6f_ASAP7_75t_L g2850 ( 
.A(n_1914),
.Y(n_2850)
);

AOI21xp5_ASAP7_75t_L g2851 ( 
.A1(n_2406),
.A2(n_2447),
.B(n_2441),
.Y(n_2851)
);

O2A1O1Ixp33_ASAP7_75t_L g2852 ( 
.A1(n_2449),
.A2(n_2469),
.B(n_2496),
.C(n_2457),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_SL g2853 ( 
.A(n_1859),
.B(n_2279),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_1990),
.B(n_2011),
.Y(n_2854)
);

AOI21xp5_ASAP7_75t_L g2855 ( 
.A1(n_2506),
.A2(n_2517),
.B(n_2510),
.Y(n_2855)
);

OAI22xp5_ASAP7_75t_L g2856 ( 
.A1(n_1859),
.A2(n_2317),
.B1(n_2318),
.B2(n_2279),
.Y(n_2856)
);

INVx4_ASAP7_75t_L g2857 ( 
.A(n_1914),
.Y(n_2857)
);

AND2x4_ASAP7_75t_L g2858 ( 
.A(n_2362),
.B(n_2386),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_1874),
.B(n_1876),
.Y(n_2859)
);

AOI21xp5_ASAP7_75t_L g2860 ( 
.A1(n_2525),
.A2(n_2531),
.B(n_2530),
.Y(n_2860)
);

OAI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2274),
.A2(n_2390),
.B(n_2365),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_1874),
.B(n_1876),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_1907),
.B(n_1913),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_1908),
.B(n_1915),
.Y(n_2864)
);

AOI21xp5_ASAP7_75t_L g2865 ( 
.A1(n_2545),
.A2(n_2584),
.B(n_2579),
.Y(n_2865)
);

BUFx6f_ASAP7_75t_L g2866 ( 
.A(n_1914),
.Y(n_2866)
);

OAI21xp5_ASAP7_75t_L g2867 ( 
.A1(n_2587),
.A2(n_2602),
.B(n_2595),
.Y(n_2867)
);

NOR2xp33_ASAP7_75t_L g2868 ( 
.A(n_1863),
.B(n_1864),
.Y(n_2868)
);

A2O1A1Ixp33_ASAP7_75t_L g2869 ( 
.A1(n_2794),
.A2(n_2318),
.B(n_2344),
.C(n_2317),
.Y(n_2869)
);

A2O1A1Ixp33_ASAP7_75t_L g2870 ( 
.A1(n_2344),
.A2(n_2393),
.B(n_2399),
.C(n_2380),
.Y(n_2870)
);

AOI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2615),
.A2(n_2644),
.B(n_2643),
.Y(n_2871)
);

AOI21xp33_ASAP7_75t_L g2872 ( 
.A1(n_2645),
.A2(n_2665),
.B(n_2652),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_1937),
.B(n_1942),
.Y(n_2873)
);

NOR2xp33_ASAP7_75t_L g2874 ( 
.A(n_1867),
.B(n_1871),
.Y(n_2874)
);

BUFx6f_ASAP7_75t_L g2875 ( 
.A(n_1986),
.Y(n_2875)
);

AND2x4_ASAP7_75t_L g2876 ( 
.A(n_2362),
.B(n_2386),
.Y(n_2876)
);

OAI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_2380),
.A2(n_2399),
.B1(n_2442),
.B2(n_2393),
.Y(n_2877)
);

OAI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2442),
.A2(n_2482),
.B1(n_2568),
.B2(n_2453),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2670),
.A2(n_2714),
.B(n_2689),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_1978),
.B(n_1992),
.Y(n_2880)
);

AO21x2_ASAP7_75t_L g2881 ( 
.A1(n_1862),
.A2(n_2283),
.B(n_1866),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_1998),
.B(n_2006),
.Y(n_2882)
);

AOI21xp5_ASAP7_75t_L g2883 ( 
.A1(n_2729),
.A2(n_2766),
.B(n_2746),
.Y(n_2883)
);

AOI21xp5_ASAP7_75t_L g2884 ( 
.A1(n_2770),
.A2(n_2044),
.B(n_2122),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2797),
.Y(n_2885)
);

AOI21xp5_ASAP7_75t_L g2886 ( 
.A1(n_2078),
.A2(n_2091),
.B(n_2079),
.Y(n_2886)
);

OAI21xp5_ASAP7_75t_L g2887 ( 
.A1(n_2453),
.A2(n_2568),
.B(n_2482),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_1875),
.B(n_1877),
.Y(n_2888)
);

AOI21xp5_ASAP7_75t_L g2889 ( 
.A1(n_2093),
.A2(n_1956),
.B(n_1946),
.Y(n_2889)
);

OAI21xp33_ASAP7_75t_L g2890 ( 
.A1(n_2613),
.A2(n_2636),
.B(n_2631),
.Y(n_2890)
);

AOI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_1960),
.A2(n_1968),
.B(n_1962),
.Y(n_2891)
);

AOI21xp5_ASAP7_75t_L g2892 ( 
.A1(n_1970),
.A2(n_1987),
.B(n_1974),
.Y(n_2892)
);

AOI21xp33_ASAP7_75t_L g2893 ( 
.A1(n_2025),
.A2(n_2038),
.B(n_2358),
.Y(n_2893)
);

BUFx6f_ASAP7_75t_L g2894 ( 
.A(n_1986),
.Y(n_2894)
);

NOR2xp33_ASAP7_75t_L g2895 ( 
.A(n_1880),
.B(n_1892),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2010),
.B(n_1965),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_1965),
.B(n_2008),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2805),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_L g2899 ( 
.A(n_1894),
.B(n_1860),
.Y(n_2899)
);

AOI21xp5_ASAP7_75t_L g2900 ( 
.A1(n_1991),
.A2(n_2018),
.B(n_2000),
.Y(n_2900)
);

OAI21xp33_ASAP7_75t_L g2901 ( 
.A1(n_2613),
.A2(n_2636),
.B(n_2631),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2805),
.Y(n_2902)
);

AOI21xp5_ASAP7_75t_L g2903 ( 
.A1(n_2020),
.A2(n_2021),
.B(n_2387),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2127),
.Y(n_2904)
);

AOI21x1_ASAP7_75t_L g2905 ( 
.A1(n_2339),
.A2(n_1883),
.B(n_1869),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2127),
.Y(n_2906)
);

AOI21xp5_ASAP7_75t_L g2907 ( 
.A1(n_2387),
.A2(n_2508),
.B(n_2433),
.Y(n_2907)
);

AOI21xp5_ASAP7_75t_L g2908 ( 
.A1(n_2387),
.A2(n_2508),
.B(n_2433),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_SL g2909 ( 
.A(n_2649),
.B(n_2659),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_SL g2910 ( 
.A(n_2649),
.B(n_2659),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_SL g2911 ( 
.A(n_1920),
.B(n_1986),
.Y(n_2911)
);

AOI21xp5_ASAP7_75t_L g2912 ( 
.A1(n_2387),
.A2(n_2508),
.B(n_2433),
.Y(n_2912)
);

HB1xp67_ASAP7_75t_L g2913 ( 
.A(n_2309),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_1908),
.Y(n_2914)
);

AOI21xp5_ASAP7_75t_L g2915 ( 
.A1(n_2387),
.A2(n_2508),
.B(n_2433),
.Y(n_2915)
);

O2A1O1Ixp33_ASAP7_75t_L g2916 ( 
.A1(n_1898),
.A2(n_2696),
.B(n_2735),
.C(n_2489),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2016),
.B(n_2003),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2016),
.B(n_2003),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_2666),
.B(n_2677),
.Y(n_2919)
);

A2O1A1Ixp33_ASAP7_75t_L g2920 ( 
.A1(n_2794),
.A2(n_2666),
.B(n_2684),
.C(n_2677),
.Y(n_2920)
);

AO21x1_ASAP7_75t_L g2921 ( 
.A1(n_2027),
.A2(n_2280),
.B(n_1868),
.Y(n_2921)
);

BUFx12f_ASAP7_75t_L g2922 ( 
.A(n_1967),
.Y(n_2922)
);

AOI21x1_ASAP7_75t_L g2923 ( 
.A1(n_1883),
.A2(n_2326),
.B(n_1869),
.Y(n_2923)
);

OAI22xp5_ASAP7_75t_L g2924 ( 
.A1(n_2684),
.A2(n_2756),
.B1(n_2758),
.B2(n_2731),
.Y(n_2924)
);

AOI21xp5_ASAP7_75t_L g2925 ( 
.A1(n_2433),
.A2(n_2675),
.B(n_2508),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2008),
.B(n_2048),
.Y(n_2926)
);

OAI21xp5_ASAP7_75t_L g2927 ( 
.A1(n_2731),
.A2(n_2758),
.B(n_2756),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_1870),
.B(n_1873),
.Y(n_2928)
);

AOI21xp5_ASAP7_75t_L g2929 ( 
.A1(n_2675),
.A2(n_2733),
.B(n_1933),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_1908),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_1870),
.B(n_1873),
.Y(n_2931)
);

NOR2xp33_ASAP7_75t_L g2932 ( 
.A(n_2275),
.B(n_2276),
.Y(n_2932)
);

BUFx3_ASAP7_75t_L g2933 ( 
.A(n_2244),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_1915),
.Y(n_2934)
);

AOI21xp5_ASAP7_75t_L g2935 ( 
.A1(n_2675),
.A2(n_2733),
.B(n_1940),
.Y(n_2935)
);

NOR2xp67_ASAP7_75t_L g2936 ( 
.A(n_2190),
.B(n_2326),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2272),
.B(n_2278),
.Y(n_2937)
);

AOI21xp5_ASAP7_75t_L g2938 ( 
.A1(n_2675),
.A2(n_2733),
.B(n_1948),
.Y(n_2938)
);

AOI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2437),
.A2(n_2281),
.B1(n_2291),
.B2(n_2277),
.Y(n_2939)
);

AOI21xp5_ASAP7_75t_L g2940 ( 
.A1(n_2675),
.A2(n_2733),
.B(n_1949),
.Y(n_2940)
);

OAI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2054),
.A2(n_2533),
.B(n_2438),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2272),
.B(n_2278),
.Y(n_2942)
);

AOI21xp5_ASAP7_75t_L g2943 ( 
.A1(n_2733),
.A2(n_1954),
.B(n_1928),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_1915),
.B(n_1958),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_L g2945 ( 
.A(n_2298),
.B(n_2301),
.Y(n_2945)
);

AOI22xp5_ASAP7_75t_L g2946 ( 
.A1(n_2437),
.A2(n_2308),
.B1(n_2319),
.B2(n_2303),
.Y(n_2946)
);

INVx11_ASAP7_75t_L g2947 ( 
.A(n_1976),
.Y(n_2947)
);

AOI21xp5_ASAP7_75t_L g2948 ( 
.A1(n_1971),
.A2(n_1988),
.B(n_1983),
.Y(n_2948)
);

HB1xp67_ASAP7_75t_L g2949 ( 
.A(n_1966),
.Y(n_2949)
);

BUFx8_ASAP7_75t_SL g2950 ( 
.A(n_2225),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_1958),
.Y(n_2951)
);

AND2x2_ASAP7_75t_L g2952 ( 
.A(n_1958),
.B(n_1964),
.Y(n_2952)
);

AOI21xp5_ASAP7_75t_L g2953 ( 
.A1(n_2005),
.A2(n_2280),
.B(n_1868),
.Y(n_2953)
);

INVx3_ASAP7_75t_L g2954 ( 
.A(n_1945),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2286),
.B(n_2311),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2286),
.B(n_2311),
.Y(n_2956)
);

NOR2xp33_ASAP7_75t_L g2957 ( 
.A(n_2322),
.B(n_2329),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_L g2958 ( 
.A(n_2331),
.B(n_2350),
.Y(n_2958)
);

OAI21xp5_ASAP7_75t_L g2959 ( 
.A1(n_2054),
.A2(n_2578),
.B(n_2570),
.Y(n_2959)
);

INVx3_ASAP7_75t_L g2960 ( 
.A(n_1945),
.Y(n_2960)
);

OAI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2734),
.A2(n_2349),
.B(n_2327),
.Y(n_2961)
);

OAI21xp33_ASAP7_75t_L g2962 ( 
.A1(n_2790),
.A2(n_2798),
.B(n_2796),
.Y(n_2962)
);

BUFx4f_ASAP7_75t_L g2963 ( 
.A(n_2801),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2332),
.B(n_2352),
.Y(n_2964)
);

INVx3_ASAP7_75t_L g2965 ( 
.A(n_1945),
.Y(n_2965)
);

AOI21xp5_ASAP7_75t_L g2966 ( 
.A1(n_2327),
.A2(n_2367),
.B(n_2349),
.Y(n_2966)
);

O2A1O1Ixp33_ASAP7_75t_L g2967 ( 
.A1(n_2306),
.A2(n_2663),
.B(n_2335),
.C(n_2042),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2332),
.B(n_2352),
.Y(n_2968)
);

AOI21xp5_ASAP7_75t_L g2969 ( 
.A1(n_2367),
.A2(n_2435),
.B(n_2402),
.Y(n_2969)
);

OAI21xp5_ASAP7_75t_L g2970 ( 
.A1(n_2402),
.A2(n_2439),
.B(n_2435),
.Y(n_2970)
);

AOI21xp5_ASAP7_75t_L g2971 ( 
.A1(n_2439),
.A2(n_2493),
.B(n_2464),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2356),
.B(n_2366),
.Y(n_2972)
);

OAI22xp5_ASAP7_75t_L g2973 ( 
.A1(n_2351),
.A2(n_2361),
.B1(n_2368),
.B2(n_2354),
.Y(n_2973)
);

OAI22xp5_ASAP7_75t_L g2974 ( 
.A1(n_2376),
.A2(n_2385),
.B1(n_2391),
.B2(n_2381),
.Y(n_2974)
);

BUFx4f_ASAP7_75t_L g2975 ( 
.A(n_2801),
.Y(n_2975)
);

A2O1A1Ixp33_ASAP7_75t_L g2976 ( 
.A1(n_1895),
.A2(n_2068),
.B(n_2052),
.C(n_2461),
.Y(n_2976)
);

AOI22xp5_ASAP7_75t_L g2977 ( 
.A1(n_2392),
.A2(n_2411),
.B1(n_2413),
.B2(n_2407),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_1964),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2356),
.B(n_2366),
.Y(n_2979)
);

AOI21xp5_ASAP7_75t_L g2980 ( 
.A1(n_2464),
.A2(n_2498),
.B(n_2493),
.Y(n_2980)
);

OAI22xp5_ASAP7_75t_L g2981 ( 
.A1(n_2416),
.A2(n_2419),
.B1(n_2426),
.B2(n_2418),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2372),
.B(n_2375),
.Y(n_2982)
);

A2O1A1Ixp33_ASAP7_75t_L g2983 ( 
.A1(n_1885),
.A2(n_2307),
.B(n_2338),
.C(n_1889),
.Y(n_2983)
);

NAND2xp33_ASAP7_75t_L g2984 ( 
.A(n_2430),
.B(n_2431),
.Y(n_2984)
);

NAND3xp33_ASAP7_75t_SL g2985 ( 
.A(n_2432),
.B(n_2445),
.C(n_2444),
.Y(n_2985)
);

OAI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2498),
.A2(n_2566),
.B(n_2549),
.Y(n_2986)
);

BUFx3_ASAP7_75t_L g2987 ( 
.A(n_2244),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2372),
.B(n_2375),
.Y(n_2988)
);

AOI21xp5_ASAP7_75t_L g2989 ( 
.A1(n_2549),
.A2(n_2628),
.B(n_2566),
.Y(n_2989)
);

OAI21xp5_ASAP7_75t_L g2990 ( 
.A1(n_2628),
.A2(n_2667),
.B(n_2641),
.Y(n_2990)
);

NOR2x1p5_ASAP7_75t_SL g2991 ( 
.A(n_1969),
.B(n_2370),
.Y(n_2991)
);

AND2x2_ASAP7_75t_L g2992 ( 
.A(n_1964),
.B(n_1977),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2379),
.B(n_2382),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2379),
.B(n_2382),
.Y(n_2994)
);

HB1xp67_ASAP7_75t_L g2995 ( 
.A(n_2420),
.Y(n_2995)
);

AOI21xp5_ASAP7_75t_L g2996 ( 
.A1(n_2641),
.A2(n_2786),
.B(n_2667),
.Y(n_2996)
);

OAI21xp5_ASAP7_75t_L g2997 ( 
.A1(n_2786),
.A2(n_2451),
.B(n_2448),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_SL g2998 ( 
.A(n_2189),
.B(n_2101),
.Y(n_2998)
);

AND2x2_ASAP7_75t_L g2999 ( 
.A(n_1977),
.B(n_1984),
.Y(n_2999)
);

BUFx3_ASAP7_75t_L g3000 ( 
.A(n_2244),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2397),
.B(n_2400),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_SL g3002 ( 
.A(n_2101),
.B(n_2697),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2397),
.B(n_2400),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2403),
.B(n_2404),
.Y(n_3004)
);

INVx3_ASAP7_75t_L g3005 ( 
.A(n_1945),
.Y(n_3005)
);

AOI21xp5_ASAP7_75t_L g3006 ( 
.A1(n_1900),
.A2(n_1909),
.B(n_1906),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_1977),
.B(n_1984),
.Y(n_3007)
);

AOI21xp5_ASAP7_75t_L g3008 ( 
.A1(n_1912),
.A2(n_1918),
.B(n_1916),
.Y(n_3008)
);

AOI21xp5_ASAP7_75t_L g3009 ( 
.A1(n_1922),
.A2(n_1927),
.B(n_1924),
.Y(n_3009)
);

A2O1A1Ixp33_ASAP7_75t_L g3010 ( 
.A1(n_2369),
.A2(n_2394),
.B(n_2401),
.C(n_2378),
.Y(n_3010)
);

NOR2xp33_ASAP7_75t_L g3011 ( 
.A(n_2456),
.B(n_2459),
.Y(n_3011)
);

AOI21xp5_ASAP7_75t_L g3012 ( 
.A1(n_1935),
.A2(n_1941),
.B(n_1938),
.Y(n_3012)
);

AND2x4_ASAP7_75t_L g3013 ( 
.A(n_2362),
.B(n_2386),
.Y(n_3013)
);

A2O1A1Ixp33_ASAP7_75t_L g3014 ( 
.A1(n_2405),
.A2(n_2417),
.B(n_2466),
.C(n_2409),
.Y(n_3014)
);

OAI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2460),
.A2(n_2465),
.B(n_2463),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2403),
.B(n_2404),
.Y(n_3016)
);

AOI21xp5_ASAP7_75t_L g3017 ( 
.A1(n_2123),
.A2(n_2099),
.B(n_1921),
.Y(n_3017)
);

INVx2_ASAP7_75t_SL g3018 ( 
.A(n_2180),
.Y(n_3018)
);

INVx2_ASAP7_75t_SL g3019 ( 
.A(n_2180),
.Y(n_3019)
);

INVx6_ASAP7_75t_L g3020 ( 
.A(n_2374),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_1984),
.Y(n_3021)
);

NOR2xp33_ASAP7_75t_L g3022 ( 
.A(n_2468),
.B(n_2476),
.Y(n_3022)
);

AOI22xp5_ASAP7_75t_L g3023 ( 
.A1(n_2477),
.A2(n_2481),
.B1(n_2484),
.B2(n_2480),
.Y(n_3023)
);

AOI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_2128),
.A2(n_2490),
.B(n_2486),
.Y(n_3024)
);

BUFx12f_ASAP7_75t_L g3025 ( 
.A(n_1976),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2414),
.B(n_2427),
.Y(n_3026)
);

AOI21xp5_ASAP7_75t_L g3027 ( 
.A1(n_2784),
.A2(n_2799),
.B(n_2499),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2414),
.B(n_2427),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2436),
.B(n_2443),
.Y(n_3029)
);

NOR2xp67_ASAP7_75t_L g3030 ( 
.A(n_1904),
.B(n_1920),
.Y(n_3030)
);

OAI22xp5_ASAP7_75t_L g3031 ( 
.A1(n_2494),
.A2(n_2502),
.B1(n_2504),
.B2(n_2501),
.Y(n_3031)
);

OAI21xp5_ASAP7_75t_L g3032 ( 
.A1(n_2509),
.A2(n_2532),
.B(n_2516),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_SL g3033 ( 
.A(n_2697),
.B(n_2534),
.Y(n_3033)
);

INVx2_ASAP7_75t_SL g3034 ( 
.A(n_2180),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_SL g3035 ( 
.A(n_2541),
.B(n_2544),
.Y(n_3035)
);

INVx4_ASAP7_75t_L g3036 ( 
.A(n_1920),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2436),
.B(n_2443),
.Y(n_3037)
);

AOI22xp5_ASAP7_75t_L g3038 ( 
.A1(n_2546),
.A2(n_2581),
.B1(n_2590),
.B2(n_2557),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_SL g3039 ( 
.A(n_2591),
.B(n_2600),
.Y(n_3039)
);

O2A1O1Ixp33_ASAP7_75t_SL g3040 ( 
.A1(n_2608),
.A2(n_2610),
.B(n_2618),
.C(n_2609),
.Y(n_3040)
);

OAI22xp5_ASAP7_75t_L g3041 ( 
.A1(n_2621),
.A2(n_2624),
.B1(n_2630),
.B2(n_2622),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_SL g3042 ( 
.A(n_2638),
.B(n_2640),
.Y(n_3042)
);

AOI22xp5_ASAP7_75t_L g3043 ( 
.A1(n_2651),
.A2(n_2657),
.B1(n_2662),
.B2(n_2654),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2450),
.B(n_2454),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_L g3045 ( 
.A(n_2668),
.B(n_2674),
.Y(n_3045)
);

OAI22xp5_ASAP7_75t_L g3046 ( 
.A1(n_2686),
.A2(n_2695),
.B1(n_2698),
.B2(n_2690),
.Y(n_3046)
);

INVx4_ASAP7_75t_L g3047 ( 
.A(n_1920),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2450),
.B(n_2454),
.Y(n_3048)
);

AOI21xp5_ASAP7_75t_L g3049 ( 
.A1(n_2699),
.A2(n_2706),
.B(n_2704),
.Y(n_3049)
);

OAI21xp5_ASAP7_75t_L g3050 ( 
.A1(n_2711),
.A2(n_2716),
.B(n_2712),
.Y(n_3050)
);

BUFx8_ASAP7_75t_L g3051 ( 
.A(n_2246),
.Y(n_3051)
);

AND2x4_ASAP7_75t_SL g3052 ( 
.A(n_2287),
.B(n_2313),
.Y(n_3052)
);

AOI21xp5_ASAP7_75t_L g3053 ( 
.A1(n_2718),
.A2(n_2723),
.B(n_2722),
.Y(n_3053)
);

AOI21xp5_ASAP7_75t_L g3054 ( 
.A1(n_2740),
.A2(n_2748),
.B(n_2743),
.Y(n_3054)
);

OAI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2750),
.A2(n_2755),
.B(n_2751),
.Y(n_3055)
);

AOI22xp5_ASAP7_75t_L g3056 ( 
.A1(n_2763),
.A2(n_2768),
.B1(n_2769),
.B2(n_2765),
.Y(n_3056)
);

AOI21xp5_ASAP7_75t_L g3057 ( 
.A1(n_2775),
.A2(n_2779),
.B(n_2249),
.Y(n_3057)
);

OAI21xp5_ASAP7_75t_L g3058 ( 
.A1(n_2049),
.A2(n_2059),
.B(n_2802),
.Y(n_3058)
);

BUFx3_ASAP7_75t_L g3059 ( 
.A(n_2244),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2009),
.Y(n_3060)
);

INVxp67_ASAP7_75t_L g3061 ( 
.A(n_2090),
.Y(n_3061)
);

O2A1O1Ixp33_ASAP7_75t_L g3062 ( 
.A1(n_2289),
.A2(n_2320),
.B(n_2792),
.C(n_2396),
.Y(n_3062)
);

AOI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_2249),
.A2(n_2037),
.B(n_2293),
.Y(n_3063)
);

AOI21xp5_ASAP7_75t_L g3064 ( 
.A1(n_2037),
.A2(n_2513),
.B(n_2072),
.Y(n_3064)
);

AOI21xp5_ASAP7_75t_L g3065 ( 
.A1(n_1904),
.A2(n_2757),
.B(n_2512),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_SL g3066 ( 
.A(n_1902),
.B(n_2112),
.Y(n_3066)
);

AOI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_1904),
.A2(n_2757),
.B(n_2512),
.Y(n_3067)
);

INVx3_ASAP7_75t_L g3068 ( 
.A(n_1945),
.Y(n_3068)
);

AOI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2512),
.A2(n_2757),
.B(n_2560),
.Y(n_3069)
);

AOI21xp5_ASAP7_75t_L g3070 ( 
.A1(n_2774),
.A2(n_2543),
.B(n_2243),
.Y(n_3070)
);

AOI21xp5_ASAP7_75t_L g3071 ( 
.A1(n_2252),
.A2(n_2255),
.B(n_2195),
.Y(n_3071)
);

BUFx8_ASAP7_75t_L g3072 ( 
.A(n_2246),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2458),
.B(n_2475),
.Y(n_3073)
);

CKINVDCx20_ASAP7_75t_R g3074 ( 
.A(n_1957),
.Y(n_3074)
);

AOI21xp5_ASAP7_75t_L g3075 ( 
.A1(n_2234),
.A2(n_2678),
.B(n_2599),
.Y(n_3075)
);

AOI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_2234),
.A2(n_2678),
.B(n_2599),
.Y(n_3076)
);

BUFx8_ASAP7_75t_SL g3077 ( 
.A(n_2225),
.Y(n_3077)
);

A2O1A1Ixp33_ASAP7_75t_L g3078 ( 
.A1(n_2467),
.A2(n_2470),
.B(n_2479),
.C(n_2478),
.Y(n_3078)
);

BUFx6f_ASAP7_75t_L g3079 ( 
.A(n_2374),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2009),
.Y(n_3080)
);

AOI21xp5_ASAP7_75t_L g3081 ( 
.A1(n_2234),
.A2(n_2678),
.B(n_2599),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_SL g3082 ( 
.A(n_2069),
.B(n_1934),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2458),
.B(n_2475),
.Y(n_3083)
);

OAI21xp33_ASAP7_75t_L g3084 ( 
.A1(n_2539),
.A2(n_2569),
.B(n_2559),
.Y(n_3084)
);

BUFx8_ASAP7_75t_L g3085 ( 
.A(n_2246),
.Y(n_3085)
);

OAI21xp5_ASAP7_75t_L g3086 ( 
.A1(n_2573),
.A2(n_2604),
.B(n_2586),
.Y(n_3086)
);

AOI21xp5_ASAP7_75t_L g3087 ( 
.A1(n_2234),
.A2(n_2678),
.B(n_2599),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2491),
.B(n_2503),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2491),
.B(n_2503),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2009),
.Y(n_3090)
);

AOI21xp5_ASAP7_75t_L g3091 ( 
.A1(n_2234),
.A2(n_2787),
.B(n_2780),
.Y(n_3091)
);

O2A1O1Ixp33_ASAP7_75t_L g3092 ( 
.A1(n_2629),
.A2(n_2639),
.B(n_2647),
.C(n_2637),
.Y(n_3092)
);

INVx3_ASAP7_75t_L g3093 ( 
.A(n_1945),
.Y(n_3093)
);

AOI21xp5_ASAP7_75t_L g3094 ( 
.A1(n_2780),
.A2(n_2787),
.B(n_2080),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2507),
.B(n_2515),
.Y(n_3095)
);

BUFx12f_ASAP7_75t_L g3096 ( 
.A(n_1976),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_2507),
.B(n_2515),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2524),
.B(n_2527),
.Y(n_3098)
);

AOI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_2780),
.A2(n_2787),
.B(n_2076),
.Y(n_3099)
);

AOI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2780),
.A2(n_2787),
.B(n_2109),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2015),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2524),
.B(n_2527),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2529),
.B(n_2536),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2529),
.B(n_2536),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_SL g3105 ( 
.A(n_2069),
.B(n_1934),
.Y(n_3105)
);

AND2x4_ASAP7_75t_L g3106 ( 
.A(n_1936),
.B(n_2015),
.Y(n_3106)
);

AOI22xp5_ASAP7_75t_L g3107 ( 
.A1(n_2655),
.A2(n_2681),
.B1(n_2685),
.B2(n_2676),
.Y(n_3107)
);

INVx4_ASAP7_75t_L g3108 ( 
.A(n_2374),
.Y(n_3108)
);

NOR2xp33_ASAP7_75t_L g3109 ( 
.A(n_2691),
.B(n_2692),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2102),
.A2(n_2115),
.B(n_2110),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2547),
.B(n_2548),
.Y(n_3111)
);

NOR2xp33_ASAP7_75t_L g3112 ( 
.A(n_2724),
.B(n_2737),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2547),
.B(n_2548),
.Y(n_3113)
);

BUFx2_ASAP7_75t_L g3114 ( 
.A(n_2089),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_2015),
.B(n_2017),
.Y(n_3115)
);

AND2x2_ASAP7_75t_L g3116 ( 
.A(n_2017),
.B(n_2023),
.Y(n_3116)
);

OAI22xp5_ASAP7_75t_L g3117 ( 
.A1(n_2764),
.A2(n_2788),
.B1(n_2777),
.B2(n_2297),
.Y(n_3117)
);

AOI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_2085),
.A2(n_2632),
.B(n_2333),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_SL g3119 ( 
.A(n_1981),
.B(n_2043),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2017),
.Y(n_3120)
);

NOR3xp33_ASAP7_75t_L g3121 ( 
.A(n_2333),
.B(n_2632),
.C(n_2271),
.Y(n_3121)
);

AOI21xp5_ASAP7_75t_L g3122 ( 
.A1(n_2374),
.A2(n_2594),
.B(n_2395),
.Y(n_3122)
);

AOI21xp5_ASAP7_75t_L g3123 ( 
.A1(n_2374),
.A2(n_2594),
.B(n_2395),
.Y(n_3123)
);

OAI321xp33_ASAP7_75t_L g3124 ( 
.A1(n_2294),
.A2(n_2363),
.A3(n_2305),
.B1(n_2412),
.B2(n_2371),
.C(n_2340),
.Y(n_3124)
);

O2A1O1Ixp33_ASAP7_75t_L g3125 ( 
.A1(n_2155),
.A2(n_2035),
.B(n_2083),
.C(n_2075),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2550),
.B(n_2552),
.Y(n_3126)
);

AOI21xp5_ASAP7_75t_L g3127 ( 
.A1(n_2395),
.A2(n_2801),
.B(n_2594),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2550),
.B(n_2552),
.Y(n_3128)
);

NOR2xp33_ASAP7_75t_L g3129 ( 
.A(n_1858),
.B(n_2342),
.Y(n_3129)
);

O2A1O1Ixp33_ASAP7_75t_L g3130 ( 
.A1(n_2077),
.A2(n_2031),
.B(n_2032),
.C(n_2029),
.Y(n_3130)
);

OAI21xp33_ASAP7_75t_L g3131 ( 
.A1(n_2485),
.A2(n_2519),
.B(n_2518),
.Y(n_3131)
);

HB1xp67_ASAP7_75t_L g3132 ( 
.A(n_2472),
.Y(n_3132)
);

AOI22xp5_ASAP7_75t_L g3133 ( 
.A1(n_2526),
.A2(n_2537),
.B1(n_2598),
.B2(n_2565),
.Y(n_3133)
);

INVx3_ASAP7_75t_L g3134 ( 
.A(n_2180),
.Y(n_3134)
);

A2O1A1Ixp33_ASAP7_75t_L g3135 ( 
.A1(n_2055),
.A2(n_2063),
.B(n_2056),
.C(n_2612),
.Y(n_3135)
);

AOI21xp5_ASAP7_75t_L g3136 ( 
.A1(n_2395),
.A2(n_2801),
.B(n_2594),
.Y(n_3136)
);

NOR2xp33_ASAP7_75t_L g3137 ( 
.A(n_2425),
.B(n_2495),
.Y(n_3137)
);

INVx4_ASAP7_75t_L g3138 ( 
.A(n_2395),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2567),
.B(n_2572),
.Y(n_3139)
);

AND2x2_ASAP7_75t_L g3140 ( 
.A(n_2023),
.B(n_2024),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2567),
.B(n_2572),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2574),
.B(n_2575),
.Y(n_3142)
);

NOR2x1_ASAP7_75t_R g3143 ( 
.A(n_1919),
.B(n_2324),
.Y(n_3143)
);

NOR2xp33_ASAP7_75t_L g3144 ( 
.A(n_2660),
.B(n_2680),
.Y(n_3144)
);

OAI22xp5_ASAP7_75t_L g3145 ( 
.A1(n_2614),
.A2(n_2616),
.B1(n_2658),
.B2(n_2648),
.Y(n_3145)
);

OAI21xp33_ASAP7_75t_L g3146 ( 
.A1(n_2679),
.A2(n_2732),
.B(n_2717),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2023),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_SL g3148 ( 
.A(n_2043),
.B(n_1917),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_SL g3149 ( 
.A(n_1917),
.B(n_1979),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_2574),
.B(n_2575),
.Y(n_3150)
);

INVxp67_ASAP7_75t_L g3151 ( 
.A(n_2033),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2577),
.B(n_2583),
.Y(n_3152)
);

OAI21xp5_ASAP7_75t_L g3153 ( 
.A1(n_1995),
.A2(n_2036),
.B(n_2268),
.Y(n_3153)
);

AOI22xp5_ASAP7_75t_L g3154 ( 
.A1(n_2741),
.A2(n_2742),
.B1(n_2785),
.B2(n_2776),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2577),
.B(n_2583),
.Y(n_3155)
);

AOI21xp5_ASAP7_75t_L g3156 ( 
.A1(n_2594),
.A2(n_2801),
.B(n_2596),
.Y(n_3156)
);

AOI21xp5_ASAP7_75t_L g3157 ( 
.A1(n_2592),
.A2(n_2603),
.B(n_2596),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2024),
.Y(n_3158)
);

AOI21xp5_ASAP7_75t_L g3159 ( 
.A1(n_2592),
.A2(n_2611),
.B(n_2603),
.Y(n_3159)
);

AOI22xp5_ASAP7_75t_L g3160 ( 
.A1(n_2791),
.A2(n_1865),
.B1(n_1899),
.B2(n_1917),
.Y(n_3160)
);

AOI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_2611),
.A2(n_2633),
.B(n_2625),
.Y(n_3161)
);

AOI21xp5_ASAP7_75t_L g3162 ( 
.A1(n_2625),
.A2(n_2683),
.B(n_2633),
.Y(n_3162)
);

NOR2xp67_ASAP7_75t_L g3163 ( 
.A(n_2683),
.B(n_2693),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_SL g3164 ( 
.A(n_2203),
.B(n_2242),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2693),
.B(n_2694),
.Y(n_3165)
);

AOI21xp5_ASAP7_75t_L g3166 ( 
.A1(n_2694),
.A2(n_2713),
.B(n_2707),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_SL g3167 ( 
.A(n_2203),
.B(n_2242),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_SL g3168 ( 
.A(n_2131),
.B(n_2094),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2707),
.B(n_2713),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_2726),
.B(n_2728),
.Y(n_3170)
);

BUFx6f_ASAP7_75t_L g3171 ( 
.A(n_2287),
.Y(n_3171)
);

O2A1O1Ixp33_ASAP7_75t_L g3172 ( 
.A1(n_2650),
.A2(n_2749),
.B(n_2710),
.C(n_2720),
.Y(n_3172)
);

OAI21x1_ASAP7_75t_L g3173 ( 
.A1(n_2292),
.A2(n_2334),
.B(n_2325),
.Y(n_3173)
);

NAND3xp33_ASAP7_75t_L g3174 ( 
.A(n_2617),
.B(n_2084),
.C(n_2268),
.Y(n_3174)
);

AND2x2_ASAP7_75t_L g3175 ( 
.A(n_2024),
.B(n_2034),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2726),
.B(n_2728),
.Y(n_3176)
);

AOI21xp5_ASAP7_75t_L g3177 ( 
.A1(n_2730),
.A2(n_2745),
.B(n_2736),
.Y(n_3177)
);

OAI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_2617),
.A2(n_2104),
.B(n_2125),
.Y(n_3178)
);

INVx3_ASAP7_75t_L g3179 ( 
.A(n_2180),
.Y(n_3179)
);

OAI22xp5_ASAP7_75t_L g3180 ( 
.A1(n_1893),
.A2(n_1932),
.B1(n_2593),
.B2(n_2007),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_2034),
.B(n_2040),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_SL g3182 ( 
.A(n_2132),
.B(n_1950),
.Y(n_3182)
);

AOI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_2730),
.A2(n_2745),
.B(n_2736),
.Y(n_3183)
);

INVx3_ASAP7_75t_L g3184 ( 
.A(n_2180),
.Y(n_3184)
);

AO21x1_ASAP7_75t_L g3185 ( 
.A1(n_2253),
.A2(n_2138),
.B(n_2135),
.Y(n_3185)
);

AOI21xp5_ASAP7_75t_L g3186 ( 
.A1(n_2753),
.A2(n_2782),
.B(n_2773),
.Y(n_3186)
);

O2A1O1Ixp33_ASAP7_75t_L g3187 ( 
.A1(n_1943),
.A2(n_2120),
.B(n_2157),
.C(n_2133),
.Y(n_3187)
);

NAND2x1_ASAP7_75t_L g3188 ( 
.A(n_2228),
.B(n_2089),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2034),
.Y(n_3189)
);

INVx3_ASAP7_75t_L g3190 ( 
.A(n_2204),
.Y(n_3190)
);

O2A1O1Ixp33_ASAP7_75t_L g3191 ( 
.A1(n_1943),
.A2(n_2133),
.B(n_2060),
.C(n_2061),
.Y(n_3191)
);

O2A1O1Ixp33_ASAP7_75t_L g3192 ( 
.A1(n_2050),
.A2(n_2064),
.B(n_2264),
.C(n_2261),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_2753),
.A2(n_2782),
.B(n_2773),
.Y(n_3193)
);

AOI21xp5_ASAP7_75t_L g3194 ( 
.A1(n_2793),
.A2(n_2800),
.B(n_2325),
.Y(n_3194)
);

INVx3_ASAP7_75t_L g3195 ( 
.A(n_2204),
.Y(n_3195)
);

CKINVDCx5p33_ASAP7_75t_R g3196 ( 
.A(n_2582),
.Y(n_3196)
);

NOR2xp33_ASAP7_75t_L g3197 ( 
.A(n_2007),
.B(n_2619),
.Y(n_3197)
);

AND2x4_ASAP7_75t_L g3198 ( 
.A(n_1936),
.B(n_2057),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_2793),
.B(n_2800),
.Y(n_3199)
);

AOI21xp5_ASAP7_75t_L g3200 ( 
.A1(n_2292),
.A2(n_2334),
.B(n_2325),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2334),
.A2(n_2346),
.B(n_2343),
.Y(n_3201)
);

AOI22xp5_ASAP7_75t_L g3202 ( 
.A1(n_2175),
.A2(n_2290),
.B1(n_2564),
.B2(n_1911),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2130),
.B(n_2183),
.Y(n_3203)
);

NAND2xp33_ASAP7_75t_L g3204 ( 
.A(n_2330),
.B(n_2705),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2058),
.Y(n_3205)
);

A2O1A1Ixp33_ASAP7_75t_L g3206 ( 
.A1(n_2290),
.A2(n_2564),
.B(n_2104),
.C(n_2130),
.Y(n_3206)
);

AOI21xp5_ASAP7_75t_L g3207 ( 
.A1(n_2343),
.A2(n_2347),
.B(n_2346),
.Y(n_3207)
);

INVx2_ASAP7_75t_SL g3208 ( 
.A(n_2287),
.Y(n_3208)
);

NOR2xp33_ASAP7_75t_SL g3209 ( 
.A(n_1969),
.B(n_2370),
.Y(n_3209)
);

AOI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_2343),
.A2(n_2347),
.B(n_2346),
.Y(n_3210)
);

AOI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_2347),
.A2(n_2388),
.B(n_2360),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2183),
.B(n_2198),
.Y(n_3212)
);

INVx3_ASAP7_75t_L g3213 ( 
.A(n_2204),
.Y(n_3213)
);

INVxp67_ASAP7_75t_L g3214 ( 
.A(n_2179),
.Y(n_3214)
);

AOI21x1_ASAP7_75t_L g3215 ( 
.A1(n_2360),
.A2(n_2410),
.B(n_2388),
.Y(n_3215)
);

INVx8_ASAP7_75t_L g3216 ( 
.A(n_2184),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2058),
.Y(n_3217)
);

BUFx2_ASAP7_75t_L g3218 ( 
.A(n_2237),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2067),
.Y(n_3219)
);

OR2x6_ASAP7_75t_L g3220 ( 
.A(n_2176),
.B(n_1997),
.Y(n_3220)
);

INVx1_ASAP7_75t_SL g3221 ( 
.A(n_1931),
.Y(n_3221)
);

NOR2xp67_ASAP7_75t_L g3222 ( 
.A(n_2360),
.B(n_2388),
.Y(n_3222)
);

OAI22xp5_ASAP7_75t_L g3223 ( 
.A1(n_1931),
.A2(n_1947),
.B1(n_1951),
.B2(n_1939),
.Y(n_3223)
);

INVx3_ASAP7_75t_L g3224 ( 
.A(n_2204),
.Y(n_3224)
);

AOI21x1_ASAP7_75t_L g3225 ( 
.A1(n_2410),
.A2(n_2440),
.B(n_2429),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2198),
.B(n_2212),
.Y(n_3226)
);

AOI21xp5_ASAP7_75t_L g3227 ( 
.A1(n_2410),
.A2(n_2440),
.B(n_2429),
.Y(n_3227)
);

AOI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_2429),
.A2(n_2446),
.B(n_2440),
.Y(n_3228)
);

OAI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_2125),
.A2(n_2145),
.B(n_2142),
.Y(n_3229)
);

AOI21xp33_ASAP7_75t_L g3230 ( 
.A1(n_2143),
.A2(n_2170),
.B(n_2462),
.Y(n_3230)
);

OAI21xp5_ASAP7_75t_L g3231 ( 
.A1(n_2147),
.A2(n_2165),
.B(n_2164),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_SL g3232 ( 
.A(n_2132),
.B(n_1950),
.Y(n_3232)
);

AOI21xp5_ASAP7_75t_L g3233 ( 
.A1(n_2446),
.A2(n_2473),
.B(n_2455),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_2212),
.B(n_2215),
.Y(n_3234)
);

AOI222xp33_ASAP7_75t_L g3235 ( 
.A1(n_2175),
.A2(n_1911),
.B1(n_2166),
.B2(n_2171),
.C1(n_2151),
.C2(n_1976),
.Y(n_3235)
);

OR2x6_ASAP7_75t_L g3236 ( 
.A(n_2176),
.B(n_1997),
.Y(n_3236)
);

AND2x2_ASAP7_75t_L g3237 ( 
.A(n_2073),
.B(n_2107),
.Y(n_3237)
);

AOI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_2455),
.A2(n_2483),
.B(n_2473),
.Y(n_3238)
);

AOI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_2455),
.A2(n_2483),
.B(n_2473),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_2747),
.B(n_2081),
.Y(n_3240)
);

OAI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_2168),
.A2(n_2107),
.B(n_1947),
.Y(n_3241)
);

AOI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_2488),
.A2(n_2500),
.B(n_2492),
.Y(n_3242)
);

AOI21xp5_ASAP7_75t_L g3243 ( 
.A1(n_2488),
.A2(n_2500),
.B(n_2492),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2215),
.B(n_2073),
.Y(n_3244)
);

AOI21xp5_ASAP7_75t_L g3245 ( 
.A1(n_2488),
.A2(n_2500),
.B(n_2492),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2073),
.B(n_2129),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2129),
.B(n_2160),
.Y(n_3247)
);

CKINVDCx5p33_ASAP7_75t_R g3248 ( 
.A(n_2194),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_2505),
.A2(n_2551),
.B(n_2542),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_2160),
.B(n_1939),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_1951),
.Y(n_3251)
);

OAI22xp5_ASAP7_75t_L g3252 ( 
.A1(n_1953),
.A2(n_1959),
.B1(n_1980),
.B2(n_1972),
.Y(n_3252)
);

NOR2xp33_ASAP7_75t_SL g3253 ( 
.A(n_1969),
.B(n_2370),
.Y(n_3253)
);

O2A1O1Ixp33_ASAP7_75t_L g3254 ( 
.A1(n_2188),
.A2(n_2117),
.B(n_2267),
.C(n_2182),
.Y(n_3254)
);

NOR2xp33_ASAP7_75t_L g3255 ( 
.A(n_2248),
.B(n_2345),
.Y(n_3255)
);

AOI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_2505),
.A2(n_2551),
.B(n_2542),
.Y(n_3256)
);

NOR2xp33_ASAP7_75t_L g3257 ( 
.A(n_2181),
.B(n_2185),
.Y(n_3257)
);

O2A1O1Ixp33_ASAP7_75t_L g3258 ( 
.A1(n_2151),
.A2(n_2166),
.B(n_2171),
.C(n_2239),
.Y(n_3258)
);

OAI22xp5_ASAP7_75t_L g3259 ( 
.A1(n_1953),
.A2(n_1959),
.B1(n_1980),
.B2(n_1972),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_1985),
.B(n_1994),
.Y(n_3260)
);

A2O1A1Ixp33_ASAP7_75t_L g3261 ( 
.A1(n_2213),
.A2(n_2232),
.B(n_2220),
.C(n_2250),
.Y(n_3261)
);

AOI21xp5_ASAP7_75t_L g3262 ( 
.A1(n_2505),
.A2(n_2551),
.B(n_2542),
.Y(n_3262)
);

BUFx4f_ASAP7_75t_L g3263 ( 
.A(n_2285),
.Y(n_3263)
);

AOI21xp5_ASAP7_75t_L g3264 ( 
.A1(n_2576),
.A2(n_2605),
.B(n_2597),
.Y(n_3264)
);

OAI22xp5_ASAP7_75t_L g3265 ( 
.A1(n_1985),
.A2(n_1996),
.B1(n_2002),
.B2(n_1994),
.Y(n_3265)
);

AOI21xp5_ASAP7_75t_L g3266 ( 
.A1(n_2576),
.A2(n_2605),
.B(n_2597),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_1996),
.B(n_2002),
.Y(n_3267)
);

AOI21xp5_ASAP7_75t_L g3268 ( 
.A1(n_2597),
.A2(n_2606),
.B(n_2605),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_2004),
.B(n_2012),
.Y(n_3269)
);

NOR2xp67_ASAP7_75t_L g3270 ( 
.A(n_2606),
.B(n_2607),
.Y(n_3270)
);

A2O1A1Ixp33_ASAP7_75t_L g3271 ( 
.A1(n_2220),
.A2(n_2250),
.B(n_2174),
.C(n_2065),
.Y(n_3271)
);

BUFx3_ASAP7_75t_L g3272 ( 
.A(n_2244),
.Y(n_3272)
);

BUFx3_ASAP7_75t_L g3273 ( 
.A(n_2244),
.Y(n_3273)
);

O2A1O1Ixp33_ASAP7_75t_L g3274 ( 
.A1(n_2240),
.A2(n_2012),
.B(n_2013),
.C(n_2004),
.Y(n_3274)
);

A2O1A1Ixp33_ASAP7_75t_L g3275 ( 
.A1(n_2137),
.A2(n_2163),
.B(n_2066),
.C(n_2013),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_2019),
.Y(n_3276)
);

O2A1O1Ixp33_ASAP7_75t_L g3277 ( 
.A1(n_2019),
.A2(n_2046),
.B(n_2051),
.C(n_2026),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2026),
.B(n_2046),
.Y(n_3278)
);

OAI22xp5_ASAP7_75t_L g3279 ( 
.A1(n_2051),
.A2(n_2062),
.B1(n_2074),
.B2(n_2053),
.Y(n_3279)
);

NAND2xp33_ASAP7_75t_L g3280 ( 
.A(n_1969),
.B(n_2370),
.Y(n_3280)
);

O2A1O1Ixp33_ASAP7_75t_L g3281 ( 
.A1(n_2053),
.A2(n_2074),
.B(n_2087),
.C(n_2062),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_SL g3282 ( 
.A(n_1950),
.B(n_2082),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_SL g3283 ( 
.A(n_1950),
.B(n_2082),
.Y(n_3283)
);

OAI21xp5_ASAP7_75t_L g3284 ( 
.A1(n_2087),
.A2(n_2111),
.B(n_2088),
.Y(n_3284)
);

AOI21xp5_ASAP7_75t_L g3285 ( 
.A1(n_2607),
.A2(n_2627),
.B(n_2626),
.Y(n_3285)
);

AOI21xp5_ASAP7_75t_L g3286 ( 
.A1(n_2607),
.A2(n_2627),
.B(n_2626),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2088),
.Y(n_3287)
);

A2O1A1Ixp33_ASAP7_75t_L g3288 ( 
.A1(n_2137),
.A2(n_2111),
.B(n_2687),
.C(n_2262),
.Y(n_3288)
);

NOR2xp33_ASAP7_75t_L g3289 ( 
.A(n_2233),
.B(n_2238),
.Y(n_3289)
);

AND2x2_ASAP7_75t_L g3290 ( 
.A(n_2208),
.B(n_1936),
.Y(n_3290)
);

AOI21xp5_ASAP7_75t_L g3291 ( 
.A1(n_2626),
.A2(n_2656),
.B(n_2627),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_2216),
.B(n_2218),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_SL g3293 ( 
.A(n_1950),
.B(n_2082),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_2216),
.B(n_2218),
.Y(n_3294)
);

AOI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_2661),
.A2(n_2719),
.B(n_2708),
.Y(n_3295)
);

BUFx4f_ASAP7_75t_L g3296 ( 
.A(n_2285),
.Y(n_3296)
);

OAI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_2262),
.A2(n_2121),
.B(n_2086),
.Y(n_3297)
);

AND2x2_ASAP7_75t_L g3298 ( 
.A(n_2208),
.B(n_1936),
.Y(n_3298)
);

AOI21xp5_ASAP7_75t_L g3299 ( 
.A1(n_2661),
.A2(n_2719),
.B(n_2708),
.Y(n_3299)
);

CKINVDCx5p33_ASAP7_75t_R g3300 ( 
.A(n_2106),
.Y(n_3300)
);

A2O1A1Ixp33_ASAP7_75t_L g3301 ( 
.A1(n_2687),
.A2(n_2202),
.B(n_2210),
.C(n_2141),
.Y(n_3301)
);

AOI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_2708),
.A2(n_2725),
.B(n_2719),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2725),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2725),
.Y(n_3304)
);

O2A1O1Ixp5_ASAP7_75t_L g3305 ( 
.A1(n_2186),
.A2(n_2196),
.B(n_2206),
.C(n_2201),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_2221),
.B(n_2231),
.Y(n_3306)
);

AOI21xp5_ASAP7_75t_L g3307 ( 
.A1(n_2727),
.A2(n_2754),
.B(n_2744),
.Y(n_3307)
);

BUFx12f_ASAP7_75t_L g3308 ( 
.A(n_2336),
.Y(n_3308)
);

AOI21xp5_ASAP7_75t_L g3309 ( 
.A1(n_2727),
.A2(n_2754),
.B(n_2744),
.Y(n_3309)
);

OAI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_2086),
.A2(n_2121),
.B(n_2257),
.Y(n_3310)
);

INVx4_ASAP7_75t_L g3311 ( 
.A(n_1969),
.Y(n_3311)
);

NAND3xp33_ASAP7_75t_L g3312 ( 
.A(n_2257),
.B(n_2233),
.C(n_1963),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_2221),
.B(n_2231),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_2727),
.Y(n_3314)
);

BUFx6f_ASAP7_75t_L g3315 ( 
.A(n_2313),
.Y(n_3315)
);

O2A1O1Ixp5_ASAP7_75t_L g3316 ( 
.A1(n_2209),
.A2(n_2219),
.B(n_2227),
.C(n_2178),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_2236),
.B(n_2251),
.Y(n_3317)
);

AOI22xp5_ASAP7_75t_L g3318 ( 
.A1(n_2118),
.A2(n_2028),
.B1(n_2124),
.B2(n_2247),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_2754),
.A2(n_2760),
.B(n_2759),
.Y(n_3319)
);

BUFx3_ASAP7_75t_L g3320 ( 
.A(n_2244),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_2236),
.B(n_2251),
.Y(n_3321)
);

AOI21xp5_ASAP7_75t_L g3322 ( 
.A1(n_2759),
.A2(n_2761),
.B(n_2760),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_2759),
.A2(n_2761),
.B(n_2760),
.Y(n_3323)
);

AO21x1_ASAP7_75t_L g3324 ( 
.A1(n_2761),
.A2(n_2767),
.B(n_2762),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_2256),
.B(n_2263),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_2256),
.B(n_2263),
.Y(n_3326)
);

AOI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_2762),
.A2(n_2772),
.B(n_2767),
.Y(n_3327)
);

OAI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_2001),
.A2(n_2228),
.B(n_2217),
.Y(n_3328)
);

AOI21xp5_ASAP7_75t_L g3329 ( 
.A1(n_2767),
.A2(n_2772),
.B(n_2228),
.Y(n_3329)
);

AOI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_2118),
.A2(n_2124),
.B1(n_2141),
.B2(n_1944),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2260),
.B(n_2154),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_L g3332 ( 
.A(n_2070),
.B(n_1872),
.Y(n_3332)
);

AND2x4_ASAP7_75t_L g3333 ( 
.A(n_2313),
.B(n_2353),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_2260),
.B(n_2154),
.Y(n_3334)
);

O2A1O1Ixp33_ASAP7_75t_L g3335 ( 
.A1(n_2270),
.A2(n_2169),
.B(n_2197),
.C(n_2193),
.Y(n_3335)
);

OAI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_2001),
.A2(n_2228),
.B(n_2687),
.Y(n_3336)
);

AOI21xp5_ASAP7_75t_L g3337 ( 
.A1(n_2772),
.A2(n_2228),
.B(n_2687),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_2260),
.B(n_2159),
.Y(n_3338)
);

OAI321xp33_ASAP7_75t_L g3339 ( 
.A1(n_1989),
.A2(n_2214),
.A3(n_2192),
.B1(n_2176),
.B2(n_2187),
.C(n_2200),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_2159),
.B(n_2341),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_2159),
.B(n_2341),
.Y(n_3341)
);

OAI21xp5_ASAP7_75t_L g3342 ( 
.A1(n_2270),
.A2(n_1903),
.B(n_2200),
.Y(n_3342)
);

NOR2xp33_ASAP7_75t_SL g3343 ( 
.A(n_1969),
.B(n_2370),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_2237),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_2341),
.B(n_2514),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_SL g3346 ( 
.A(n_1950),
.B(n_2082),
.Y(n_3346)
);

AOI21xp5_ASAP7_75t_L g3347 ( 
.A1(n_2269),
.A2(n_2119),
.B(n_2191),
.Y(n_3347)
);

OAI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_1903),
.A2(n_2103),
.B(n_2095),
.Y(n_3348)
);

BUFx6f_ASAP7_75t_L g3349 ( 
.A(n_2313),
.Y(n_3349)
);

BUFx6f_ASAP7_75t_L g3350 ( 
.A(n_2313),
.Y(n_3350)
);

NOR2xp33_ASAP7_75t_L g3351 ( 
.A(n_2070),
.B(n_1872),
.Y(n_3351)
);

AND2x2_ASAP7_75t_L g3352 ( 
.A(n_2191),
.B(n_2092),
.Y(n_3352)
);

AOI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_2269),
.A2(n_2119),
.B(n_2191),
.Y(n_3353)
);

AOI21xp5_ASAP7_75t_L g3354 ( 
.A1(n_2269),
.A2(n_2119),
.B(n_2191),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_2341),
.B(n_2514),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_SL g3356 ( 
.A(n_2082),
.B(n_2113),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_2341),
.B(n_2514),
.Y(n_3357)
);

NAND2xp33_ASAP7_75t_L g3358 ( 
.A(n_1969),
.B(n_2370),
.Y(n_3358)
);

BUFx3_ASAP7_75t_L g3359 ( 
.A(n_2341),
.Y(n_3359)
);

AND2x6_ASAP7_75t_L g3360 ( 
.A(n_2014),
.B(n_2030),
.Y(n_3360)
);

OAI321xp33_ASAP7_75t_L g3361 ( 
.A1(n_2192),
.A2(n_2176),
.A3(n_2672),
.B1(n_2434),
.B2(n_2285),
.C(n_2804),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_2341),
.B(n_2514),
.Y(n_3362)
);

OR2x2_ASAP7_75t_SL g3363 ( 
.A(n_2173),
.B(n_2353),
.Y(n_3363)
);

AOI21xp5_ASAP7_75t_L g3364 ( 
.A1(n_2269),
.A2(n_2119),
.B(n_2353),
.Y(n_3364)
);

O2A1O1Ixp5_ASAP7_75t_L g3365 ( 
.A1(n_2116),
.A2(n_2156),
.B(n_2134),
.C(n_2148),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_2092),
.B(n_2139),
.Y(n_3366)
);

BUFx6f_ASAP7_75t_L g3367 ( 
.A(n_2353),
.Y(n_3367)
);

HB1xp67_ASAP7_75t_L g3368 ( 
.A(n_2241),
.Y(n_3368)
);

OAI22xp5_ASAP7_75t_L g3369 ( 
.A1(n_2184),
.A2(n_2561),
.B1(n_2553),
.B2(n_2664),
.Y(n_3369)
);

OAI22xp5_ASAP7_75t_L g3370 ( 
.A1(n_2184),
.A2(n_2462),
.B1(n_2553),
.B2(n_2561),
.Y(n_3370)
);

AND2x4_ASAP7_75t_L g3371 ( 
.A(n_2353),
.B(n_2474),
.Y(n_3371)
);

INVx2_ASAP7_75t_SL g3372 ( 
.A(n_2353),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_2092),
.B(n_2139),
.Y(n_3373)
);

AOI21xp5_ASAP7_75t_L g3374 ( 
.A1(n_2269),
.A2(n_2558),
.B(n_2789),
.Y(n_3374)
);

NOR2xp33_ASAP7_75t_L g3375 ( 
.A(n_1884),
.B(n_1887),
.Y(n_3375)
);

OAI21xp5_ASAP7_75t_L g3376 ( 
.A1(n_2144),
.A2(n_2162),
.B(n_2158),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_2092),
.B(n_2139),
.Y(n_3377)
);

HB1xp67_ASAP7_75t_L g3378 ( 
.A(n_2241),
.Y(n_3378)
);

CKINVDCx20_ASAP7_75t_R g3379 ( 
.A(n_1929),
.Y(n_3379)
);

BUFx3_ASAP7_75t_L g3380 ( 
.A(n_2514),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_2514),
.B(n_2139),
.Y(n_3381)
);

BUFx12f_ASAP7_75t_L g3382 ( 
.A(n_2336),
.Y(n_3382)
);

AOI21xp5_ASAP7_75t_L g3383 ( 
.A1(n_2474),
.A2(n_2688),
.B(n_2789),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_2514),
.B(n_2152),
.Y(n_3384)
);

INVx3_ASAP7_75t_L g3385 ( 
.A(n_2246),
.Y(n_3385)
);

AOI21xp5_ASAP7_75t_L g3386 ( 
.A1(n_2474),
.A2(n_2688),
.B(n_2789),
.Y(n_3386)
);

AND2x2_ASAP7_75t_L g3387 ( 
.A(n_2152),
.B(n_2167),
.Y(n_3387)
);

NOR2xp33_ASAP7_75t_L g3388 ( 
.A(n_1884),
.B(n_1887),
.Y(n_3388)
);

AOI22xp5_ASAP7_75t_L g3389 ( 
.A1(n_1969),
.A2(n_2370),
.B1(n_2771),
.B2(n_2184),
.Y(n_3389)
);

INVx2_ASAP7_75t_SL g3390 ( 
.A(n_2474),
.Y(n_3390)
);

O2A1O1Ixp33_ASAP7_75t_L g3391 ( 
.A1(n_2169),
.A2(n_2211),
.B(n_2664),
.C(n_2161),
.Y(n_3391)
);

BUFx3_ASAP7_75t_L g3392 ( 
.A(n_2014),
.Y(n_3392)
);

NOR2xp33_ASAP7_75t_L g3393 ( 
.A(n_1901),
.B(n_1930),
.Y(n_3393)
);

AOI21xp33_ASAP7_75t_L g3394 ( 
.A1(n_2176),
.A2(n_2105),
.B(n_2022),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_2152),
.B(n_2167),
.Y(n_3395)
);

INVx4_ASAP7_75t_L g3396 ( 
.A(n_1969),
.Y(n_3396)
);

AOI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_2474),
.A2(n_2789),
.B(n_2721),
.Y(n_3397)
);

BUFx6f_ASAP7_75t_L g3398 ( 
.A(n_2474),
.Y(n_3398)
);

AOI21xp5_ASAP7_75t_L g3399 ( 
.A1(n_2555),
.A2(n_2789),
.B(n_2721),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_2152),
.B(n_2167),
.Y(n_3400)
);

AOI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_2555),
.A2(n_2789),
.B(n_2721),
.Y(n_3401)
);

BUFx3_ASAP7_75t_L g3402 ( 
.A(n_2014),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_2555),
.A2(n_2558),
.B(n_2721),
.Y(n_3403)
);

AOI21xp5_ASAP7_75t_L g3404 ( 
.A1(n_2555),
.A2(n_2558),
.B(n_2721),
.Y(n_3404)
);

O2A1O1Ixp33_ASAP7_75t_L g3405 ( 
.A1(n_1901),
.A2(n_2295),
.B(n_1930),
.C(n_2783),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_2167),
.B(n_2222),
.Y(n_3406)
);

AOI21xp5_ASAP7_75t_L g3407 ( 
.A1(n_2555),
.A2(n_2721),
.B(n_2688),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_2222),
.B(n_2226),
.Y(n_3408)
);

AND3x1_ASAP7_75t_L g3409 ( 
.A(n_1993),
.B(n_2487),
.C(n_2783),
.Y(n_3409)
);

OAI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_2229),
.A2(n_2207),
.B(n_2205),
.Y(n_3410)
);

AOI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_2555),
.A2(n_2688),
.B(n_2558),
.Y(n_3411)
);

INVx3_ASAP7_75t_L g3412 ( 
.A(n_2370),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_SL g3413 ( 
.A(n_2082),
.B(n_2113),
.Y(n_3413)
);

A2O1A1Ixp33_ASAP7_75t_L g3414 ( 
.A1(n_2229),
.A2(n_2153),
.B(n_2288),
.C(n_2296),
.Y(n_3414)
);

OR2x6_ASAP7_75t_L g3415 ( 
.A(n_1999),
.B(n_2022),
.Y(n_3415)
);

AOI21xp5_ASAP7_75t_L g3416 ( 
.A1(n_2558),
.A2(n_2688),
.B(n_1973),
.Y(n_3416)
);

NOR2xp67_ASAP7_75t_L g3417 ( 
.A(n_1973),
.B(n_1982),
.Y(n_3417)
);

OAI21xp33_ASAP7_75t_L g3418 ( 
.A1(n_2241),
.A2(n_2804),
.B(n_2434),
.Y(n_3418)
);

AOI21x1_ASAP7_75t_L g3419 ( 
.A1(n_2229),
.A2(n_2226),
.B(n_2265),
.Y(n_3419)
);

AOI21xp5_ASAP7_75t_L g3420 ( 
.A1(n_2558),
.A2(n_2688),
.B(n_1973),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_2226),
.B(n_2199),
.Y(n_3421)
);

AOI21xp5_ASAP7_75t_L g3422 ( 
.A1(n_1973),
.A2(n_1982),
.B(n_2672),
.Y(n_3422)
);

NOR3xp33_ASAP7_75t_L g3423 ( 
.A(n_1999),
.B(n_2096),
.C(n_2105),
.Y(n_3423)
);

BUFx6f_ASAP7_75t_L g3424 ( 
.A(n_2113),
.Y(n_3424)
);

NOR2xp67_ASAP7_75t_L g3425 ( 
.A(n_1982),
.B(n_2273),
.Y(n_3425)
);

O2A1O1Ixp33_ASAP7_75t_L g3426 ( 
.A1(n_1993),
.A2(n_2321),
.B(n_2715),
.C(n_2702),
.Y(n_3426)
);

OAI21xp5_ASAP7_75t_L g3427 ( 
.A1(n_2229),
.A2(n_2804),
.B(n_2434),
.Y(n_3427)
);

AOI21xp5_ASAP7_75t_L g3428 ( 
.A1(n_1982),
.A2(n_2672),
.B(n_2153),
.Y(n_3428)
);

AOI21xp5_ASAP7_75t_L g3429 ( 
.A1(n_2273),
.A2(n_2296),
.B(n_2522),
.Y(n_3429)
);

AOI21xp5_ASAP7_75t_L g3430 ( 
.A1(n_2273),
.A2(n_2296),
.B(n_2522),
.Y(n_3430)
);

BUFx6f_ASAP7_75t_SL g3431 ( 
.A(n_1929),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_L g3432 ( 
.A(n_2295),
.B(n_2300),
.Y(n_3432)
);

A2O1A1Ixp33_ASAP7_75t_L g3433 ( 
.A1(n_2273),
.A2(n_2288),
.B(n_2296),
.C(n_2709),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_L g3434 ( 
.A(n_2300),
.B(n_2321),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_2265),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_2224),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_2199),
.B(n_2224),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_2288),
.A2(n_2646),
.B(n_2682),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_2245),
.B(n_2259),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_2245),
.B(n_2259),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_2288),
.B(n_2421),
.Y(n_3441)
);

BUFx6f_ASAP7_75t_L g3442 ( 
.A(n_2113),
.Y(n_3442)
);

OAI22xp5_ASAP7_75t_L g3443 ( 
.A1(n_2030),
.A2(n_2071),
.B1(n_2096),
.B2(n_2041),
.Y(n_3443)
);

AOI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_2421),
.A2(n_2709),
.B(n_2682),
.Y(n_3444)
);

AOI21xp5_ASAP7_75t_L g3445 ( 
.A1(n_2421),
.A2(n_2709),
.B(n_2682),
.Y(n_3445)
);

A2O1A1Ixp33_ASAP7_75t_L g3446 ( 
.A1(n_2421),
.A2(n_2682),
.B(n_2522),
.C(n_2709),
.Y(n_3446)
);

AND2x2_ASAP7_75t_L g3447 ( 
.A(n_2172),
.B(n_2646),
.Y(n_3447)
);

INVx3_ASAP7_75t_L g3448 ( 
.A(n_2370),
.Y(n_3448)
);

A2O1A1Ixp33_ASAP7_75t_L g3449 ( 
.A1(n_2522),
.A2(n_2646),
.B(n_2348),
.C(n_2041),
.Y(n_3449)
);

OAI22xp5_ASAP7_75t_L g3450 ( 
.A1(n_2030),
.A2(n_2071),
.B1(n_1955),
.B2(n_1975),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_2646),
.B(n_2071),
.Y(n_3451)
);

OAI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_2047),
.A2(n_2150),
.B(n_2149),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_2172),
.B(n_2771),
.Y(n_3453)
);

AND2x4_ASAP7_75t_L g3454 ( 
.A(n_2348),
.B(n_2172),
.Y(n_3454)
);

AOI21x1_ASAP7_75t_L g3455 ( 
.A1(n_2223),
.A2(n_2266),
.B(n_2258),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_2172),
.B(n_2771),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_SL g3457 ( 
.A(n_2113),
.B(n_2146),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_SL g3458 ( 
.A(n_2113),
.B(n_2146),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_2235),
.Y(n_3459)
);

BUFx6f_ASAP7_75t_L g3460 ( 
.A(n_2146),
.Y(n_3460)
);

AO22x1_ASAP7_75t_L g3461 ( 
.A1(n_1929),
.A2(n_1955),
.B1(n_1975),
.B2(n_2781),
.Y(n_3461)
);

NOR2xp33_ASAP7_75t_L g3462 ( 
.A(n_2364),
.B(n_2589),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_2771),
.B(n_2146),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_SL g3464 ( 
.A(n_2146),
.B(n_2771),
.Y(n_3464)
);

AOI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_2146),
.A2(n_2348),
.B(n_2771),
.Y(n_3465)
);

BUFx6f_ASAP7_75t_L g3466 ( 
.A(n_1955),
.Y(n_3466)
);

AOI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_2771),
.A2(n_2140),
.B(n_2098),
.Y(n_3467)
);

O2A1O1Ixp33_ASAP7_75t_L g3468 ( 
.A1(n_2364),
.A2(n_2715),
.B(n_2702),
.C(n_2487),
.Y(n_3468)
);

BUFx4f_ASAP7_75t_L g3469 ( 
.A(n_2373),
.Y(n_3469)
);

O2A1O1Ixp33_ASAP7_75t_L g3470 ( 
.A1(n_2373),
.A2(n_2671),
.B(n_2642),
.C(n_2424),
.Y(n_3470)
);

AND2x4_ASAP7_75t_L g3471 ( 
.A(n_1975),
.B(n_2795),
.Y(n_3471)
);

OAI22xp5_ASAP7_75t_L g3472 ( 
.A1(n_2315),
.A2(n_2528),
.B1(n_2781),
.B2(n_2700),
.Y(n_3472)
);

A2O1A1Ixp33_ASAP7_75t_L g3473 ( 
.A1(n_2377),
.A2(n_2523),
.B(n_2671),
.C(n_2642),
.Y(n_3473)
);

OAI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_2100),
.A2(n_2108),
.B(n_2114),
.Y(n_3474)
);

OAI21xp33_ASAP7_75t_L g3475 ( 
.A1(n_2315),
.A2(n_2528),
.B(n_2781),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_2771),
.B(n_2230),
.Y(n_3476)
);

AOI21xp5_ASAP7_75t_L g3477 ( 
.A1(n_2771),
.A2(n_2523),
.B(n_2563),
.Y(n_3477)
);

AOI21xp5_ASAP7_75t_L g3478 ( 
.A1(n_2377),
.A2(n_2634),
.B(n_2563),
.Y(n_3478)
);

NOR2xp33_ASAP7_75t_L g3479 ( 
.A(n_2415),
.B(n_2424),
.Y(n_3479)
);

AO21x1_ASAP7_75t_L g3480 ( 
.A1(n_2471),
.A2(n_2701),
.B(n_2673),
.Y(n_3480)
);

CKINVDCx10_ASAP7_75t_R g3481 ( 
.A(n_2106),
.Y(n_3481)
);

NOR2xp33_ASAP7_75t_L g3482 ( 
.A(n_2415),
.B(n_2589),
.Y(n_3482)
);

A2O1A1Ixp33_ASAP7_75t_L g3483 ( 
.A1(n_2422),
.A2(n_2634),
.B(n_2601),
.C(n_2623),
.Y(n_3483)
);

AOI22xp33_ASAP7_75t_L g3484 ( 
.A1(n_2177),
.A2(n_2315),
.B1(n_2355),
.B2(n_2700),
.Y(n_3484)
);

AOI21xp5_ASAP7_75t_L g3485 ( 
.A1(n_2422),
.A2(n_2623),
.B(n_2601),
.Y(n_3485)
);

AOI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_2355),
.A2(n_2428),
.B(n_2700),
.Y(n_3486)
);

AND2x2_ASAP7_75t_L g3487 ( 
.A(n_2355),
.B(n_2428),
.Y(n_3487)
);

NOR3xp33_ASAP7_75t_L g3488 ( 
.A(n_2428),
.B(n_2795),
.C(n_2580),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_2520),
.B(n_2795),
.Y(n_3489)
);

AOI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_2520),
.A2(n_2580),
.B(n_2528),
.Y(n_3490)
);

AOI21xp5_ASAP7_75t_L g3491 ( 
.A1(n_2520),
.A2(n_2580),
.B(n_2497),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_SL g3492 ( 
.A(n_2471),
.B(n_2497),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_2511),
.B(n_2673),
.Y(n_3493)
);

OR2x2_ASAP7_75t_L g3494 ( 
.A(n_2511),
.B(n_2701),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_2562),
.B(n_2045),
.Y(n_3495)
);

AOI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3496)
);

OAI21xp5_ASAP7_75t_L g3497 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_SL g3498 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3498)
);

OAI22xp5_ASAP7_75t_L g3499 ( 
.A1(n_1859),
.A2(n_2317),
.B1(n_2318),
.B2(n_2279),
.Y(n_3499)
);

AOI21xp5_ASAP7_75t_L g3500 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3500)
);

AOI22xp5_ASAP7_75t_L g3501 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3501)
);

AOI21xp5_ASAP7_75t_L g3502 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3502)
);

NOR2x1_ASAP7_75t_L g3503 ( 
.A(n_2389),
.B(n_2408),
.Y(n_3503)
);

CKINVDCx20_ASAP7_75t_R g3504 ( 
.A(n_1905),
.Y(n_3504)
);

A2O1A1Ixp33_ASAP7_75t_L g3505 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3506)
);

AOI21xp5_ASAP7_75t_L g3507 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3508)
);

OR2x6_ASAP7_75t_L g3509 ( 
.A(n_2387),
.B(n_2433),
.Y(n_3509)
);

A2O1A1Ixp33_ASAP7_75t_L g3510 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3510)
);

OAI21xp5_ASAP7_75t_L g3511 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3515)
);

INVx2_ASAP7_75t_SL g3516 ( 
.A(n_2180),
.Y(n_3516)
);

AND2x4_ASAP7_75t_L g3517 ( 
.A(n_2362),
.B(n_2386),
.Y(n_3517)
);

AND2x4_ASAP7_75t_L g3518 ( 
.A(n_2362),
.B(n_2386),
.Y(n_3518)
);

O2A1O1Ixp33_ASAP7_75t_L g3519 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_SL g3520 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3520)
);

AOI21xp5_ASAP7_75t_L g3521 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3521)
);

AOI22xp5_ASAP7_75t_L g3522 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3523)
);

NOR2xp33_ASAP7_75t_L g3524 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3525)
);

INVx4_ASAP7_75t_SL g3526 ( 
.A(n_2387),
.Y(n_3526)
);

AOI21xp5_ASAP7_75t_L g3527 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3527)
);

INVx3_ASAP7_75t_L g3528 ( 
.A(n_2554),
.Y(n_3528)
);

AOI22xp5_ASAP7_75t_L g3529 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_SL g3530 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3531)
);

OAI22xp5_ASAP7_75t_L g3532 ( 
.A1(n_1859),
.A2(n_2317),
.B1(n_2318),
.B2(n_2279),
.Y(n_3532)
);

NAND3xp33_ASAP7_75t_SL g3533 ( 
.A(n_1859),
.B(n_2317),
.C(n_2279),
.Y(n_3533)
);

O2A1O1Ixp33_ASAP7_75t_L g3534 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3535)
);

AO21x1_ASAP7_75t_L g3536 ( 
.A1(n_1882),
.A2(n_2357),
.B(n_2284),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_SL g3537 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3537)
);

AOI21xp5_ASAP7_75t_L g3538 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3538)
);

AOI21xp5_ASAP7_75t_L g3539 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3540)
);

AOI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3541)
);

AOI21xp5_ASAP7_75t_L g3542 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3542)
);

AOI21xp5_ASAP7_75t_L g3543 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3543)
);

A2O1A1Ixp33_ASAP7_75t_L g3544 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3545)
);

CKINVDCx10_ASAP7_75t_R g3546 ( 
.A(n_2184),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3547)
);

AOI21xp5_ASAP7_75t_L g3548 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3548)
);

A2O1A1Ixp33_ASAP7_75t_L g3549 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3549)
);

HB1xp67_ASAP7_75t_L g3550 ( 
.A(n_2309),
.Y(n_3550)
);

AOI21xp5_ASAP7_75t_L g3551 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3552)
);

OAI21xp5_ASAP7_75t_L g3553 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3554)
);

AOI22xp5_ASAP7_75t_L g3555 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3556)
);

AOI21xp5_ASAP7_75t_L g3557 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3557)
);

NAND2xp33_ASAP7_75t_L g3558 ( 
.A(n_2489),
.B(n_1603),
.Y(n_3558)
);

AND2x4_ASAP7_75t_L g3559 ( 
.A(n_2362),
.B(n_2386),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3560)
);

AOI21xp5_ASAP7_75t_L g3561 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_L g3562 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3562)
);

OAI22xp5_ASAP7_75t_L g3563 ( 
.A1(n_1859),
.A2(n_2317),
.B1(n_2318),
.B2(n_2279),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_L g3565 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_SL g3568 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3568)
);

AOI21xp33_ASAP7_75t_L g3569 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3569)
);

NOR2xp33_ASAP7_75t_L g3570 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3571)
);

AOI21xp5_ASAP7_75t_L g3572 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3572)
);

AOI21xp5_ASAP7_75t_L g3573 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3573)
);

AOI21xp5_ASAP7_75t_L g3574 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3574)
);

OAI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3575)
);

INVx4_ASAP7_75t_L g3576 ( 
.A(n_1914),
.Y(n_3576)
);

AND2x2_ASAP7_75t_L g3577 ( 
.A(n_1878),
.B(n_1897),
.Y(n_3577)
);

NOR2xp33_ASAP7_75t_L g3578 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3578)
);

AOI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3579)
);

OAI21xp33_ASAP7_75t_L g3580 ( 
.A1(n_1859),
.A2(n_2317),
.B(n_2279),
.Y(n_3580)
);

O2A1O1Ixp33_ASAP7_75t_L g3581 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_SL g3582 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3582)
);

AOI21xp5_ASAP7_75t_L g3583 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3583)
);

NAND2x1p5_ASAP7_75t_L g3584 ( 
.A(n_1914),
.B(n_2617),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3585)
);

AOI21xp5_ASAP7_75t_L g3586 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3586)
);

AOI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_1878),
.B(n_1897),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3590)
);

INVx4_ASAP7_75t_L g3591 ( 
.A(n_1914),
.Y(n_3591)
);

OAI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3593)
);

BUFx4f_ASAP7_75t_L g3594 ( 
.A(n_1986),
.Y(n_3594)
);

AND2x4_ASAP7_75t_L g3595 ( 
.A(n_2362),
.B(n_2386),
.Y(n_3595)
);

O2A1O1Ixp33_ASAP7_75t_L g3596 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3596)
);

A2O1A1Ixp33_ASAP7_75t_L g3597 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3597)
);

INVx1_ASAP7_75t_SL g3598 ( 
.A(n_1893),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3599)
);

NOR2xp33_ASAP7_75t_L g3600 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3600)
);

AO21x1_ASAP7_75t_L g3601 ( 
.A1(n_1882),
.A2(n_2357),
.B(n_2284),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_2797),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_SL g3604 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3604)
);

OAI21xp33_ASAP7_75t_L g3605 ( 
.A1(n_1859),
.A2(n_2317),
.B(n_2279),
.Y(n_3605)
);

INVx11_ASAP7_75t_L g3606 ( 
.A(n_1976),
.Y(n_3606)
);

AOI21xp5_ASAP7_75t_L g3607 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3607)
);

A2O1A1Ixp33_ASAP7_75t_L g3608 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3608)
);

NOR2xp33_ASAP7_75t_L g3609 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3609)
);

OAI21xp5_ASAP7_75t_L g3610 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_2136),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_SL g3612 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3612)
);

O2A1O1Ixp33_ASAP7_75t_L g3613 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_2797),
.Y(n_3614)
);

NOR2xp33_ASAP7_75t_L g3615 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3615)
);

AOI22xp33_ASAP7_75t_L g3616 ( 
.A1(n_2294),
.A2(n_1311),
.B1(n_2305),
.B2(n_2297),
.Y(n_3616)
);

AOI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3617)
);

O2A1O1Ixp33_ASAP7_75t_L g3618 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_2797),
.Y(n_3619)
);

AOI21xp5_ASAP7_75t_L g3620 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3620)
);

OAI21xp5_ASAP7_75t_L g3621 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3621)
);

AOI21xp5_ASAP7_75t_L g3622 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3623)
);

OR2x6_ASAP7_75t_L g3624 ( 
.A(n_2387),
.B(n_2433),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_2797),
.Y(n_3625)
);

AND2x6_ASAP7_75t_SL g3626 ( 
.A(n_1898),
.B(n_1896),
.Y(n_3626)
);

OAI21xp33_ASAP7_75t_L g3627 ( 
.A1(n_1859),
.A2(n_2317),
.B(n_2279),
.Y(n_3627)
);

A2O1A1Ixp33_ASAP7_75t_L g3628 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3628)
);

AOI21xp5_ASAP7_75t_L g3629 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3629)
);

AOI22xp5_ASAP7_75t_L g3630 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3630)
);

AOI21xp5_ASAP7_75t_L g3631 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3631)
);

AOI21xp5_ASAP7_75t_L g3632 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3632)
);

NOR2xp33_ASAP7_75t_L g3633 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_1878),
.B(n_1897),
.Y(n_3634)
);

AOI21xp5_ASAP7_75t_L g3635 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3635)
);

AOI21xp5_ASAP7_75t_L g3636 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3637)
);

AOI21xp5_ASAP7_75t_L g3638 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3638)
);

A2O1A1Ixp33_ASAP7_75t_L g3639 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3639)
);

AOI21xp5_ASAP7_75t_L g3640 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_2797),
.Y(n_3641)
);

NAND2xp33_ASAP7_75t_L g3642 ( 
.A(n_2489),
.B(n_1603),
.Y(n_3642)
);

AOI22xp5_ASAP7_75t_L g3643 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3643)
);

AOI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_SL g3647 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3647)
);

AOI22xp5_ASAP7_75t_L g3648 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3649)
);

NAND2xp33_ASAP7_75t_L g3650 ( 
.A(n_2489),
.B(n_1603),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3651)
);

NOR2xp33_ASAP7_75t_L g3652 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3652)
);

O2A1O1Ixp33_ASAP7_75t_L g3653 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3653)
);

AOI21xp5_ASAP7_75t_L g3654 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3654)
);

AOI21xp5_ASAP7_75t_L g3655 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3655)
);

AOI21xp5_ASAP7_75t_L g3656 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3657)
);

AOI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3658)
);

AOI21xp5_ASAP7_75t_L g3659 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3659)
);

BUFx6f_ASAP7_75t_L g3660 ( 
.A(n_1914),
.Y(n_3660)
);

INVx2_ASAP7_75t_SL g3661 ( 
.A(n_2180),
.Y(n_3661)
);

BUFx6f_ASAP7_75t_L g3662 ( 
.A(n_1914),
.Y(n_3662)
);

NOR2xp33_ASAP7_75t_L g3663 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3663)
);

AOI21xp5_ASAP7_75t_L g3664 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3664)
);

O2A1O1Ixp33_ASAP7_75t_L g3665 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3666)
);

NOR2xp33_ASAP7_75t_L g3667 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3668)
);

HB1xp67_ASAP7_75t_L g3669 ( 
.A(n_2309),
.Y(n_3669)
);

NOR2x1_ASAP7_75t_L g3670 ( 
.A(n_2389),
.B(n_2408),
.Y(n_3670)
);

AOI21xp5_ASAP7_75t_L g3671 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3671)
);

NAND3xp33_ASAP7_75t_L g3672 ( 
.A(n_1882),
.B(n_2357),
.C(n_2284),
.Y(n_3672)
);

AOI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3673)
);

NOR2xp33_ASAP7_75t_L g3674 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3674)
);

OAI321xp33_ASAP7_75t_L g3675 ( 
.A1(n_1882),
.A2(n_2284),
.A3(n_2359),
.B1(n_2635),
.B2(n_2538),
.C(n_2357),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3676)
);

O2A1O1Ixp5_ASAP7_75t_L g3677 ( 
.A1(n_1882),
.A2(n_1220),
.B(n_2357),
.C(n_2284),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_2797),
.Y(n_3679)
);

AOI21xp5_ASAP7_75t_L g3680 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3680)
);

O2A1O1Ixp33_ASAP7_75t_L g3681 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3681)
);

O2A1O1Ixp33_ASAP7_75t_SL g3682 ( 
.A1(n_1898),
.A2(n_1220),
.B(n_2299),
.C(n_2282),
.Y(n_3682)
);

A2O1A1Ixp33_ASAP7_75t_L g3683 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3684)
);

A2O1A1Ixp33_ASAP7_75t_L g3685 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3685)
);

A2O1A1Ixp33_ASAP7_75t_L g3686 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3686)
);

CKINVDCx5p33_ASAP7_75t_R g3687 ( 
.A(n_1905),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_SL g3688 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3688)
);

OAI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3689)
);

AOI21xp5_ASAP7_75t_L g3690 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3690)
);

INVx3_ASAP7_75t_L g3691 ( 
.A(n_2554),
.Y(n_3691)
);

CKINVDCx5p33_ASAP7_75t_R g3692 ( 
.A(n_1905),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3693)
);

INVx3_ASAP7_75t_L g3694 ( 
.A(n_2554),
.Y(n_3694)
);

OAI22xp5_ASAP7_75t_L g3695 ( 
.A1(n_1859),
.A2(n_2317),
.B1(n_2318),
.B2(n_2279),
.Y(n_3695)
);

O2A1O1Ixp33_ASAP7_75t_SL g3696 ( 
.A1(n_1898),
.A2(n_1220),
.B(n_2299),
.C(n_2282),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3697)
);

A2O1A1Ixp33_ASAP7_75t_L g3698 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3698)
);

OAI21xp33_ASAP7_75t_L g3699 ( 
.A1(n_1859),
.A2(n_2317),
.B(n_2279),
.Y(n_3699)
);

CKINVDCx20_ASAP7_75t_R g3700 ( 
.A(n_1905),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3701)
);

NOR2xp33_ASAP7_75t_L g3702 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3702)
);

BUFx3_ASAP7_75t_L g3703 ( 
.A(n_2244),
.Y(n_3703)
);

O2A1O1Ixp33_ASAP7_75t_L g3704 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3704)
);

BUFx3_ASAP7_75t_L g3705 ( 
.A(n_2244),
.Y(n_3705)
);

NOR2xp33_ASAP7_75t_L g3706 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3706)
);

O2A1O1Ixp33_ASAP7_75t_L g3707 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_2797),
.Y(n_3709)
);

AOI22xp5_ASAP7_75t_L g3710 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3710)
);

AOI21xp5_ASAP7_75t_L g3711 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3711)
);

OAI21xp5_ASAP7_75t_L g3712 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3712)
);

INVx1_ASAP7_75t_SL g3713 ( 
.A(n_1893),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_2797),
.Y(n_3714)
);

OAI22xp5_ASAP7_75t_L g3715 ( 
.A1(n_1859),
.A2(n_2317),
.B1(n_2318),
.B2(n_2279),
.Y(n_3715)
);

AOI21xp5_ASAP7_75t_L g3716 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3716)
);

AOI22xp5_ASAP7_75t_L g3717 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3718)
);

AOI21xp5_ASAP7_75t_L g3719 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3720)
);

INVx2_ASAP7_75t_SL g3721 ( 
.A(n_2180),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3722)
);

AOI21xp5_ASAP7_75t_L g3723 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3723)
);

AOI21xp5_ASAP7_75t_L g3724 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3724)
);

AO21x1_ASAP7_75t_L g3725 ( 
.A1(n_1882),
.A2(n_2357),
.B(n_2284),
.Y(n_3725)
);

AOI21xp5_ASAP7_75t_L g3726 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3726)
);

AOI21xp5_ASAP7_75t_L g3727 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3727)
);

A2O1A1Ixp33_ASAP7_75t_L g3728 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3730)
);

AOI21xp5_ASAP7_75t_L g3731 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3731)
);

OAI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_1859),
.A2(n_2317),
.B1(n_2318),
.B2(n_2279),
.Y(n_3732)
);

AOI21xp5_ASAP7_75t_L g3733 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3733)
);

CKINVDCx5p33_ASAP7_75t_R g3734 ( 
.A(n_1905),
.Y(n_3734)
);

NOR2xp67_ASAP7_75t_L g3735 ( 
.A(n_2284),
.B(n_1273),
.Y(n_3735)
);

AOI21xp5_ASAP7_75t_L g3736 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3736)
);

A2O1A1Ixp33_ASAP7_75t_L g3737 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3737)
);

O2A1O1Ixp33_ASAP7_75t_SL g3738 ( 
.A1(n_1898),
.A2(n_1220),
.B(n_2299),
.C(n_2282),
.Y(n_3738)
);

NOR2xp33_ASAP7_75t_L g3739 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3739)
);

NOR2xp33_ASAP7_75t_L g3740 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3740)
);

AND2x2_ASAP7_75t_L g3741 ( 
.A(n_1878),
.B(n_1897),
.Y(n_3741)
);

AOI21xp33_ASAP7_75t_L g3742 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_2797),
.Y(n_3743)
);

AOI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3744)
);

AND2x2_ASAP7_75t_L g3745 ( 
.A(n_1878),
.B(n_1897),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3746)
);

BUFx3_ASAP7_75t_L g3747 ( 
.A(n_2244),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_SL g3748 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3748)
);

A2O1A1Ixp33_ASAP7_75t_L g3749 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_2797),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3751)
);

A2O1A1Ixp33_ASAP7_75t_L g3752 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3752)
);

NOR2x1_ASAP7_75t_L g3753 ( 
.A(n_2389),
.B(n_2408),
.Y(n_3753)
);

AOI21xp5_ASAP7_75t_L g3754 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3756)
);

O2A1O1Ixp33_ASAP7_75t_L g3757 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3757)
);

NOR2xp33_ASAP7_75t_SL g3758 ( 
.A(n_1920),
.B(n_1914),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_SL g3760 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3760)
);

NOR2xp33_ASAP7_75t_L g3761 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_1878),
.B(n_1897),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3764)
);

AOI22xp5_ASAP7_75t_L g3765 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3765)
);

AOI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3766)
);

NOR2xp33_ASAP7_75t_L g3767 ( 
.A(n_1896),
.B(n_1886),
.Y(n_3767)
);

CKINVDCx10_ASAP7_75t_R g3768 ( 
.A(n_2184),
.Y(n_3768)
);

AOI21xp5_ASAP7_75t_L g3769 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3769)
);

AOI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_1878),
.B(n_1897),
.Y(n_3771)
);

BUFx2_ASAP7_75t_L g3772 ( 
.A(n_2387),
.Y(n_3772)
);

OAI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3774)
);

AND2x2_ASAP7_75t_L g3775 ( 
.A(n_1878),
.B(n_1897),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_SL g3776 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3776)
);

NOR2xp33_ASAP7_75t_SL g3777 ( 
.A(n_1920),
.B(n_1914),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3778)
);

BUFx6f_ASAP7_75t_L g3779 ( 
.A(n_1914),
.Y(n_3779)
);

INVx6_ASAP7_75t_L g3780 ( 
.A(n_2374),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3781)
);

AOI21x1_ASAP7_75t_L g3782 ( 
.A1(n_2254),
.A2(n_2585),
.B(n_2304),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3783)
);

INVx1_ASAP7_75t_SL g3784 ( 
.A(n_1893),
.Y(n_3784)
);

AOI21xp5_ASAP7_75t_L g3785 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3785)
);

AOI21xp5_ASAP7_75t_L g3786 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3786)
);

O2A1O1Ixp33_ASAP7_75t_SL g3787 ( 
.A1(n_1898),
.A2(n_1220),
.B(n_2299),
.C(n_2282),
.Y(n_3787)
);

OAI221xp5_ASAP7_75t_L g3788 ( 
.A1(n_1859),
.A2(n_2279),
.B1(n_2344),
.B2(n_2318),
.C(n_2317),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_2797),
.Y(n_3790)
);

INVx4_ASAP7_75t_L g3791 ( 
.A(n_1914),
.Y(n_3791)
);

AND3x2_ASAP7_75t_L g3792 ( 
.A(n_2118),
.B(n_1804),
.C(n_1299),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_SL g3793 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3793)
);

INVx4_ASAP7_75t_L g3794 ( 
.A(n_1914),
.Y(n_3794)
);

AOI22xp5_ASAP7_75t_L g3795 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3795)
);

A2O1A1Ixp33_ASAP7_75t_L g3796 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3796)
);

OAI22xp5_ASAP7_75t_L g3797 ( 
.A1(n_1859),
.A2(n_2317),
.B1(n_2318),
.B2(n_2279),
.Y(n_3797)
);

OAI22xp5_ASAP7_75t_L g3798 ( 
.A1(n_1859),
.A2(n_2317),
.B1(n_2318),
.B2(n_2279),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_2136),
.Y(n_3799)
);

AOI22xp5_ASAP7_75t_L g3800 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3800)
);

O2A1O1Ixp33_ASAP7_75t_L g3801 ( 
.A1(n_2282),
.A2(n_1220),
.B(n_2302),
.C(n_2299),
.Y(n_3801)
);

AOI22xp5_ASAP7_75t_L g3802 ( 
.A1(n_1896),
.A2(n_1859),
.B1(n_2317),
.B2(n_2279),
.Y(n_3802)
);

AND2x2_ASAP7_75t_L g3803 ( 
.A(n_1878),
.B(n_1897),
.Y(n_3803)
);

NOR2xp33_ASAP7_75t_SL g3804 ( 
.A(n_1920),
.B(n_1914),
.Y(n_3804)
);

OAI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3805)
);

INVxp67_ASAP7_75t_L g3806 ( 
.A(n_2090),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3807)
);

BUFx6f_ASAP7_75t_L g3808 ( 
.A(n_1914),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_1878),
.B(n_1897),
.Y(n_3809)
);

AOI21xp5_ASAP7_75t_L g3810 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3810)
);

OAI21xp5_ASAP7_75t_L g3811 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3811)
);

BUFx6f_ASAP7_75t_L g3812 ( 
.A(n_1914),
.Y(n_3812)
);

OAI21xp5_ASAP7_75t_L g3813 ( 
.A1(n_2284),
.A2(n_2359),
.B(n_2357),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3814)
);

AND2x2_ASAP7_75t_L g3815 ( 
.A(n_1878),
.B(n_1897),
.Y(n_3815)
);

AOI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3816)
);

AOI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3817)
);

BUFx6f_ASAP7_75t_L g3818 ( 
.A(n_1914),
.Y(n_3818)
);

BUFx2_ASAP7_75t_SL g3819 ( 
.A(n_1869),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_2045),
.B(n_1879),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_2304),
.A2(n_2703),
.B(n_2585),
.Y(n_3822)
);

BUFx6f_ASAP7_75t_L g3823 ( 
.A(n_1914),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_SL g3824 ( 
.A(n_1859),
.B(n_2279),
.Y(n_3824)
);

A2O1A1Ixp33_ASAP7_75t_L g3825 ( 
.A1(n_2535),
.A2(n_2669),
.B(n_2752),
.C(n_2556),
.Y(n_3825)
);

CKINVDCx5p33_ASAP7_75t_R g3826 ( 
.A(n_1905),
.Y(n_3826)
);

AND2x4_ASAP7_75t_SL g3827 ( 
.A(n_1920),
.B(n_2387),
.Y(n_3827)
);

INVx11_ASAP7_75t_L g3828 ( 
.A(n_1976),
.Y(n_3828)
);

INVxp67_ASAP7_75t_L g3829 ( 
.A(n_3218),
.Y(n_3829)
);

INVx2_ASAP7_75t_SL g3830 ( 
.A(n_2823),
.Y(n_3830)
);

AND2x4_ASAP7_75t_SL g3831 ( 
.A(n_2857),
.B(n_3576),
.Y(n_3831)
);

AOI22xp5_ASAP7_75t_L g3832 ( 
.A1(n_2890),
.A2(n_3580),
.B1(n_3605),
.B2(n_2901),
.Y(n_3832)
);

HB1xp67_ASAP7_75t_L g3833 ( 
.A(n_2913),
.Y(n_3833)
);

AOI22xp33_ASAP7_75t_L g3834 ( 
.A1(n_2890),
.A2(n_3605),
.B1(n_3627),
.B2(n_2901),
.Y(n_3834)
);

BUFx6f_ASAP7_75t_L g3835 ( 
.A(n_3782),
.Y(n_3835)
);

BUFx3_ASAP7_75t_L g3836 ( 
.A(n_3359),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_2896),
.B(n_2926),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_2896),
.B(n_2926),
.Y(n_3838)
);

BUFx12f_ASAP7_75t_L g3839 ( 
.A(n_3025),
.Y(n_3839)
);

INVx4_ASAP7_75t_L g3840 ( 
.A(n_3594),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_2832),
.B(n_2858),
.Y(n_3841)
);

AND2x4_ASAP7_75t_L g3842 ( 
.A(n_2823),
.B(n_2954),
.Y(n_3842)
);

BUFx2_ASAP7_75t_L g3843 ( 
.A(n_2823),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_2897),
.B(n_2917),
.Y(n_3844)
);

AND2x2_ASAP7_75t_L g3845 ( 
.A(n_2832),
.B(n_2858),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_2914),
.Y(n_3846)
);

CKINVDCx6p67_ASAP7_75t_R g3847 ( 
.A(n_3481),
.Y(n_3847)
);

BUFx6f_ASAP7_75t_L g3848 ( 
.A(n_3782),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_2897),
.B(n_2917),
.Y(n_3849)
);

CKINVDCx20_ASAP7_75t_R g3850 ( 
.A(n_2950),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_2914),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_2930),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_2930),
.Y(n_3853)
);

OR2x2_ASAP7_75t_L g3854 ( 
.A(n_3598),
.B(n_3713),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_2918),
.B(n_2827),
.Y(n_3855)
);

INVx6_ASAP7_75t_L g3856 ( 
.A(n_3526),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_2918),
.B(n_2836),
.Y(n_3857)
);

AND2x4_ASAP7_75t_L g3858 ( 
.A(n_2954),
.B(n_2960),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_2934),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_2837),
.B(n_2838),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_2840),
.B(n_2841),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_2845),
.B(n_2815),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_SL g3863 ( 
.A(n_3675),
.B(n_2807),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_2815),
.B(n_2819),
.Y(n_3864)
);

INVx5_ASAP7_75t_L g3865 ( 
.A(n_3509),
.Y(n_3865)
);

BUFx2_ASAP7_75t_L g3866 ( 
.A(n_2954),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_2832),
.B(n_2858),
.Y(n_3867)
);

INVxp67_ASAP7_75t_SL g3868 ( 
.A(n_2819),
.Y(n_3868)
);

INVx3_ASAP7_75t_L g3869 ( 
.A(n_2960),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3506),
.B(n_3508),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_SL g3871 ( 
.A(n_3675),
.B(n_2807),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_3506),
.B(n_3508),
.Y(n_3872)
);

HB1xp67_ASAP7_75t_L g3873 ( 
.A(n_3550),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_2934),
.Y(n_3874)
);

AND3x1_ASAP7_75t_SL g3875 ( 
.A(n_3788),
.B(n_3481),
.C(n_3626),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_2951),
.Y(n_3876)
);

OAI22xp5_ASAP7_75t_SL g3877 ( 
.A1(n_2809),
.A2(n_3562),
.B1(n_3570),
.B2(n_3524),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_2951),
.Y(n_3878)
);

BUFx3_ASAP7_75t_L g3879 ( 
.A(n_3359),
.Y(n_3879)
);

HB1xp67_ASAP7_75t_L g3880 ( 
.A(n_3669),
.Y(n_3880)
);

AOI22xp33_ASAP7_75t_L g3881 ( 
.A1(n_3580),
.A2(n_3627),
.B1(n_3699),
.B2(n_3788),
.Y(n_3881)
);

INVx4_ASAP7_75t_L g3882 ( 
.A(n_3594),
.Y(n_3882)
);

BUFx6f_ASAP7_75t_L g3883 ( 
.A(n_2810),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_2978),
.Y(n_3884)
);

A2O1A1Ixp33_ASAP7_75t_L g3885 ( 
.A1(n_2811),
.A2(n_2814),
.B(n_3699),
.C(n_3511),
.Y(n_3885)
);

INVx6_ASAP7_75t_L g3886 ( 
.A(n_3526),
.Y(n_3886)
);

INVxp67_ASAP7_75t_SL g3887 ( 
.A(n_3512),
.Y(n_3887)
);

HB1xp67_ASAP7_75t_L g3888 ( 
.A(n_3114),
.Y(n_3888)
);

AND2x4_ASAP7_75t_L g3889 ( 
.A(n_2960),
.B(n_2965),
.Y(n_3889)
);

INVx3_ASAP7_75t_L g3890 ( 
.A(n_2960),
.Y(n_3890)
);

OAI221xp5_ASAP7_75t_L g3891 ( 
.A1(n_3501),
.A2(n_3555),
.B1(n_3630),
.B2(n_3529),
.C(n_3522),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_SL g3892 ( 
.A(n_3497),
.B(n_3511),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_2978),
.Y(n_3893)
);

INVxp67_ASAP7_75t_L g3894 ( 
.A(n_3218),
.Y(n_3894)
);

INVx1_ASAP7_75t_SL g3895 ( 
.A(n_3819),
.Y(n_3895)
);

OR2x2_ASAP7_75t_SL g3896 ( 
.A(n_3533),
.B(n_3672),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3021),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3021),
.Y(n_3898)
);

OAI22xp33_ASAP7_75t_L g3899 ( 
.A1(n_3501),
.A2(n_3529),
.B1(n_3555),
.B2(n_3522),
.Y(n_3899)
);

INVx3_ASAP7_75t_L g3900 ( 
.A(n_2965),
.Y(n_3900)
);

BUFx2_ASAP7_75t_L g3901 ( 
.A(n_2965),
.Y(n_3901)
);

AND2x2_ASAP7_75t_L g3902 ( 
.A(n_2832),
.B(n_2858),
.Y(n_3902)
);

INVxp67_ASAP7_75t_L g3903 ( 
.A(n_3344),
.Y(n_3903)
);

AND3x1_ASAP7_75t_SL g3904 ( 
.A(n_3626),
.B(n_3600),
.C(n_3578),
.Y(n_3904)
);

BUFx6f_ASAP7_75t_L g3905 ( 
.A(n_2810),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3512),
.B(n_3513),
.Y(n_3906)
);

BUFx2_ASAP7_75t_L g3907 ( 
.A(n_3005),
.Y(n_3907)
);

NOR2xp33_ASAP7_75t_SL g3908 ( 
.A(n_3672),
.B(n_3497),
.Y(n_3908)
);

INVx1_ASAP7_75t_SL g3909 ( 
.A(n_3819),
.Y(n_3909)
);

CKINVDCx20_ASAP7_75t_R g3910 ( 
.A(n_3077),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3513),
.B(n_3514),
.Y(n_3911)
);

NOR2xp33_ASAP7_75t_L g3912 ( 
.A(n_3609),
.B(n_3615),
.Y(n_3912)
);

BUFx2_ASAP7_75t_SL g3913 ( 
.A(n_3536),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3514),
.B(n_3515),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3060),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_SL g3916 ( 
.A(n_3553),
.B(n_3575),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3060),
.Y(n_3917)
);

HB1xp67_ASAP7_75t_L g3918 ( 
.A(n_3114),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3080),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3080),
.Y(n_3920)
);

BUFx6f_ASAP7_75t_L g3921 ( 
.A(n_3171),
.Y(n_3921)
);

AO22x1_ASAP7_75t_L g3922 ( 
.A1(n_2887),
.A2(n_2927),
.B1(n_3592),
.B2(n_3575),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3515),
.B(n_3523),
.Y(n_3923)
);

BUFx6f_ASAP7_75t_L g3924 ( 
.A(n_3171),
.Y(n_3924)
);

CKINVDCx5p33_ASAP7_75t_R g3925 ( 
.A(n_3074),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3090),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3090),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3523),
.B(n_3525),
.Y(n_3928)
);

AO22x1_ASAP7_75t_L g3929 ( 
.A1(n_2887),
.A2(n_2927),
.B1(n_3592),
.B2(n_3553),
.Y(n_3929)
);

NOR2xp33_ASAP7_75t_L g3930 ( 
.A(n_3633),
.B(n_3652),
.Y(n_3930)
);

CKINVDCx5p33_ASAP7_75t_R g3931 ( 
.A(n_2813),
.Y(n_3931)
);

INVx2_ASAP7_75t_SL g3932 ( 
.A(n_3068),
.Y(n_3932)
);

NOR2x1p5_ASAP7_75t_L g3933 ( 
.A(n_2857),
.B(n_3576),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3525),
.B(n_3535),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3535),
.B(n_3540),
.Y(n_3935)
);

AOI22xp33_ASAP7_75t_L g3936 ( 
.A1(n_3131),
.A2(n_3146),
.B1(n_2856),
.B2(n_2878),
.Y(n_3936)
);

INVx5_ASAP7_75t_L g3937 ( 
.A(n_3509),
.Y(n_3937)
);

NAND2x1p5_ASAP7_75t_L g3938 ( 
.A(n_3311),
.B(n_3396),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3540),
.B(n_3547),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3547),
.B(n_3554),
.Y(n_3940)
);

NOR2x1_ASAP7_75t_R g3941 ( 
.A(n_2922),
.B(n_3025),
.Y(n_3941)
);

BUFx2_ASAP7_75t_L g3942 ( 
.A(n_3068),
.Y(n_3942)
);

HB1xp67_ASAP7_75t_L g3943 ( 
.A(n_2844),
.Y(n_3943)
);

NAND2x1p5_ASAP7_75t_L g3944 ( 
.A(n_3311),
.B(n_3396),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3554),
.B(n_3556),
.Y(n_3945)
);

INVx2_ASAP7_75t_SL g3946 ( 
.A(n_3093),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3101),
.Y(n_3947)
);

AND2x4_ASAP7_75t_L g3948 ( 
.A(n_3093),
.B(n_2876),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3101),
.Y(n_3949)
);

AND2x4_ASAP7_75t_L g3950 ( 
.A(n_3093),
.B(n_2876),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3556),
.B(n_3560),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3120),
.Y(n_3952)
);

CKINVDCx16_ASAP7_75t_R g3953 ( 
.A(n_3025),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3120),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3147),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3560),
.B(n_3564),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3147),
.Y(n_3957)
);

BUFx12f_ASAP7_75t_L g3958 ( 
.A(n_3096),
.Y(n_3958)
);

NOR2x1_ASAP7_75t_L g3959 ( 
.A(n_3174),
.B(n_2941),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3158),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3158),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3564),
.B(n_3566),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3189),
.Y(n_3963)
);

INVx5_ASAP7_75t_L g3964 ( 
.A(n_3509),
.Y(n_3964)
);

AND3x1_ASAP7_75t_SL g3965 ( 
.A(n_3663),
.B(n_3674),
.C(n_3667),
.Y(n_3965)
);

AOI22x1_ASAP7_75t_L g3966 ( 
.A1(n_3070),
.A2(n_3586),
.B1(n_3587),
.B2(n_3585),
.Y(n_3966)
);

NOR2xp33_ASAP7_75t_L g3967 ( 
.A(n_3702),
.B(n_3706),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_L g3968 ( 
.A(n_3566),
.B(n_3567),
.Y(n_3968)
);

BUFx2_ASAP7_75t_R g3969 ( 
.A(n_3002),
.Y(n_3969)
);

INVx2_ASAP7_75t_SL g3970 ( 
.A(n_2816),
.Y(n_3970)
);

INVx1_ASAP7_75t_SL g3971 ( 
.A(n_3598),
.Y(n_3971)
);

INVx3_ASAP7_75t_L g3972 ( 
.A(n_2816),
.Y(n_3972)
);

AND2x4_ASAP7_75t_L g3973 ( 
.A(n_2876),
.B(n_3013),
.Y(n_3973)
);

BUFx2_ASAP7_75t_L g3974 ( 
.A(n_2816),
.Y(n_3974)
);

AOI22xp5_ASAP7_75t_L g3975 ( 
.A1(n_2856),
.A2(n_2878),
.B1(n_2924),
.B2(n_2877),
.Y(n_3975)
);

BUFx3_ASAP7_75t_L g3976 ( 
.A(n_3359),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3567),
.B(n_3571),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3571),
.B(n_3588),
.Y(n_3978)
);

AOI22xp33_ASAP7_75t_L g3979 ( 
.A1(n_3131),
.A2(n_3146),
.B1(n_2877),
.B2(n_2924),
.Y(n_3979)
);

INVx4_ASAP7_75t_L g3980 ( 
.A(n_3594),
.Y(n_3980)
);

BUFx4f_ASAP7_75t_L g3981 ( 
.A(n_3584),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3205),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_SL g3983 ( 
.A(n_3610),
.B(n_3621),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3205),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3217),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3217),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3588),
.B(n_3590),
.Y(n_3987)
);

BUFx3_ASAP7_75t_L g3988 ( 
.A(n_3380),
.Y(n_3988)
);

OR2x2_ASAP7_75t_L g3989 ( 
.A(n_3713),
.B(n_3784),
.Y(n_3989)
);

INVx2_ASAP7_75t_SL g3990 ( 
.A(n_2816),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_3590),
.B(n_3593),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3593),
.B(n_3599),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3219),
.Y(n_3993)
);

BUFx2_ASAP7_75t_L g3994 ( 
.A(n_3528),
.Y(n_3994)
);

CKINVDCx5p33_ASAP7_75t_R g3995 ( 
.A(n_3300),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3599),
.B(n_3602),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_2843),
.Y(n_3997)
);

NOR2xp67_ASAP7_75t_L g3998 ( 
.A(n_3528),
.B(n_3691),
.Y(n_3998)
);

AOI22xp33_ASAP7_75t_L g3999 ( 
.A1(n_3499),
.A2(n_3563),
.B1(n_3695),
.B2(n_3532),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3219),
.Y(n_4000)
);

NAND2x1p5_ASAP7_75t_L g4001 ( 
.A(n_3311),
.B(n_3396),
.Y(n_4001)
);

BUFx8_ASAP7_75t_L g4002 ( 
.A(n_3431),
.Y(n_4002)
);

INVx2_ASAP7_75t_SL g4003 ( 
.A(n_3528),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_L g4004 ( 
.A(n_3602),
.B(n_3623),
.Y(n_4004)
);

AND2x4_ASAP7_75t_L g4005 ( 
.A(n_2876),
.B(n_3013),
.Y(n_4005)
);

OR2x2_ASAP7_75t_L g4006 ( 
.A(n_3784),
.B(n_2844),
.Y(n_4006)
);

INVx2_ASAP7_75t_L g4007 ( 
.A(n_2843),
.Y(n_4007)
);

A2O1A1Ixp33_ASAP7_75t_L g4008 ( 
.A1(n_3610),
.A2(n_3689),
.B(n_3712),
.C(n_3621),
.Y(n_4008)
);

INVxp67_ASAP7_75t_SL g4009 ( 
.A(n_3623),
.Y(n_4009)
);

HB1xp67_ASAP7_75t_L g4010 ( 
.A(n_3637),
.Y(n_4010)
);

AND2x2_ASAP7_75t_SL g4011 ( 
.A(n_3594),
.B(n_3772),
.Y(n_4011)
);

INVx4_ASAP7_75t_L g4012 ( 
.A(n_2850),
.Y(n_4012)
);

CKINVDCx5p33_ASAP7_75t_R g4013 ( 
.A(n_3196),
.Y(n_4013)
);

NOR2xp33_ASAP7_75t_SL g4014 ( 
.A(n_3689),
.B(n_3712),
.Y(n_4014)
);

AOI22xp5_ASAP7_75t_L g4015 ( 
.A1(n_3499),
.A2(n_3563),
.B1(n_3695),
.B2(n_3532),
.Y(n_4015)
);

BUFx2_ASAP7_75t_L g4016 ( 
.A(n_3528),
.Y(n_4016)
);

BUFx2_ASAP7_75t_L g4017 ( 
.A(n_3691),
.Y(n_4017)
);

INVx1_ASAP7_75t_SL g4018 ( 
.A(n_3368),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3637),
.B(n_3645),
.Y(n_4019)
);

AND2x4_ASAP7_75t_L g4020 ( 
.A(n_3013),
.B(n_3517),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_SL g4021 ( 
.A(n_3773),
.B(n_3805),
.Y(n_4021)
);

OAI221xp5_ASAP7_75t_L g4022 ( 
.A1(n_3630),
.A2(n_3710),
.B1(n_3717),
.B2(n_3648),
.C(n_3643),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3645),
.B(n_3646),
.Y(n_4023)
);

HB1xp67_ASAP7_75t_L g4024 ( 
.A(n_3646),
.Y(n_4024)
);

NOR2xp33_ASAP7_75t_L g4025 ( 
.A(n_3739),
.B(n_3740),
.Y(n_4025)
);

INVx3_ASAP7_75t_L g4026 ( 
.A(n_3691),
.Y(n_4026)
);

AOI22xp5_ASAP7_75t_L g4027 ( 
.A1(n_3715),
.A2(n_3732),
.B1(n_3798),
.B2(n_3797),
.Y(n_4027)
);

OAI22xp5_ASAP7_75t_L g4028 ( 
.A1(n_3643),
.A2(n_3710),
.B1(n_3717),
.B2(n_3648),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_L g4029 ( 
.A(n_3649),
.B(n_3651),
.Y(n_4029)
);

BUFx2_ASAP7_75t_L g4030 ( 
.A(n_3691),
.Y(n_4030)
);

BUFx4f_ASAP7_75t_L g4031 ( 
.A(n_3584),
.Y(n_4031)
);

NAND2xp33_ASAP7_75t_L g4032 ( 
.A(n_3773),
.B(n_3805),
.Y(n_4032)
);

INVx3_ASAP7_75t_L g4033 ( 
.A(n_3694),
.Y(n_4033)
);

HB1xp67_ASAP7_75t_L g4034 ( 
.A(n_3649),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3651),
.B(n_3657),
.Y(n_4035)
);

NOR2xp33_ASAP7_75t_L g4036 ( 
.A(n_3761),
.B(n_3767),
.Y(n_4036)
);

INVx2_ASAP7_75t_L g4037 ( 
.A(n_2885),
.Y(n_4037)
);

NAND2x1p5_ASAP7_75t_L g4038 ( 
.A(n_3311),
.B(n_3396),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3246),
.Y(n_4039)
);

NOR2xp33_ASAP7_75t_L g4040 ( 
.A(n_3765),
.B(n_3795),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3657),
.B(n_3666),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_3666),
.B(n_3668),
.Y(n_4042)
);

AOI221xp5_ASAP7_75t_L g4043 ( 
.A1(n_3715),
.A2(n_3732),
.B1(n_3798),
.B2(n_3797),
.C(n_3117),
.Y(n_4043)
);

AND2x4_ASAP7_75t_L g4044 ( 
.A(n_3013),
.B(n_3517),
.Y(n_4044)
);

INVx2_ASAP7_75t_L g4045 ( 
.A(n_2885),
.Y(n_4045)
);

INVx2_ASAP7_75t_L g4046 ( 
.A(n_2898),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3246),
.Y(n_4047)
);

AOI22x1_ASAP7_75t_L g4048 ( 
.A1(n_3585),
.A2(n_3587),
.B1(n_3607),
.B2(n_3586),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3247),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3668),
.B(n_3676),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3676),
.B(n_3678),
.Y(n_4051)
);

AND2x6_ASAP7_75t_L g4052 ( 
.A(n_2933),
.B(n_3000),
.Y(n_4052)
);

INVx2_ASAP7_75t_L g4053 ( 
.A(n_2898),
.Y(n_4053)
);

NOR2xp33_ASAP7_75t_L g4054 ( 
.A(n_3765),
.B(n_3795),
.Y(n_4054)
);

INVx1_ASAP7_75t_SL g4055 ( 
.A(n_3378),
.Y(n_4055)
);

BUFx3_ASAP7_75t_L g4056 ( 
.A(n_3380),
.Y(n_4056)
);

AOI22xp5_ASAP7_75t_L g4057 ( 
.A1(n_3802),
.A2(n_3800),
.B1(n_2853),
.B2(n_2910),
.Y(n_4057)
);

INVx4_ASAP7_75t_L g4058 ( 
.A(n_2850),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_3517),
.B(n_3518),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3247),
.Y(n_4060)
);

INVx1_ASAP7_75t_SL g4061 ( 
.A(n_3489),
.Y(n_4061)
);

INVx2_ASAP7_75t_L g4062 ( 
.A(n_2898),
.Y(n_4062)
);

BUFx2_ASAP7_75t_L g4063 ( 
.A(n_3694),
.Y(n_4063)
);

AND2x4_ASAP7_75t_L g4064 ( 
.A(n_3517),
.B(n_3518),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3678),
.B(n_3684),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_3518),
.B(n_3559),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3684),
.B(n_3693),
.Y(n_4067)
);

BUFx6f_ASAP7_75t_L g4068 ( 
.A(n_3171),
.Y(n_4068)
);

INVx5_ASAP7_75t_L g4069 ( 
.A(n_3509),
.Y(n_4069)
);

AND3x1_ASAP7_75t_L g4070 ( 
.A(n_2869),
.B(n_2920),
.C(n_2870),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3251),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3693),
.B(n_3697),
.Y(n_4072)
);

A2O1A1Ixp33_ASAP7_75t_L g4073 ( 
.A1(n_3811),
.A2(n_3813),
.B(n_3677),
.C(n_2846),
.Y(n_4073)
);

BUFx2_ASAP7_75t_L g4074 ( 
.A(n_3694),
.Y(n_4074)
);

BUFx2_ASAP7_75t_L g4075 ( 
.A(n_3694),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_SL g4076 ( 
.A(n_3811),
.B(n_3813),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3251),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3276),
.Y(n_4078)
);

AOI221x1_ASAP7_75t_L g4079 ( 
.A1(n_3569),
.A2(n_3742),
.B1(n_2820),
.B2(n_2849),
.C(n_2818),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_2902),
.Y(n_4080)
);

AOI22xp5_ASAP7_75t_L g4081 ( 
.A1(n_3800),
.A2(n_3802),
.B1(n_2919),
.B2(n_3498),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3697),
.B(n_3701),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_SL g4083 ( 
.A(n_3536),
.B(n_3601),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3701),
.B(n_3708),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3708),
.B(n_3718),
.Y(n_4085)
);

BUFx6f_ASAP7_75t_L g4086 ( 
.A(n_3171),
.Y(n_4086)
);

BUFx3_ASAP7_75t_L g4087 ( 
.A(n_3380),
.Y(n_4087)
);

BUFx3_ASAP7_75t_L g4088 ( 
.A(n_3518),
.Y(n_4088)
);

INVx3_ASAP7_75t_L g4089 ( 
.A(n_2857),
.Y(n_4089)
);

OR2x6_ASAP7_75t_L g4090 ( 
.A(n_3509),
.B(n_3624),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_SL g4091 ( 
.A(n_3601),
.B(n_3725),
.Y(n_4091)
);

INVx3_ASAP7_75t_L g4092 ( 
.A(n_2857),
.Y(n_4092)
);

NOR2xp33_ASAP7_75t_L g4093 ( 
.A(n_2998),
.B(n_2909),
.Y(n_4093)
);

BUFx12f_ASAP7_75t_L g4094 ( 
.A(n_3096),
.Y(n_4094)
);

NOR2xp33_ASAP7_75t_L g4095 ( 
.A(n_3520),
.B(n_3530),
.Y(n_4095)
);

BUFx4f_ASAP7_75t_L g4096 ( 
.A(n_3584),
.Y(n_4096)
);

BUFx4f_ASAP7_75t_L g4097 ( 
.A(n_3079),
.Y(n_4097)
);

CKINVDCx8_ASAP7_75t_R g4098 ( 
.A(n_2850),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3718),
.B(n_3722),
.Y(n_4099)
);

INVx1_ASAP7_75t_SL g4100 ( 
.A(n_3489),
.Y(n_4100)
);

AOI22xp5_ASAP7_75t_L g4101 ( 
.A1(n_3537),
.A2(n_3568),
.B1(n_3604),
.B2(n_3582),
.Y(n_4101)
);

AND2x2_ASAP7_75t_SL g4102 ( 
.A(n_3772),
.B(n_3758),
.Y(n_4102)
);

INVx3_ASAP7_75t_L g4103 ( 
.A(n_3576),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3722),
.B(n_3729),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3276),
.Y(n_4105)
);

HB1xp67_ASAP7_75t_SL g4106 ( 
.A(n_3051),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_SL g4107 ( 
.A(n_3725),
.B(n_3569),
.Y(n_4107)
);

HB1xp67_ASAP7_75t_L g4108 ( 
.A(n_3729),
.Y(n_4108)
);

AOI22xp5_ASAP7_75t_L g4109 ( 
.A1(n_3612),
.A2(n_3647),
.B1(n_3748),
.B2(n_3688),
.Y(n_4109)
);

HB1xp67_ASAP7_75t_L g4110 ( 
.A(n_3730),
.Y(n_4110)
);

HB1xp67_ASAP7_75t_L g4111 ( 
.A(n_3730),
.Y(n_4111)
);

AOI22xp5_ASAP7_75t_L g4112 ( 
.A1(n_3760),
.A2(n_3776),
.B1(n_3824),
.B2(n_3793),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_3287),
.Y(n_4113)
);

NOR2x1_ASAP7_75t_L g4114 ( 
.A(n_3174),
.B(n_2941),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3751),
.B(n_3755),
.Y(n_4115)
);

A2O1A1Ixp33_ASAP7_75t_L g4116 ( 
.A1(n_3742),
.A2(n_2821),
.B(n_3534),
.C(n_3519),
.Y(n_4116)
);

BUFx4f_ASAP7_75t_L g4117 ( 
.A(n_3079),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_3751),
.B(n_3755),
.Y(n_4118)
);

A2O1A1Ixp33_ASAP7_75t_L g4119 ( 
.A1(n_3581),
.A2(n_3613),
.B(n_3618),
.C(n_3596),
.Y(n_4119)
);

HB1xp67_ASAP7_75t_L g4120 ( 
.A(n_3756),
.Y(n_4120)
);

NOR2xp33_ASAP7_75t_L g4121 ( 
.A(n_3682),
.B(n_3696),
.Y(n_4121)
);

BUFx12f_ASAP7_75t_L g4122 ( 
.A(n_3096),
.Y(n_4122)
);

CKINVDCx8_ASAP7_75t_R g4123 ( 
.A(n_2850),
.Y(n_4123)
);

AOI22xp5_ASAP7_75t_L g4124 ( 
.A1(n_3117),
.A2(n_3145),
.B1(n_3154),
.B2(n_3133),
.Y(n_4124)
);

NOR2xp33_ASAP7_75t_L g4125 ( 
.A(n_3738),
.B(n_3787),
.Y(n_4125)
);

AND2x2_ASAP7_75t_L g4126 ( 
.A(n_3559),
.B(n_3595),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_3756),
.B(n_3759),
.Y(n_4127)
);

A2O1A1Ixp33_ASAP7_75t_L g4128 ( 
.A1(n_3653),
.A2(n_3681),
.B(n_3704),
.C(n_3665),
.Y(n_4128)
);

INVx2_ASAP7_75t_SL g4129 ( 
.A(n_3559),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_L g4130 ( 
.A(n_3759),
.B(n_3762),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3287),
.Y(n_4131)
);

CKINVDCx11_ASAP7_75t_R g4132 ( 
.A(n_2812),
.Y(n_4132)
);

AND2x4_ASAP7_75t_L g4133 ( 
.A(n_3595),
.B(n_2991),
.Y(n_4133)
);

A2O1A1Ixp33_ASAP7_75t_L g4134 ( 
.A1(n_3707),
.A2(n_3801),
.B(n_3757),
.C(n_2835),
.Y(n_4134)
);

AOI22xp33_ASAP7_75t_SL g4135 ( 
.A1(n_3145),
.A2(n_3180),
.B1(n_2867),
.B2(n_2828),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3762),
.B(n_3764),
.Y(n_4136)
);

AOI221x1_ASAP7_75t_L g4137 ( 
.A1(n_3607),
.A2(n_3622),
.B1(n_3629),
.B2(n_3620),
.C(n_3617),
.Y(n_4137)
);

INVx2_ASAP7_75t_SL g4138 ( 
.A(n_3595),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3764),
.B(n_3774),
.Y(n_4139)
);

NOR2xp33_ASAP7_75t_R g4140 ( 
.A(n_2923),
.B(n_2911),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_3774),
.B(n_3778),
.Y(n_4141)
);

CKINVDCx20_ASAP7_75t_R g4142 ( 
.A(n_3504),
.Y(n_4142)
);

INVx4_ASAP7_75t_L g4143 ( 
.A(n_2850),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_3778),
.B(n_3781),
.Y(n_4144)
);

NOR2xp33_ASAP7_75t_R g4145 ( 
.A(n_2923),
.B(n_2911),
.Y(n_4145)
);

INVx4_ASAP7_75t_L g4146 ( 
.A(n_2850),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_3781),
.B(n_3783),
.Y(n_4147)
);

HB1xp67_ASAP7_75t_L g4148 ( 
.A(n_3783),
.Y(n_4148)
);

AOI22xp33_ASAP7_75t_L g4149 ( 
.A1(n_3133),
.A2(n_3154),
.B1(n_3616),
.B2(n_2872),
.Y(n_4149)
);

AO22x1_ASAP7_75t_L g4150 ( 
.A1(n_3051),
.A2(n_3085),
.B1(n_3072),
.B2(n_2861),
.Y(n_4150)
);

BUFx4f_ASAP7_75t_L g4151 ( 
.A(n_3079),
.Y(n_4151)
);

OR2x6_ASAP7_75t_L g4152 ( 
.A(n_3624),
.B(n_2907),
.Y(n_4152)
);

INVxp67_ASAP7_75t_L g4153 ( 
.A(n_3344),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_2864),
.Y(n_4154)
);

INVx4_ASAP7_75t_L g4155 ( 
.A(n_2866),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_2864),
.Y(n_4156)
);

NOR2xp33_ASAP7_75t_L g4157 ( 
.A(n_3084),
.B(n_2872),
.Y(n_4157)
);

BUFx4f_ASAP7_75t_L g4158 ( 
.A(n_3079),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_2944),
.Y(n_4159)
);

INVxp67_ASAP7_75t_L g4160 ( 
.A(n_3503),
.Y(n_4160)
);

CKINVDCx5p33_ASAP7_75t_R g4161 ( 
.A(n_3248),
.Y(n_4161)
);

NAND3xp33_ASAP7_75t_L g4162 ( 
.A(n_2833),
.B(n_2852),
.C(n_2867),
.Y(n_4162)
);

HB1xp67_ASAP7_75t_L g4163 ( 
.A(n_3789),
.Y(n_4163)
);

HB1xp67_ASAP7_75t_L g4164 ( 
.A(n_3789),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_SL g4165 ( 
.A(n_3735),
.B(n_2830),
.Y(n_4165)
);

NAND2x1p5_ASAP7_75t_L g4166 ( 
.A(n_3036),
.B(n_3047),
.Y(n_4166)
);

AND2x2_ASAP7_75t_L g4167 ( 
.A(n_2970),
.B(n_2986),
.Y(n_4167)
);

INVx6_ASAP7_75t_L g4168 ( 
.A(n_3526),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_SL g4169 ( 
.A(n_3735),
.B(n_2921),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_3807),
.B(n_3814),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_2944),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_SL g4172 ( 
.A(n_2921),
.B(n_2839),
.Y(n_4172)
);

CKINVDCx20_ASAP7_75t_R g4173 ( 
.A(n_3700),
.Y(n_4173)
);

OR2x2_ASAP7_75t_L g4174 ( 
.A(n_3807),
.B(n_3814),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_3820),
.B(n_3821),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_2952),
.Y(n_4176)
);

AOI22x1_ASAP7_75t_L g4177 ( 
.A1(n_3617),
.A2(n_3622),
.B1(n_3629),
.B2(n_3620),
.Y(n_4177)
);

AND2x4_ASAP7_75t_L g4178 ( 
.A(n_2991),
.B(n_3526),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_3820),
.B(n_3821),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_2952),
.Y(n_4180)
);

NOR2xp33_ASAP7_75t_L g4181 ( 
.A(n_3084),
.B(n_2976),
.Y(n_4181)
);

OR2x2_ASAP7_75t_L g4182 ( 
.A(n_3223),
.B(n_2854),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_2992),
.Y(n_4183)
);

INVx2_ASAP7_75t_SL g4184 ( 
.A(n_3188),
.Y(n_4184)
);

BUFx2_ASAP7_75t_R g4185 ( 
.A(n_3492),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_2886),
.B(n_2903),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_2970),
.B(n_2986),
.Y(n_4187)
);

INVxp33_ASAP7_75t_SL g4188 ( 
.A(n_3143),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_3503),
.B(n_3670),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_3670),
.B(n_3753),
.Y(n_4190)
);

OAI21xp5_ASAP7_75t_L g4191 ( 
.A1(n_2851),
.A2(n_2860),
.B(n_2855),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_2992),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_2999),
.Y(n_4193)
);

AOI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_3109),
.A2(n_3112),
.B1(n_3105),
.B2(n_3082),
.Y(n_4194)
);

BUFx3_ASAP7_75t_L g4195 ( 
.A(n_2933),
.Y(n_4195)
);

CKINVDCx16_ASAP7_75t_R g4196 ( 
.A(n_3379),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_2999),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_3753),
.B(n_2889),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_3250),
.Y(n_4199)
);

HB1xp67_ASAP7_75t_L g4200 ( 
.A(n_3163),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_3057),
.B(n_3186),
.Y(n_4201)
);

NOR2x1p5_ASAP7_75t_L g4202 ( 
.A(n_3576),
.B(n_3591),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_L g4203 ( 
.A(n_3186),
.B(n_3193),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_3193),
.B(n_2997),
.Y(n_4204)
);

NAND2xp33_ASAP7_75t_R g4205 ( 
.A(n_3792),
.B(n_3624),
.Y(n_4205)
);

AND2x4_ASAP7_75t_L g4206 ( 
.A(n_3526),
.B(n_3412),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_2997),
.B(n_2966),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_2969),
.B(n_2971),
.Y(n_4208)
);

BUFx3_ASAP7_75t_L g4209 ( 
.A(n_2933),
.Y(n_4209)
);

A2O1A1Ixp33_ASAP7_75t_L g4210 ( 
.A1(n_3062),
.A2(n_3118),
.B(n_2871),
.C(n_2879),
.Y(n_4210)
);

BUFx2_ASAP7_75t_L g4211 ( 
.A(n_3624),
.Y(n_4211)
);

AOI22xp5_ASAP7_75t_L g4212 ( 
.A1(n_2939),
.A2(n_2946),
.B1(n_3107),
.B2(n_2883),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_2980),
.B(n_2989),
.Y(n_4213)
);

BUFx2_ASAP7_75t_L g4214 ( 
.A(n_3624),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_3250),
.Y(n_4215)
);

HB1xp67_ASAP7_75t_L g4216 ( 
.A(n_3163),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_2996),
.B(n_2891),
.Y(n_4217)
);

INVx3_ASAP7_75t_L g4218 ( 
.A(n_3591),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_SL g4219 ( 
.A(n_2839),
.B(n_2861),
.Y(n_4219)
);

INVx3_ASAP7_75t_L g4220 ( 
.A(n_3591),
.Y(n_4220)
);

AND2x4_ASAP7_75t_L g4221 ( 
.A(n_3412),
.B(n_3448),
.Y(n_4221)
);

INVx1_ASAP7_75t_SL g4222 ( 
.A(n_3487),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_SL g4223 ( 
.A(n_2884),
.B(n_3631),
.Y(n_4223)
);

AND2x2_ASAP7_75t_L g4224 ( 
.A(n_2990),
.B(n_3237),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_3244),
.Y(n_4225)
);

NOR2xp67_ASAP7_75t_L g4226 ( 
.A(n_3591),
.B(n_3791),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_2892),
.B(n_2900),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_3244),
.Y(n_4228)
);

BUFx12f_ASAP7_75t_L g4229 ( 
.A(n_3051),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_SL g4230 ( 
.A(n_3631),
.B(n_3632),
.Y(n_4230)
);

BUFx2_ASAP7_75t_L g4231 ( 
.A(n_3791),
.Y(n_4231)
);

BUFx8_ASAP7_75t_L g4232 ( 
.A(n_3431),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_2817),
.Y(n_4233)
);

CKINVDCx5p33_ASAP7_75t_R g4234 ( 
.A(n_2947),
.Y(n_4234)
);

AOI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_2939),
.A2(n_2946),
.B1(n_3107),
.B2(n_2865),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_2822),
.B(n_2829),
.Y(n_4236)
);

AND2x4_ASAP7_75t_L g4237 ( 
.A(n_3412),
.B(n_3448),
.Y(n_4237)
);

AND2x6_ASAP7_75t_L g4238 ( 
.A(n_2987),
.B(n_3000),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_2822),
.B(n_2829),
.Y(n_4239)
);

AND2x4_ASAP7_75t_L g4240 ( 
.A(n_3412),
.B(n_3448),
.Y(n_4240)
);

BUFx2_ASAP7_75t_L g4241 ( 
.A(n_3791),
.Y(n_4241)
);

INVx4_ASAP7_75t_L g4242 ( 
.A(n_2866),
.Y(n_4242)
);

INVx2_ASAP7_75t_SL g4243 ( 
.A(n_3188),
.Y(n_4243)
);

HB1xp67_ASAP7_75t_L g4244 ( 
.A(n_3252),
.Y(n_4244)
);

A2O1A1Ixp33_ASAP7_75t_L g4245 ( 
.A1(n_2916),
.A2(n_2961),
.B(n_3635),
.C(n_3632),
.Y(n_4245)
);

AOI22xp5_ASAP7_75t_L g4246 ( 
.A1(n_3160),
.A2(n_3180),
.B1(n_3119),
.B2(n_2932),
.Y(n_4246)
);

AOI22xp5_ASAP7_75t_L g4247 ( 
.A1(n_3160),
.A2(n_2945),
.B1(n_2958),
.B2(n_2957),
.Y(n_4247)
);

INVx4_ASAP7_75t_L g4248 ( 
.A(n_2866),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_L g4249 ( 
.A(n_2847),
.B(n_3577),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_SL g4250 ( 
.A(n_3635),
.B(n_3636),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_2847),
.B(n_3577),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_2817),
.Y(n_4252)
);

BUFx2_ASAP7_75t_L g4253 ( 
.A(n_3791),
.Y(n_4253)
);

BUFx3_ASAP7_75t_L g4254 ( 
.A(n_2987),
.Y(n_4254)
);

BUFx3_ASAP7_75t_L g4255 ( 
.A(n_2987),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_3589),
.B(n_3634),
.Y(n_4256)
);

BUFx2_ASAP7_75t_L g4257 ( 
.A(n_3794),
.Y(n_4257)
);

CKINVDCx5p33_ASAP7_75t_R g4258 ( 
.A(n_2947),
.Y(n_4258)
);

AOI22xp33_ASAP7_75t_L g4259 ( 
.A1(n_3121),
.A2(n_3033),
.B1(n_3058),
.B2(n_3086),
.Y(n_4259)
);

AOI22xp33_ASAP7_75t_L g4260 ( 
.A1(n_3058),
.A2(n_3086),
.B1(n_3312),
.B2(n_3235),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_3007),
.Y(n_4261)
);

BUFx3_ASAP7_75t_L g4262 ( 
.A(n_3000),
.Y(n_4262)
);

AND2x2_ASAP7_75t_L g4263 ( 
.A(n_2990),
.B(n_3237),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_3007),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_3115),
.Y(n_4265)
);

INVx2_ASAP7_75t_SL g4266 ( 
.A(n_3385),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_3589),
.B(n_3634),
.Y(n_4267)
);

AND2x4_ASAP7_75t_L g4268 ( 
.A(n_3448),
.B(n_3075),
.Y(n_4268)
);

NOR2xp67_ASAP7_75t_SL g4269 ( 
.A(n_3636),
.B(n_3638),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_3741),
.B(n_3745),
.Y(n_4270)
);

AND2x2_ASAP7_75t_L g4271 ( 
.A(n_3741),
.B(n_3745),
.Y(n_4271)
);

INVx3_ASAP7_75t_L g4272 ( 
.A(n_3794),
.Y(n_4272)
);

A2O1A1Ixp33_ASAP7_75t_L g4273 ( 
.A1(n_2961),
.A2(n_3640),
.B(n_3644),
.C(n_3638),
.Y(n_4273)
);

OA22x2_ASAP7_75t_L g4274 ( 
.A1(n_3202),
.A2(n_3495),
.B1(n_3330),
.B2(n_3178),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_SL g4275 ( 
.A(n_3640),
.B(n_3644),
.Y(n_4275)
);

HB1xp67_ASAP7_75t_L g4276 ( 
.A(n_3252),
.Y(n_4276)
);

AOI22x1_ASAP7_75t_L g4277 ( 
.A1(n_3654),
.A2(n_3656),
.B1(n_3658),
.B2(n_3655),
.Y(n_4277)
);

NAND2x1p5_ASAP7_75t_L g4278 ( 
.A(n_3036),
.B(n_3047),
.Y(n_4278)
);

AND2x2_ASAP7_75t_L g4279 ( 
.A(n_3763),
.B(n_3771),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_SL g4280 ( 
.A(n_3654),
.B(n_3655),
.Y(n_4280)
);

A2O1A1Ixp33_ASAP7_75t_L g4281 ( 
.A1(n_3656),
.A2(n_3659),
.B(n_3658),
.C(n_2967),
.Y(n_4281)
);

NOR2xp33_ASAP7_75t_R g4282 ( 
.A(n_3758),
.B(n_3777),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_3115),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3116),
.Y(n_4284)
);

BUFx4f_ASAP7_75t_SL g4285 ( 
.A(n_2922),
.Y(n_4285)
);

HB1xp67_ASAP7_75t_L g4286 ( 
.A(n_3259),
.Y(n_4286)
);

NOR2xp33_ASAP7_75t_L g4287 ( 
.A(n_3066),
.B(n_2973),
.Y(n_4287)
);

HB1xp67_ASAP7_75t_L g4288 ( 
.A(n_3259),
.Y(n_4288)
);

BUFx3_ASAP7_75t_L g4289 ( 
.A(n_3059),
.Y(n_4289)
);

AND2x4_ASAP7_75t_L g4290 ( 
.A(n_3076),
.B(n_3081),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_3763),
.B(n_3771),
.Y(n_4291)
);

BUFx3_ASAP7_75t_L g4292 ( 
.A(n_3059),
.Y(n_4292)
);

AND2x4_ASAP7_75t_L g4293 ( 
.A(n_3087),
.B(n_3091),
.Y(n_4293)
);

CKINVDCx16_ASAP7_75t_R g4294 ( 
.A(n_2922),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_3116),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_3775),
.B(n_3803),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_3775),
.B(n_3803),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_SL g4298 ( 
.A(n_3659),
.B(n_2808),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_3140),
.Y(n_4299)
);

NOR2xp33_ASAP7_75t_L g4300 ( 
.A(n_2973),
.B(n_2974),
.Y(n_4300)
);

OAI22xp5_ASAP7_75t_L g4301 ( 
.A1(n_2983),
.A2(n_3014),
.B1(n_3078),
.B2(n_3010),
.Y(n_4301)
);

INVx1_ASAP7_75t_SL g4302 ( 
.A(n_3487),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_3140),
.Y(n_4303)
);

OR2x6_ASAP7_75t_L g4304 ( 
.A(n_2908),
.B(n_2912),
.Y(n_4304)
);

NAND2xp33_ASAP7_75t_L g4305 ( 
.A(n_2806),
.B(n_3505),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_3175),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_3175),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_SL g4308 ( 
.A(n_3496),
.B(n_3500),
.Y(n_4308)
);

BUFx4f_ASAP7_75t_L g4309 ( 
.A(n_3079),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_SL g4310 ( 
.A(n_3502),
.B(n_3507),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_3809),
.B(n_3815),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_3181),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_3809),
.B(n_3815),
.Y(n_4313)
);

NOR2xp33_ASAP7_75t_R g4314 ( 
.A(n_3777),
.B(n_3804),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_3064),
.B(n_3100),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_L g4316 ( 
.A(n_2859),
.B(n_2862),
.Y(n_4316)
);

NOR2xp33_ASAP7_75t_L g4317 ( 
.A(n_2974),
.B(n_2981),
.Y(n_4317)
);

NOR2xp33_ASAP7_75t_R g4318 ( 
.A(n_3804),
.B(n_3558),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_SL g4319 ( 
.A(n_3521),
.B(n_3527),
.Y(n_4319)
);

INVx5_ASAP7_75t_L g4320 ( 
.A(n_2866),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_2859),
.B(n_2862),
.Y(n_4321)
);

HB1xp67_ASAP7_75t_L g4322 ( 
.A(n_3265),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_SL g4323 ( 
.A(n_3531),
.B(n_3538),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_3006),
.B(n_3008),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_3009),
.B(n_3012),
.Y(n_4325)
);

BUFx8_ASAP7_75t_L g4326 ( 
.A(n_3431),
.Y(n_4326)
);

OR2x2_ASAP7_75t_L g4327 ( 
.A(n_3223),
.B(n_2854),
.Y(n_4327)
);

HB1xp67_ASAP7_75t_L g4328 ( 
.A(n_3265),
.Y(n_4328)
);

AOI22xp33_ASAP7_75t_L g4329 ( 
.A1(n_3312),
.A2(n_3235),
.B1(n_3495),
.B2(n_3031),
.Y(n_4329)
);

NOR2xp33_ASAP7_75t_L g4330 ( 
.A(n_2981),
.B(n_3031),
.Y(n_4330)
);

BUFx3_ASAP7_75t_L g4331 ( 
.A(n_3059),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_SL g4332 ( 
.A(n_3539),
.B(n_3541),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_3157),
.B(n_3159),
.Y(n_4333)
);

HB1xp67_ASAP7_75t_L g4334 ( 
.A(n_3279),
.Y(n_4334)
);

AND2x4_ASAP7_75t_L g4335 ( 
.A(n_3106),
.B(n_3198),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_L g4336 ( 
.A(n_3161),
.B(n_3162),
.Y(n_4336)
);

HB1xp67_ASAP7_75t_L g4337 ( 
.A(n_3279),
.Y(n_4337)
);

NOR2xp33_ASAP7_75t_L g4338 ( 
.A(n_3041),
.B(n_3046),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_2904),
.Y(n_4339)
);

BUFx3_ASAP7_75t_L g4340 ( 
.A(n_3272),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_3166),
.B(n_3177),
.Y(n_4341)
);

BUFx2_ASAP7_75t_L g4342 ( 
.A(n_3794),
.Y(n_4342)
);

OR2x2_ASAP7_75t_L g4343 ( 
.A(n_3241),
.B(n_3221),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_2906),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_SL g4345 ( 
.A(n_3542),
.B(n_3543),
.Y(n_4345)
);

INVxp67_ASAP7_75t_SL g4346 ( 
.A(n_3185),
.Y(n_4346)
);

OR2x2_ASAP7_75t_SL g4347 ( 
.A(n_2866),
.B(n_3660),
.Y(n_4347)
);

BUFx2_ASAP7_75t_L g4348 ( 
.A(n_2866),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_3183),
.B(n_2824),
.Y(n_4349)
);

INVxp33_ASAP7_75t_L g4350 ( 
.A(n_3332),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_2824),
.B(n_2825),
.Y(n_4351)
);

AND2x2_ASAP7_75t_L g4352 ( 
.A(n_3290),
.B(n_3298),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_2825),
.B(n_2826),
.Y(n_4353)
);

OAI22xp5_ASAP7_75t_SL g4354 ( 
.A1(n_3202),
.A2(n_3046),
.B1(n_3041),
.B2(n_3494),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_3290),
.B(n_3298),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_L g4356 ( 
.A(n_2826),
.B(n_2831),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_L g4357 ( 
.A(n_2831),
.B(n_2842),
.Y(n_4357)
);

BUFx2_ASAP7_75t_L g4358 ( 
.A(n_3660),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_2842),
.B(n_2848),
.Y(n_4359)
);

CKINVDCx6p67_ASAP7_75t_R g4360 ( 
.A(n_3546),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_2848),
.B(n_2928),
.Y(n_4361)
);

AOI22xp33_ASAP7_75t_L g4362 ( 
.A1(n_3480),
.A2(n_2863),
.B1(n_2880),
.B2(n_2873),
.Y(n_4362)
);

BUFx12f_ASAP7_75t_L g4363 ( 
.A(n_3051),
.Y(n_4363)
);

NAND2xp5_ASAP7_75t_L g4364 ( 
.A(n_2928),
.B(n_2931),
.Y(n_4364)
);

AOI22xp5_ASAP7_75t_L g4365 ( 
.A1(n_3011),
.A2(n_3022),
.B1(n_3045),
.B2(n_2899),
.Y(n_4365)
);

AND3x1_ASAP7_75t_SL g4366 ( 
.A(n_3606),
.B(n_3828),
.C(n_3092),
.Y(n_4366)
);

OR2x2_ASAP7_75t_L g4367 ( 
.A(n_3241),
.B(n_3221),
.Y(n_4367)
);

HB1xp67_ASAP7_75t_L g4368 ( 
.A(n_3284),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_L g4369 ( 
.A(n_2931),
.B(n_2937),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_L g4370 ( 
.A(n_2937),
.B(n_2942),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_SL g4371 ( 
.A(n_3545),
.B(n_3548),
.Y(n_4371)
);

NOR2xp33_ASAP7_75t_L g4372 ( 
.A(n_2962),
.B(n_2863),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_2942),
.B(n_2955),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_2955),
.B(n_2956),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_SL g4375 ( 
.A(n_3551),
.B(n_3552),
.Y(n_4375)
);

NAND2x1p5_ASAP7_75t_L g4376 ( 
.A(n_3036),
.B(n_3047),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_L g4377 ( 
.A(n_2956),
.B(n_2964),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_2964),
.B(n_2968),
.Y(n_4378)
);

BUFx2_ASAP7_75t_L g4379 ( 
.A(n_3660),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_2968),
.B(n_2972),
.Y(n_4380)
);

AOI22xp5_ASAP7_75t_L g4381 ( 
.A1(n_2868),
.A2(n_2874),
.B1(n_2895),
.B2(n_2888),
.Y(n_4381)
);

CKINVDCx5p33_ASAP7_75t_R g4382 ( 
.A(n_3606),
.Y(n_4382)
);

INVxp67_ASAP7_75t_L g4383 ( 
.A(n_2949),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_L g4384 ( 
.A(n_2972),
.B(n_2979),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_2979),
.B(n_2982),
.Y(n_4385)
);

BUFx3_ASAP7_75t_L g4386 ( 
.A(n_3272),
.Y(n_4386)
);

NOR2xp33_ASAP7_75t_L g4387 ( 
.A(n_2962),
.B(n_2873),
.Y(n_4387)
);

HB1xp67_ASAP7_75t_L g4388 ( 
.A(n_3284),
.Y(n_4388)
);

NAND2xp5_ASAP7_75t_L g4389 ( 
.A(n_2982),
.B(n_2988),
.Y(n_4389)
);

OAI22xp5_ASAP7_75t_L g4390 ( 
.A1(n_2977),
.A2(n_3038),
.B1(n_3043),
.B2(n_3023),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_L g4391 ( 
.A(n_2988),
.B(n_2993),
.Y(n_4391)
);

INVx2_ASAP7_75t_SL g4392 ( 
.A(n_3385),
.Y(n_4392)
);

NOR2xp33_ASAP7_75t_SL g4393 ( 
.A(n_3072),
.B(n_3085),
.Y(n_4393)
);

OR2x6_ASAP7_75t_L g4394 ( 
.A(n_2915),
.B(n_2925),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_L g4395 ( 
.A(n_2993),
.B(n_2994),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_L g4396 ( 
.A(n_2994),
.B(n_3001),
.Y(n_4396)
);

CKINVDCx6p67_ASAP7_75t_R g4397 ( 
.A(n_3546),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_3001),
.B(n_3003),
.Y(n_4398)
);

INVx2_ASAP7_75t_SL g4399 ( 
.A(n_3385),
.Y(n_4399)
);

INVxp67_ASAP7_75t_SL g4400 ( 
.A(n_3185),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_3003),
.B(n_3004),
.Y(n_4401)
);

INVx5_ASAP7_75t_L g4402 ( 
.A(n_3660),
.Y(n_4402)
);

INVxp67_ASAP7_75t_L g4403 ( 
.A(n_2995),
.Y(n_4403)
);

INVx1_ASAP7_75t_SL g4404 ( 
.A(n_3052),
.Y(n_4404)
);

BUFx3_ASAP7_75t_L g4405 ( 
.A(n_3272),
.Y(n_4405)
);

NOR2xp33_ASAP7_75t_L g4406 ( 
.A(n_2880),
.B(n_2882),
.Y(n_4406)
);

OR2x2_ASAP7_75t_L g4407 ( 
.A(n_3229),
.B(n_3260),
.Y(n_4407)
);

NOR2xp67_ASAP7_75t_L g4408 ( 
.A(n_3557),
.B(n_3561),
.Y(n_4408)
);

NOR2xp33_ASAP7_75t_L g4409 ( 
.A(n_2882),
.B(n_3040),
.Y(n_4409)
);

NAND2xp5_ASAP7_75t_L g4410 ( 
.A(n_3004),
.B(n_3016),
.Y(n_4410)
);

HB1xp67_ASAP7_75t_L g4411 ( 
.A(n_3260),
.Y(n_4411)
);

OAI21xp5_ASAP7_75t_L g4412 ( 
.A1(n_3510),
.A2(n_3549),
.B(n_3544),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_3016),
.B(n_3026),
.Y(n_4413)
);

CKINVDCx5p33_ASAP7_75t_R g4414 ( 
.A(n_3828),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_3026),
.B(n_3028),
.Y(n_4415)
);

NAND2xp5_ASAP7_75t_L g4416 ( 
.A(n_3028),
.B(n_3029),
.Y(n_4416)
);

NAND2xp5_ASAP7_75t_L g4417 ( 
.A(n_3029),
.B(n_3037),
.Y(n_4417)
);

INVx2_ASAP7_75t_SL g4418 ( 
.A(n_3385),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_3037),
.B(n_3044),
.Y(n_4419)
);

NAND2x1p5_ASAP7_75t_L g4420 ( 
.A(n_3036),
.B(n_3047),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_L g4421 ( 
.A(n_3044),
.B(n_3048),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_3048),
.B(n_3073),
.Y(n_4422)
);

AND2x4_ASAP7_75t_L g4423 ( 
.A(n_3106),
.B(n_3198),
.Y(n_4423)
);

BUFx3_ASAP7_75t_L g4424 ( 
.A(n_3273),
.Y(n_4424)
);

BUFx4f_ASAP7_75t_L g4425 ( 
.A(n_3079),
.Y(n_4425)
);

OR2x2_ASAP7_75t_L g4426 ( 
.A(n_3229),
.B(n_3267),
.Y(n_4426)
);

AOI22xp5_ASAP7_75t_L g4427 ( 
.A1(n_2984),
.A2(n_2977),
.B1(n_3038),
.B2(n_3023),
.Y(n_4427)
);

AND2x4_ASAP7_75t_L g4428 ( 
.A(n_3106),
.B(n_3198),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_3073),
.B(n_3083),
.Y(n_4429)
);

BUFx2_ASAP7_75t_L g4430 ( 
.A(n_3660),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_SL g4431 ( 
.A(n_3565),
.B(n_3572),
.Y(n_4431)
);

AND2x2_ASAP7_75t_SL g4432 ( 
.A(n_3827),
.B(n_3280),
.Y(n_4432)
);

A2O1A1Ixp33_ASAP7_75t_L g4433 ( 
.A1(n_3069),
.A2(n_3573),
.B(n_3579),
.C(n_3574),
.Y(n_4433)
);

HB1xp67_ASAP7_75t_L g4434 ( 
.A(n_3267),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_SL g4435 ( 
.A(n_3583),
.B(n_3664),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_3083),
.B(n_3088),
.Y(n_4436)
);

OR2x2_ASAP7_75t_L g4437 ( 
.A(n_3269),
.B(n_3278),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_SL g4438 ( 
.A(n_3671),
.B(n_3673),
.Y(n_4438)
);

BUFx2_ASAP7_75t_L g4439 ( 
.A(n_3662),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_L g4440 ( 
.A(n_3088),
.B(n_3089),
.Y(n_4440)
);

BUFx3_ASAP7_75t_L g4441 ( 
.A(n_3273),
.Y(n_4441)
);

INVx6_ASAP7_75t_L g4442 ( 
.A(n_3072),
.Y(n_4442)
);

AND2x4_ASAP7_75t_L g4443 ( 
.A(n_3345),
.B(n_3355),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_3611),
.Y(n_4444)
);

NAND2xp5_ASAP7_75t_L g4445 ( 
.A(n_3089),
.B(n_3095),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_L g4446 ( 
.A(n_3095),
.B(n_3097),
.Y(n_4446)
);

CKINVDCx5p33_ASAP7_75t_R g4447 ( 
.A(n_3687),
.Y(n_4447)
);

OR2x2_ASAP7_75t_L g4448 ( 
.A(n_3269),
.B(n_3278),
.Y(n_4448)
);

AND2x4_ASAP7_75t_L g4449 ( 
.A(n_3345),
.B(n_3355),
.Y(n_4449)
);

AND2x4_ASAP7_75t_L g4450 ( 
.A(n_3357),
.B(n_3362),
.Y(n_4450)
);

AND2x2_ASAP7_75t_SL g4451 ( 
.A(n_3827),
.B(n_3358),
.Y(n_4451)
);

OR2x2_ASAP7_75t_L g4452 ( 
.A(n_3097),
.B(n_3098),
.Y(n_4452)
);

AND3x1_ASAP7_75t_SL g4453 ( 
.A(n_3642),
.B(n_3650),
.C(n_3692),
.Y(n_4453)
);

NOR2xp33_ASAP7_75t_SL g4454 ( 
.A(n_3072),
.B(n_3085),
.Y(n_4454)
);

CKINVDCx8_ASAP7_75t_R g4455 ( 
.A(n_3662),
.Y(n_4455)
);

NOR2xp33_ASAP7_75t_L g4456 ( 
.A(n_2985),
.B(n_3043),
.Y(n_4456)
);

INVxp67_ASAP7_75t_L g4457 ( 
.A(n_3132),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_3098),
.B(n_3102),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_SL g4459 ( 
.A(n_3680),
.B(n_3690),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_L g4460 ( 
.A(n_3102),
.B(n_3103),
.Y(n_4460)
);

INVx2_ASAP7_75t_SL g4461 ( 
.A(n_3424),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_L g4462 ( 
.A(n_3103),
.B(n_3104),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_L g4463 ( 
.A(n_3104),
.B(n_3111),
.Y(n_4463)
);

AOI22xp5_ASAP7_75t_L g4464 ( 
.A1(n_3056),
.A2(n_3135),
.B1(n_3148),
.B2(n_3035),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_L g4465 ( 
.A(n_3111),
.B(n_3113),
.Y(n_4465)
);

AOI221xp5_ASAP7_75t_L g4466 ( 
.A1(n_3027),
.A2(n_3049),
.B1(n_3054),
.B2(n_3053),
.C(n_3124),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_3113),
.B(n_3126),
.Y(n_4467)
);

INVx2_ASAP7_75t_SL g4468 ( 
.A(n_3424),
.Y(n_4468)
);

AOI22xp5_ASAP7_75t_L g4469 ( 
.A1(n_3056),
.A2(n_3042),
.B1(n_3039),
.B2(n_3015),
.Y(n_4469)
);

NOR2x1_ASAP7_75t_L g4470 ( 
.A(n_2959),
.B(n_3153),
.Y(n_4470)
);

NOR2xp33_ASAP7_75t_L g4471 ( 
.A(n_3168),
.B(n_3125),
.Y(n_4471)
);

AND2x4_ASAP7_75t_L g4472 ( 
.A(n_3357),
.B(n_3362),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_L g4473 ( 
.A(n_3126),
.B(n_3128),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_SL g4474 ( 
.A(n_3711),
.B(n_3716),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_3128),
.B(n_3139),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_3139),
.B(n_3141),
.Y(n_4476)
);

NOR2xp33_ASAP7_75t_L g4477 ( 
.A(n_2953),
.B(n_3061),
.Y(n_4477)
);

AND2x2_ASAP7_75t_L g4478 ( 
.A(n_3799),
.B(n_3779),
.Y(n_4478)
);

HB1xp67_ASAP7_75t_L g4479 ( 
.A(n_2834),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_3141),
.B(n_3142),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_L g4481 ( 
.A(n_3142),
.B(n_3150),
.Y(n_4481)
);

NAND2xp33_ASAP7_75t_L g4482 ( 
.A(n_3597),
.B(n_3608),
.Y(n_4482)
);

OAI21xp5_ASAP7_75t_L g4483 ( 
.A1(n_3628),
.A2(n_3683),
.B(n_3639),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_3435),
.Y(n_4484)
);

AND2x6_ASAP7_75t_L g4485 ( 
.A(n_3273),
.B(n_3320),
.Y(n_4485)
);

BUFx2_ASAP7_75t_SL g4486 ( 
.A(n_2936),
.Y(n_4486)
);

AND2x4_ASAP7_75t_L g4487 ( 
.A(n_3320),
.B(n_3703),
.Y(n_4487)
);

BUFx2_ASAP7_75t_L g4488 ( 
.A(n_3779),
.Y(n_4488)
);

INVx2_ASAP7_75t_SL g4489 ( 
.A(n_3424),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_3435),
.Y(n_4490)
);

NAND2xp33_ASAP7_75t_SL g4491 ( 
.A(n_3779),
.B(n_3808),
.Y(n_4491)
);

INVx5_ASAP7_75t_L g4492 ( 
.A(n_3779),
.Y(n_4492)
);

AOI21xp5_ASAP7_75t_L g4493 ( 
.A1(n_3719),
.A2(n_3723),
.B(n_3720),
.Y(n_4493)
);

O2A1O1Ixp33_ASAP7_75t_L g4494 ( 
.A1(n_3685),
.A2(n_3686),
.B(n_3728),
.C(n_3698),
.Y(n_4494)
);

INVxp67_ASAP7_75t_SL g4495 ( 
.A(n_3194),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_L g4496 ( 
.A(n_3150),
.B(n_3152),
.Y(n_4496)
);

BUFx2_ASAP7_75t_L g4497 ( 
.A(n_3808),
.Y(n_4497)
);

NOR2xp33_ASAP7_75t_SL g4498 ( 
.A(n_3085),
.B(n_2963),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_3277),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_SL g4500 ( 
.A(n_3724),
.B(n_3726),
.Y(n_4500)
);

INVxp67_ASAP7_75t_L g4501 ( 
.A(n_3063),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_SL g4502 ( 
.A(n_3727),
.B(n_3731),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_3281),
.Y(n_4503)
);

AOI221xp5_ASAP7_75t_L g4504 ( 
.A1(n_3124),
.A2(n_3015),
.B1(n_3055),
.B2(n_3050),
.C(n_3032),
.Y(n_4504)
);

AND3x1_ASAP7_75t_SL g4505 ( 
.A(n_3734),
.B(n_3826),
.C(n_3143),
.Y(n_4505)
);

BUFx2_ASAP7_75t_L g4506 ( 
.A(n_3808),
.Y(n_4506)
);

BUFx2_ASAP7_75t_L g4507 ( 
.A(n_3812),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_3152),
.B(n_3155),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_3155),
.B(n_3165),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_3165),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_SL g4511 ( 
.A(n_3733),
.B(n_3736),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_3169),
.B(n_3170),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_L g4513 ( 
.A(n_3169),
.B(n_3170),
.Y(n_4513)
);

NAND2x1p5_ASAP7_75t_L g4514 ( 
.A(n_3389),
.B(n_3320),
.Y(n_4514)
);

HB1xp67_ASAP7_75t_L g4515 ( 
.A(n_2834),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_L g4516 ( 
.A(n_3176),
.B(n_3199),
.Y(n_4516)
);

INVx5_ASAP7_75t_L g4517 ( 
.A(n_3812),
.Y(n_4517)
);

AOI21xp5_ASAP7_75t_L g4518 ( 
.A1(n_3744),
.A2(n_3754),
.B(n_3746),
.Y(n_4518)
);

HB1xp67_ASAP7_75t_L g4519 ( 
.A(n_3406),
.Y(n_4519)
);

BUFx2_ASAP7_75t_L g4520 ( 
.A(n_3812),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_3176),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_3199),
.B(n_3203),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_L g4523 ( 
.A(n_3203),
.B(n_3110),
.Y(n_4523)
);

NAND2xp5_ASAP7_75t_L g4524 ( 
.A(n_3292),
.B(n_3294),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_3212),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_3212),
.Y(n_4526)
);

INVxp33_ASAP7_75t_L g4527 ( 
.A(n_3351),
.Y(n_4527)
);

AOI22xp5_ASAP7_75t_L g4528 ( 
.A1(n_3032),
.A2(n_3050),
.B1(n_3055),
.B2(n_3151),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_3292),
.B(n_3294),
.Y(n_4529)
);

INVxp67_ASAP7_75t_SL g4530 ( 
.A(n_3194),
.Y(n_4530)
);

INVx1_ASAP7_75t_L g4531 ( 
.A(n_3226),
.Y(n_4531)
);

BUFx3_ASAP7_75t_L g4532 ( 
.A(n_3703),
.Y(n_4532)
);

HB1xp67_ASAP7_75t_L g4533 ( 
.A(n_3406),
.Y(n_4533)
);

AND2x4_ASAP7_75t_L g4534 ( 
.A(n_3703),
.B(n_3705),
.Y(n_4534)
);

NAND2xp5_ASAP7_75t_SL g4535 ( 
.A(n_3766),
.B(n_3769),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_3226),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_3234),
.Y(n_4537)
);

CKINVDCx14_ASAP7_75t_R g4538 ( 
.A(n_3240),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_3306),
.B(n_3313),
.Y(n_4539)
);

CKINVDCx5p33_ASAP7_75t_R g4540 ( 
.A(n_3289),
.Y(n_4540)
);

AND2x2_ASAP7_75t_L g4541 ( 
.A(n_3818),
.B(n_3823),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_L g4542 ( 
.A(n_3306),
.B(n_3313),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_SL g4543 ( 
.A(n_3770),
.B(n_3785),
.Y(n_4543)
);

NOR2xp33_ASAP7_75t_L g4544 ( 
.A(n_3806),
.B(n_3024),
.Y(n_4544)
);

OAI22xp5_ASAP7_75t_L g4545 ( 
.A1(n_3737),
.A2(n_3752),
.B1(n_3796),
.B2(n_3749),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_SL g4546 ( 
.A(n_3786),
.B(n_3810),
.Y(n_4546)
);

CKINVDCx5p33_ASAP7_75t_R g4547 ( 
.A(n_3768),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_3234),
.Y(n_4548)
);

OR2x6_ASAP7_75t_L g4549 ( 
.A(n_3705),
.B(n_3747),
.Y(n_4549)
);

NAND2xp5_ASAP7_75t_L g4550 ( 
.A(n_3317),
.B(n_3321),
.Y(n_4550)
);

OR2x2_ASAP7_75t_L g4551 ( 
.A(n_3094),
.B(n_3099),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_3408),
.Y(n_4552)
);

BUFx3_ASAP7_75t_L g4553 ( 
.A(n_3705),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_3317),
.B(n_3321),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_3325),
.B(n_3326),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_3408),
.Y(n_4556)
);

INVx1_ASAP7_75t_SL g4557 ( 
.A(n_3052),
.Y(n_4557)
);

BUFx3_ASAP7_75t_L g4558 ( 
.A(n_3747),
.Y(n_4558)
);

A2O1A1Ixp33_ASAP7_75t_L g4559 ( 
.A1(n_3816),
.A2(n_3817),
.B(n_3822),
.C(n_3825),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_SL g4560 ( 
.A(n_2959),
.B(n_2936),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_3325),
.B(n_3326),
.Y(n_4561)
);

INVx1_ASAP7_75t_SL g4562 ( 
.A(n_3052),
.Y(n_4562)
);

NAND2xp5_ASAP7_75t_L g4563 ( 
.A(n_3017),
.B(n_3231),
.Y(n_4563)
);

NOR2xp33_ASAP7_75t_L g4564 ( 
.A(n_3206),
.B(n_3153),
.Y(n_4564)
);

AO221x1_ASAP7_75t_L g4565 ( 
.A1(n_2875),
.A2(n_2894),
.B1(n_3823),
.B2(n_3818),
.C(n_3472),
.Y(n_4565)
);

AND3x1_ASAP7_75t_SL g4566 ( 
.A(n_3204),
.B(n_3480),
.C(n_3197),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_SL g4567 ( 
.A(n_2875),
.B(n_2894),
.Y(n_4567)
);

AND2x4_ASAP7_75t_L g4568 ( 
.A(n_3747),
.B(n_3827),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_3231),
.B(n_2943),
.Y(n_4569)
);

NAND2xp5_ASAP7_75t_L g4570 ( 
.A(n_3178),
.B(n_3258),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_L g4571 ( 
.A(n_2948),
.B(n_3410),
.Y(n_4571)
);

NAND2xp5_ASAP7_75t_SL g4572 ( 
.A(n_2875),
.B(n_2894),
.Y(n_4572)
);

AOI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_3310),
.A2(n_3071),
.B(n_3282),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_3303),
.Y(n_4574)
);

NAND2x1p5_ASAP7_75t_L g4575 ( 
.A(n_3389),
.B(n_3823),
.Y(n_4575)
);

CKINVDCx11_ASAP7_75t_R g4576 ( 
.A(n_3308),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_SL g4577 ( 
.A(n_2875),
.B(n_2894),
.Y(n_4577)
);

NAND2xp5_ASAP7_75t_L g4578 ( 
.A(n_3410),
.B(n_2929),
.Y(n_4578)
);

NAND3xp33_ASAP7_75t_L g4579 ( 
.A(n_2893),
.B(n_3191),
.C(n_3130),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_L g4580 ( 
.A(n_2935),
.B(n_2938),
.Y(n_4580)
);

BUFx3_ASAP7_75t_L g4581 ( 
.A(n_2875),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_2940),
.B(n_3436),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_SL g4583 ( 
.A(n_2875),
.B(n_2894),
.Y(n_4583)
);

AOI21xp5_ASAP7_75t_L g4584 ( 
.A1(n_3310),
.A2(n_3293),
.B(n_3283),
.Y(n_4584)
);

INVx2_ASAP7_75t_SL g4585 ( 
.A(n_3424),
.Y(n_4585)
);

HB1xp67_ASAP7_75t_L g4586 ( 
.A(n_2905),
.Y(n_4586)
);

CKINVDCx5p33_ASAP7_75t_R g4587 ( 
.A(n_3768),
.Y(n_4587)
);

AND3x2_ASAP7_75t_SL g4588 ( 
.A(n_3363),
.B(n_3339),
.C(n_3361),
.Y(n_4588)
);

BUFx2_ASAP7_75t_L g4589 ( 
.A(n_3424),
.Y(n_4589)
);

OAI22xp5_ASAP7_75t_L g4590 ( 
.A1(n_3330),
.A2(n_3318),
.B1(n_3137),
.B2(n_3144),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_SL g4591 ( 
.A(n_2894),
.B(n_2893),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_3303),
.Y(n_4592)
);

AOI22xp5_ASAP7_75t_L g4593 ( 
.A1(n_3318),
.A2(n_3149),
.B1(n_3167),
.B2(n_3164),
.Y(n_4593)
);

NAND2xp5_ASAP7_75t_SL g4594 ( 
.A(n_3297),
.B(n_3065),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_3304),
.Y(n_4595)
);

AND2x2_ASAP7_75t_L g4596 ( 
.A(n_3366),
.B(n_3373),
.Y(n_4596)
);

AOI22xp33_ASAP7_75t_L g4597 ( 
.A1(n_3308),
.A2(n_3382),
.B1(n_3494),
.B2(n_3493),
.Y(n_4597)
);

INVxp33_ASAP7_75t_L g4598 ( 
.A(n_3466),
.Y(n_4598)
);

INVx2_ASAP7_75t_SL g4599 ( 
.A(n_3424),
.Y(n_4599)
);

INVx2_ASAP7_75t_SL g4600 ( 
.A(n_3442),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_3366),
.B(n_3373),
.Y(n_4601)
);

NOR2xp33_ASAP7_75t_L g4602 ( 
.A(n_3172),
.B(n_3271),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_SL g4603 ( 
.A(n_3297),
.B(n_3067),
.Y(n_4603)
);

INVx2_ASAP7_75t_SL g4604 ( 
.A(n_3442),
.Y(n_4604)
);

BUFx3_ASAP7_75t_L g4605 ( 
.A(n_3363),
.Y(n_4605)
);

CKINVDCx5p33_ASAP7_75t_R g4606 ( 
.A(n_3129),
.Y(n_4606)
);

HB1xp67_ASAP7_75t_L g4607 ( 
.A(n_2905),
.Y(n_4607)
);

INVx4_ASAP7_75t_L g4608 ( 
.A(n_3442),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_3304),
.Y(n_4609)
);

BUFx3_ASAP7_75t_L g4610 ( 
.A(n_3392),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_SL g4611 ( 
.A(n_3409),
.B(n_3342),
.Y(n_4611)
);

NAND3xp33_ASAP7_75t_L g4612 ( 
.A(n_3192),
.B(n_3274),
.C(n_3275),
.Y(n_4612)
);

NAND2x1p5_ASAP7_75t_L g4613 ( 
.A(n_3464),
.B(n_3030),
.Y(n_4613)
);

INVx3_ASAP7_75t_L g4614 ( 
.A(n_3442),
.Y(n_4614)
);

CKINVDCx5p33_ASAP7_75t_R g4615 ( 
.A(n_3308),
.Y(n_4615)
);

INVx3_ASAP7_75t_SL g4616 ( 
.A(n_3442),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_3314),
.Y(n_4617)
);

NAND2xp5_ASAP7_75t_L g4618 ( 
.A(n_3421),
.B(n_3459),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_L g4619 ( 
.A(n_3459),
.B(n_3437),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_3314),
.Y(n_4620)
);

NAND2xp5_ASAP7_75t_L g4621 ( 
.A(n_3437),
.B(n_3439),
.Y(n_4621)
);

INVx4_ASAP7_75t_L g4622 ( 
.A(n_3442),
.Y(n_4622)
);

NAND2xp5_ASAP7_75t_L g4623 ( 
.A(n_3439),
.B(n_3440),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_3440),
.B(n_3261),
.Y(n_4624)
);

BUFx3_ASAP7_75t_L g4625 ( 
.A(n_3392),
.Y(n_4625)
);

AOI22xp5_ASAP7_75t_L g4626 ( 
.A1(n_3214),
.A2(n_3257),
.B1(n_3493),
.B2(n_3382),
.Y(n_4626)
);

CKINVDCx5p33_ASAP7_75t_R g4627 ( 
.A(n_3382),
.Y(n_4627)
);

NOR2xp33_ASAP7_75t_L g4628 ( 
.A(n_3187),
.B(n_3254),
.Y(n_4628)
);

OAI22xp5_ASAP7_75t_L g4629 ( 
.A1(n_3469),
.A2(n_2975),
.B1(n_2963),
.B2(n_3409),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_3331),
.B(n_3334),
.Y(n_4630)
);

INVxp67_ASAP7_75t_SL g4631 ( 
.A(n_3324),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_SL g4632 ( 
.A(n_3342),
.B(n_3475),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_3324),
.Y(n_4633)
);

NOR2xp33_ASAP7_75t_R g4634 ( 
.A(n_2963),
.B(n_2975),
.Y(n_4634)
);

AOI22xp33_ASAP7_75t_L g4635 ( 
.A1(n_3230),
.A2(n_3474),
.B1(n_3452),
.B2(n_3370),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_SL g4636 ( 
.A(n_3475),
.B(n_3335),
.Y(n_4636)
);

INVx4_ASAP7_75t_L g4637 ( 
.A(n_3460),
.Y(n_4637)
);

NOR2xp33_ASAP7_75t_L g4638 ( 
.A(n_3472),
.B(n_3255),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_3340),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_3331),
.B(n_3334),
.Y(n_4640)
);

AOI22xp5_ASAP7_75t_L g4641 ( 
.A1(n_3369),
.A2(n_3370),
.B1(n_3450),
.B2(n_3020),
.Y(n_4641)
);

NAND2xp5_ASAP7_75t_L g4642 ( 
.A(n_3338),
.B(n_3395),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_3340),
.Y(n_4643)
);

BUFx4f_ASAP7_75t_L g4644 ( 
.A(n_3020),
.Y(n_4644)
);

HB1xp67_ASAP7_75t_L g4645 ( 
.A(n_2881),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_3338),
.B(n_3395),
.Y(n_4646)
);

NAND2xp5_ASAP7_75t_L g4647 ( 
.A(n_3400),
.B(n_3369),
.Y(n_4647)
);

A2O1A1Ixp33_ASAP7_75t_L g4648 ( 
.A1(n_3339),
.A2(n_3288),
.B(n_3156),
.C(n_3361),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_3341),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_3400),
.B(n_3451),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_3419),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_3341),
.Y(n_4652)
);

NAND2xp5_ASAP7_75t_L g4653 ( 
.A(n_3451),
.B(n_3030),
.Y(n_4653)
);

HB1xp67_ASAP7_75t_L g4654 ( 
.A(n_2881),
.Y(n_4654)
);

INVx2_ASAP7_75t_SL g4655 ( 
.A(n_3460),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_L g4656 ( 
.A(n_3328),
.B(n_3377),
.Y(n_4656)
);

BUFx4f_ASAP7_75t_L g4657 ( 
.A(n_3020),
.Y(n_4657)
);

BUFx3_ASAP7_75t_L g4658 ( 
.A(n_3402),
.Y(n_4658)
);

AND2x2_ASAP7_75t_L g4659 ( 
.A(n_3377),
.B(n_3387),
.Y(n_4659)
);

BUFx2_ASAP7_75t_SL g4660 ( 
.A(n_3460),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_3387),
.B(n_3603),
.Y(n_4661)
);

AOI22xp5_ASAP7_75t_L g4662 ( 
.A1(n_3450),
.A2(n_3780),
.B1(n_3020),
.B2(n_3230),
.Y(n_4662)
);

AND2x4_ASAP7_75t_L g4663 ( 
.A(n_3381),
.B(n_3384),
.Y(n_4663)
);

AOI22xp33_ASAP7_75t_L g4664 ( 
.A1(n_3452),
.A2(n_3474),
.B1(n_3360),
.B2(n_3020),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_SL g4665 ( 
.A(n_3391),
.B(n_3336),
.Y(n_4665)
);

OR2x2_ASAP7_75t_L g4666 ( 
.A(n_3329),
.B(n_3603),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_3419),
.Y(n_4667)
);

AOI22xp33_ASAP7_75t_L g4668 ( 
.A1(n_3360),
.A2(n_3780),
.B1(n_3467),
.B2(n_2975),
.Y(n_4668)
);

NAND2xp5_ASAP7_75t_L g4669 ( 
.A(n_3328),
.B(n_3352),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_3352),
.B(n_3460),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_3614),
.Y(n_4671)
);

INVx5_ASAP7_75t_L g4672 ( 
.A(n_3780),
.Y(n_4672)
);

OAI22xp33_ASAP7_75t_L g4673 ( 
.A1(n_2963),
.A2(n_2975),
.B1(n_3138),
.B2(n_3108),
.Y(n_4673)
);

OAI22xp5_ASAP7_75t_L g4674 ( 
.A1(n_3469),
.A2(n_3301),
.B1(n_3484),
.B2(n_3473),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_3619),
.Y(n_4675)
);

AOI21xp5_ASAP7_75t_L g4676 ( 
.A1(n_4165),
.A2(n_3356),
.B(n_3346),
.Y(n_4676)
);

OA21x2_ASAP7_75t_L g4677 ( 
.A1(n_4137),
.A2(n_3201),
.B(n_3200),
.Y(n_4677)
);

AND2x4_ASAP7_75t_L g4678 ( 
.A(n_4133),
.B(n_3381),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4071),
.Y(n_4679)
);

AOI22xp33_ASAP7_75t_L g4680 ( 
.A1(n_4135),
.A2(n_3360),
.B1(n_3780),
.B2(n_3476),
.Y(n_4680)
);

INVx3_ASAP7_75t_L g4681 ( 
.A(n_3842),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4071),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_4077),
.Y(n_4683)
);

BUFx2_ASAP7_75t_L g4684 ( 
.A(n_4244),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4077),
.Y(n_4685)
);

BUFx3_ASAP7_75t_L g4686 ( 
.A(n_4229),
.Y(n_4686)
);

HB1xp67_ASAP7_75t_L g4687 ( 
.A(n_3888),
.Y(n_4687)
);

CKINVDCx6p67_ASAP7_75t_R g4688 ( 
.A(n_4229),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4078),
.Y(n_4689)
);

INVx2_ASAP7_75t_L g4690 ( 
.A(n_3997),
.Y(n_4690)
);

INVxp67_ASAP7_75t_SL g4691 ( 
.A(n_4186),
.Y(n_4691)
);

BUFx6f_ASAP7_75t_L g4692 ( 
.A(n_3883),
.Y(n_4692)
);

NOR2xp33_ASAP7_75t_L g4693 ( 
.A(n_3877),
.B(n_3466),
.Y(n_4693)
);

NOR2xp33_ASAP7_75t_L g4694 ( 
.A(n_3877),
.B(n_3466),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4078),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_4010),
.B(n_3337),
.Y(n_4696)
);

NOR2xp33_ASAP7_75t_L g4697 ( 
.A(n_3912),
.B(n_3466),
.Y(n_4697)
);

INVx3_ASAP7_75t_L g4698 ( 
.A(n_3842),
.Y(n_4698)
);

O2A1O1Ixp33_ASAP7_75t_L g4699 ( 
.A1(n_4305),
.A2(n_3483),
.B(n_3470),
.C(n_3468),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_SL g4700 ( 
.A(n_4043),
.B(n_3315),
.Y(n_4700)
);

NOR2xp33_ASAP7_75t_L g4701 ( 
.A(n_3912),
.B(n_3466),
.Y(n_4701)
);

AND2x2_ASAP7_75t_L g4702 ( 
.A(n_4167),
.B(n_3619),
.Y(n_4702)
);

HB1xp67_ASAP7_75t_L g4703 ( 
.A(n_3888),
.Y(n_4703)
);

INVx3_ASAP7_75t_L g4704 ( 
.A(n_3842),
.Y(n_4704)
);

AOI21xp5_ASAP7_75t_L g4705 ( 
.A1(n_4165),
.A2(n_3457),
.B(n_3413),
.Y(n_4705)
);

AOI21xp5_ASAP7_75t_L g4706 ( 
.A1(n_4493),
.A2(n_3458),
.B(n_3386),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4105),
.Y(n_4707)
);

INVx6_ASAP7_75t_L g4708 ( 
.A(n_4002),
.Y(n_4708)
);

A2O1A1Ixp33_ASAP7_75t_L g4709 ( 
.A1(n_4124),
.A2(n_3127),
.B(n_3136),
.C(n_3123),
.Y(n_4709)
);

INVx1_ASAP7_75t_SL g4710 ( 
.A(n_3895),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4010),
.B(n_3337),
.Y(n_4711)
);

A2O1A1Ixp33_ASAP7_75t_SL g4712 ( 
.A1(n_4412),
.A2(n_4483),
.B(n_4317),
.C(n_4330),
.Y(n_4712)
);

AOI21xp5_ASAP7_75t_L g4713 ( 
.A1(n_4493),
.A2(n_3397),
.B(n_3383),
.Y(n_4713)
);

INVx2_ASAP7_75t_SL g4714 ( 
.A(n_4320),
.Y(n_4714)
);

AOI22xp5_ASAP7_75t_L g4715 ( 
.A1(n_4014),
.A2(n_3360),
.B1(n_3780),
.B2(n_3418),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_3997),
.Y(n_4716)
);

AND2x4_ASAP7_75t_L g4717 ( 
.A(n_4133),
.B(n_3384),
.Y(n_4717)
);

INVx2_ASAP7_75t_L g4718 ( 
.A(n_3997),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4105),
.Y(n_4719)
);

AND2x2_ASAP7_75t_L g4720 ( 
.A(n_4167),
.B(n_3619),
.Y(n_4720)
);

INVx5_ASAP7_75t_L g4721 ( 
.A(n_3883),
.Y(n_4721)
);

OAI22xp5_ASAP7_75t_L g4722 ( 
.A1(n_3999),
.A2(n_3469),
.B1(n_3108),
.B2(n_3138),
.Y(n_4722)
);

INVx2_ASAP7_75t_SL g4723 ( 
.A(n_4320),
.Y(n_4723)
);

BUFx3_ASAP7_75t_L g4724 ( 
.A(n_4229),
.Y(n_4724)
);

AND2x2_ASAP7_75t_L g4725 ( 
.A(n_4167),
.B(n_3625),
.Y(n_4725)
);

INVx2_ASAP7_75t_L g4726 ( 
.A(n_3997),
.Y(n_4726)
);

AOI22xp5_ASAP7_75t_L g4727 ( 
.A1(n_4014),
.A2(n_3360),
.B1(n_3418),
.B2(n_3491),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4113),
.Y(n_4728)
);

O2A1O1Ixp5_ASAP7_75t_SL g4729 ( 
.A1(n_4083),
.A2(n_4091),
.B(n_4219),
.C(n_4479),
.Y(n_4729)
);

CKINVDCx5p33_ASAP7_75t_R g4730 ( 
.A(n_4132),
.Y(n_4730)
);

BUFx2_ASAP7_75t_L g4731 ( 
.A(n_4244),
.Y(n_4731)
);

NOR2xp33_ASAP7_75t_L g4732 ( 
.A(n_3930),
.B(n_3967),
.Y(n_4732)
);

NAND3xp33_ASAP7_75t_L g4733 ( 
.A(n_4305),
.B(n_3376),
.C(n_3365),
.Y(n_4733)
);

O2A1O1Ixp5_ASAP7_75t_L g4734 ( 
.A1(n_3863),
.A2(n_3463),
.B(n_3477),
.C(n_3232),
.Y(n_4734)
);

NAND3xp33_ASAP7_75t_L g4735 ( 
.A(n_4482),
.B(n_3376),
.C(n_3488),
.Y(n_4735)
);

INVx2_ASAP7_75t_SL g4736 ( 
.A(n_4320),
.Y(n_4736)
);

O2A1O1Ixp33_ASAP7_75t_L g4737 ( 
.A1(n_4482),
.A2(n_3426),
.B(n_3405),
.C(n_3316),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4113),
.Y(n_4738)
);

INVx4_ASAP7_75t_L g4739 ( 
.A(n_4432),
.Y(n_4739)
);

AND2x4_ASAP7_75t_L g4740 ( 
.A(n_4133),
.B(n_3463),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_SL g4741 ( 
.A(n_4043),
.B(n_3349),
.Y(n_4741)
);

AOI21xp5_ASAP7_75t_L g4742 ( 
.A1(n_4518),
.A2(n_3401),
.B(n_3399),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4131),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_SL g4744 ( 
.A(n_3930),
.B(n_3349),
.Y(n_4744)
);

BUFx6f_ASAP7_75t_L g4745 ( 
.A(n_3883),
.Y(n_4745)
);

OAI21x1_ASAP7_75t_L g4746 ( 
.A1(n_4048),
.A2(n_4277),
.B(n_4177),
.Y(n_4746)
);

INVx2_ASAP7_75t_L g4747 ( 
.A(n_4007),
.Y(n_4747)
);

AOI22xp5_ASAP7_75t_L g4748 ( 
.A1(n_4070),
.A2(n_3360),
.B1(n_3454),
.B2(n_3431),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4131),
.Y(n_4749)
);

O2A1O1Ixp5_ASAP7_75t_SL g4750 ( 
.A1(n_4083),
.A2(n_3182),
.B(n_3184),
.C(n_3179),
.Y(n_4750)
);

CKINVDCx5p33_ASAP7_75t_R g4751 ( 
.A(n_4132),
.Y(n_4751)
);

NOR2xp33_ASAP7_75t_L g4752 ( 
.A(n_3967),
.B(n_3466),
.Y(n_4752)
);

CKINVDCx20_ASAP7_75t_R g4753 ( 
.A(n_3850),
.Y(n_4753)
);

BUFx12f_ASAP7_75t_L g4754 ( 
.A(n_3925),
.Y(n_4754)
);

NOR2xp33_ASAP7_75t_L g4755 ( 
.A(n_4025),
.B(n_3375),
.Y(n_4755)
);

AND2x2_ASAP7_75t_L g4756 ( 
.A(n_4187),
.B(n_3625),
.Y(n_4756)
);

BUFx3_ASAP7_75t_L g4757 ( 
.A(n_4229),
.Y(n_4757)
);

AOI22xp5_ASAP7_75t_L g4758 ( 
.A1(n_4070),
.A2(n_3360),
.B1(n_3454),
.B2(n_3108),
.Y(n_4758)
);

INVx2_ASAP7_75t_L g4759 ( 
.A(n_4007),
.Y(n_4759)
);

INVxp67_ASAP7_75t_SL g4760 ( 
.A(n_4186),
.Y(n_4760)
);

INVx3_ASAP7_75t_L g4761 ( 
.A(n_3842),
.Y(n_4761)
);

NOR2x1_ASAP7_75t_L g4762 ( 
.A(n_4227),
.B(n_3134),
.Y(n_4762)
);

O2A1O1Ixp33_ASAP7_75t_L g4763 ( 
.A1(n_4545),
.A2(n_3305),
.B(n_3446),
.C(n_3433),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4484),
.Y(n_4764)
);

NOR2xp67_ASAP7_75t_SL g4765 ( 
.A(n_3913),
.B(n_3891),
.Y(n_4765)
);

INVx3_ASAP7_75t_L g4766 ( 
.A(n_3842),
.Y(n_4766)
);

AND2x2_ASAP7_75t_L g4767 ( 
.A(n_4187),
.B(n_3625),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4007),
.Y(n_4768)
);

O2A1O1Ixp5_ASAP7_75t_L g4769 ( 
.A1(n_3863),
.A2(n_3438),
.B(n_3429),
.C(n_3445),
.Y(n_4769)
);

HB1xp67_ASAP7_75t_L g4770 ( 
.A(n_3918),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4484),
.Y(n_4771)
);

AND3x1_ASAP7_75t_SL g4772 ( 
.A(n_3891),
.B(n_3469),
.C(n_3461),
.Y(n_4772)
);

A2O1A1Ixp33_ASAP7_75t_L g4773 ( 
.A1(n_4124),
.A2(n_3122),
.B(n_3296),
.C(n_3263),
.Y(n_4773)
);

AOI22xp5_ASAP7_75t_L g4774 ( 
.A1(n_4135),
.A2(n_3360),
.B1(n_3454),
.B2(n_3108),
.Y(n_4774)
);

OR2x6_ASAP7_75t_L g4775 ( 
.A(n_4090),
.B(n_3216),
.Y(n_4775)
);

AOI22xp33_ASAP7_75t_L g4776 ( 
.A1(n_3871),
.A2(n_3476),
.B1(n_3216),
.B2(n_3138),
.Y(n_4776)
);

NAND2xp5_ASAP7_75t_L g4777 ( 
.A(n_4024),
.B(n_3134),
.Y(n_4777)
);

AOI22xp5_ASAP7_75t_L g4778 ( 
.A1(n_4246),
.A2(n_3454),
.B1(n_3138),
.B2(n_3453),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4490),
.Y(n_4779)
);

O2A1O1Ixp33_ASAP7_75t_L g4780 ( 
.A1(n_4545),
.A2(n_3336),
.B(n_3490),
.C(n_3486),
.Y(n_4780)
);

INVx3_ASAP7_75t_SL g4781 ( 
.A(n_4611),
.Y(n_4781)
);

BUFx3_ASAP7_75t_L g4782 ( 
.A(n_4363),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4490),
.Y(n_4783)
);

CKINVDCx14_ASAP7_75t_R g4784 ( 
.A(n_3847),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_3851),
.Y(n_4785)
);

AND2x2_ASAP7_75t_L g4786 ( 
.A(n_4187),
.B(n_3641),
.Y(n_4786)
);

INVx4_ASAP7_75t_L g4787 ( 
.A(n_4432),
.Y(n_4787)
);

BUFx6f_ASAP7_75t_L g4788 ( 
.A(n_3883),
.Y(n_4788)
);

OR2x6_ASAP7_75t_L g4789 ( 
.A(n_4090),
.B(n_3216),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_3851),
.Y(n_4790)
);

A2O1A1Ixp33_ASAP7_75t_L g4791 ( 
.A1(n_4494),
.A2(n_3263),
.B(n_3296),
.C(n_3253),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_SL g4792 ( 
.A(n_4025),
.B(n_3349),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_3851),
.Y(n_4793)
);

AOI21xp5_ASAP7_75t_L g4794 ( 
.A1(n_4518),
.A2(n_4250),
.B(n_4230),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_L g4795 ( 
.A(n_4024),
.B(n_3134),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_3852),
.Y(n_4796)
);

BUFx6f_ASAP7_75t_L g4797 ( 
.A(n_3883),
.Y(n_4797)
);

AND2x2_ASAP7_75t_L g4798 ( 
.A(n_4271),
.B(n_3641),
.Y(n_4798)
);

INVx2_ASAP7_75t_L g4799 ( 
.A(n_4007),
.Y(n_4799)
);

AOI21xp5_ASAP7_75t_SL g4800 ( 
.A1(n_4073),
.A2(n_3414),
.B(n_3449),
.Y(n_4800)
);

AND2x2_ASAP7_75t_L g4801 ( 
.A(n_4271),
.B(n_3641),
.Y(n_4801)
);

O2A1O1Ixp33_ASAP7_75t_L g4802 ( 
.A1(n_4301),
.A2(n_3441),
.B(n_3348),
.C(n_3479),
.Y(n_4802)
);

NOR2xp33_ASAP7_75t_L g4803 ( 
.A(n_4036),
.B(n_3388),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_3852),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_3852),
.Y(n_4805)
);

BUFx2_ASAP7_75t_L g4806 ( 
.A(n_4276),
.Y(n_4806)
);

OA21x2_ASAP7_75t_L g4807 ( 
.A1(n_4137),
.A2(n_3295),
.B(n_3262),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_SL g4808 ( 
.A(n_4036),
.B(n_3349),
.Y(n_4808)
);

AOI22xp33_ASAP7_75t_L g4809 ( 
.A1(n_3871),
.A2(n_3216),
.B1(n_3456),
.B2(n_3453),
.Y(n_4809)
);

BUFx2_ASAP7_75t_L g4810 ( 
.A(n_4276),
.Y(n_4810)
);

INVxp67_ASAP7_75t_L g4811 ( 
.A(n_4034),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_SL g4812 ( 
.A(n_3832),
.B(n_3349),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_SL g4813 ( 
.A(n_3832),
.B(n_3349),
.Y(n_4813)
);

AOI22xp5_ASAP7_75t_L g4814 ( 
.A1(n_4246),
.A2(n_3908),
.B1(n_4054),
.B2(n_4040),
.Y(n_4814)
);

OAI21xp33_ASAP7_75t_L g4815 ( 
.A1(n_4300),
.A2(n_3393),
.B(n_3432),
.Y(n_4815)
);

NOR2xp33_ASAP7_75t_L g4816 ( 
.A(n_4300),
.B(n_3434),
.Y(n_4816)
);

BUFx6f_ASAP7_75t_L g4817 ( 
.A(n_3883),
.Y(n_4817)
);

BUFx12f_ASAP7_75t_L g4818 ( 
.A(n_3925),
.Y(n_4818)
);

NOR2xp33_ASAP7_75t_L g4819 ( 
.A(n_4317),
.B(n_3462),
.Y(n_4819)
);

HB1xp67_ASAP7_75t_L g4820 ( 
.A(n_3918),
.Y(n_4820)
);

NAND2xp5_ASAP7_75t_SL g4821 ( 
.A(n_3975),
.B(n_3350),
.Y(n_4821)
);

HB1xp67_ASAP7_75t_L g4822 ( 
.A(n_4034),
.Y(n_4822)
);

AOI21xp5_ASAP7_75t_L g4823 ( 
.A1(n_4230),
.A2(n_3411),
.B(n_3403),
.Y(n_4823)
);

AOI21xp5_ASAP7_75t_L g4824 ( 
.A1(n_4250),
.A2(n_3404),
.B(n_3407),
.Y(n_4824)
);

NAND2x1p5_ASAP7_75t_L g4825 ( 
.A(n_4672),
.B(n_3840),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_SL g4826 ( 
.A(n_3975),
.B(n_3350),
.Y(n_4826)
);

AOI22xp33_ASAP7_75t_L g4827 ( 
.A1(n_4040),
.A2(n_3216),
.B1(n_3456),
.B2(n_3402),
.Y(n_4827)
);

BUFx2_ASAP7_75t_L g4828 ( 
.A(n_4286),
.Y(n_4828)
);

BUFx6f_ASAP7_75t_L g4829 ( 
.A(n_3883),
.Y(n_4829)
);

NAND2xp5_ASAP7_75t_L g4830 ( 
.A(n_4108),
.B(n_3179),
.Y(n_4830)
);

OAI22xp5_ASAP7_75t_L g4831 ( 
.A1(n_3999),
.A2(n_3471),
.B1(n_3296),
.B2(n_3263),
.Y(n_4831)
);

BUFx6f_ASAP7_75t_L g4832 ( 
.A(n_3905),
.Y(n_4832)
);

AOI22xp33_ASAP7_75t_L g4833 ( 
.A1(n_4054),
.A2(n_3471),
.B1(n_3447),
.B2(n_3423),
.Y(n_4833)
);

INVx3_ASAP7_75t_L g4834 ( 
.A(n_3842),
.Y(n_4834)
);

BUFx3_ASAP7_75t_L g4835 ( 
.A(n_4363),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_3853),
.Y(n_4836)
);

AOI21xp5_ASAP7_75t_L g4837 ( 
.A1(n_4275),
.A2(n_3364),
.B(n_3354),
.Y(n_4837)
);

AOI21xp5_ASAP7_75t_L g4838 ( 
.A1(n_4275),
.A2(n_3353),
.B(n_3347),
.Y(n_4838)
);

INVxp33_ASAP7_75t_L g4839 ( 
.A(n_4638),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_L g4840 ( 
.A(n_4108),
.B(n_3184),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_4110),
.B(n_3184),
.Y(n_4841)
);

BUFx3_ASAP7_75t_L g4842 ( 
.A(n_4363),
.Y(n_4842)
);

AOI22xp33_ASAP7_75t_L g4843 ( 
.A1(n_3936),
.A2(n_3471),
.B1(n_3447),
.B2(n_3443),
.Y(n_4843)
);

OAI21xp5_ASAP7_75t_L g4844 ( 
.A1(n_4008),
.A2(n_3374),
.B(n_3430),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4110),
.B(n_3184),
.Y(n_4845)
);

HB1xp67_ASAP7_75t_L g4846 ( 
.A(n_4111),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_3853),
.Y(n_4847)
);

NAND2xp5_ASAP7_75t_L g4848 ( 
.A(n_4111),
.B(n_3018),
.Y(n_4848)
);

AND2x2_ASAP7_75t_L g4849 ( 
.A(n_4271),
.B(n_3679),
.Y(n_4849)
);

INVx5_ASAP7_75t_L g4850 ( 
.A(n_3905),
.Y(n_4850)
);

OR2x6_ASAP7_75t_L g4851 ( 
.A(n_4090),
.B(n_3220),
.Y(n_4851)
);

CKINVDCx16_ASAP7_75t_R g4852 ( 
.A(n_4196),
.Y(n_4852)
);

BUFx8_ASAP7_75t_L g4853 ( 
.A(n_4363),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_3853),
.Y(n_4854)
);

OR2x6_ASAP7_75t_L g4855 ( 
.A(n_4090),
.B(n_3220),
.Y(n_4855)
);

NAND2x1_ASAP7_75t_L g4856 ( 
.A(n_3840),
.B(n_3190),
.Y(n_4856)
);

BUFx2_ASAP7_75t_L g4857 ( 
.A(n_4286),
.Y(n_4857)
);

NOR2xp33_ASAP7_75t_L g4858 ( 
.A(n_4330),
.B(n_3482),
.Y(n_4858)
);

INVx2_ASAP7_75t_SL g4859 ( 
.A(n_4320),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_3859),
.Y(n_4860)
);

AOI21xp5_ASAP7_75t_L g4861 ( 
.A1(n_4280),
.A2(n_3253),
.B(n_3343),
.Y(n_4861)
);

NAND2x1p5_ASAP7_75t_L g4862 ( 
.A(n_4672),
.B(n_3263),
.Y(n_4862)
);

A2O1A1Ixp33_ASAP7_75t_L g4863 ( 
.A1(n_4494),
.A2(n_3296),
.B(n_3343),
.C(n_3209),
.Y(n_4863)
);

AOI21xp5_ASAP7_75t_L g4864 ( 
.A1(n_4280),
.A2(n_3209),
.B(n_3465),
.Y(n_4864)
);

AND2x4_ASAP7_75t_L g4865 ( 
.A(n_4178),
.B(n_3333),
.Y(n_4865)
);

CKINVDCx20_ASAP7_75t_R g4866 ( 
.A(n_3850),
.Y(n_4866)
);

AND2x2_ASAP7_75t_L g4867 ( 
.A(n_4279),
.B(n_4291),
.Y(n_4867)
);

HB1xp67_ASAP7_75t_L g4868 ( 
.A(n_4120),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_SL g4869 ( 
.A(n_4015),
.B(n_3350),
.Y(n_4869)
);

BUFx3_ASAP7_75t_L g4870 ( 
.A(n_4347),
.Y(n_4870)
);

O2A1O1Ixp33_ASAP7_75t_L g4871 ( 
.A1(n_4301),
.A2(n_4483),
.B(n_4412),
.C(n_4390),
.Y(n_4871)
);

INVx2_ASAP7_75t_SL g4872 ( 
.A(n_4320),
.Y(n_4872)
);

AOI21xp5_ASAP7_75t_L g4873 ( 
.A1(n_4273),
.A2(n_3441),
.B(n_3420),
.Y(n_4873)
);

AND2x2_ASAP7_75t_L g4874 ( 
.A(n_4279),
.B(n_3679),
.Y(n_4874)
);

O2A1O1Ixp33_ASAP7_75t_L g4875 ( 
.A1(n_4390),
.A2(n_3348),
.B(n_3485),
.C(n_3478),
.Y(n_4875)
);

AOI21xp5_ASAP7_75t_L g4876 ( 
.A1(n_4273),
.A2(n_3416),
.B(n_3350),
.Y(n_4876)
);

NAND2xp5_ASAP7_75t_L g4877 ( 
.A(n_4120),
.B(n_3018),
.Y(n_4877)
);

O2A1O1Ixp33_ASAP7_75t_L g4878 ( 
.A1(n_4008),
.A2(n_3471),
.B(n_3224),
.C(n_3213),
.Y(n_4878)
);

HB1xp67_ASAP7_75t_L g4879 ( 
.A(n_4148),
.Y(n_4879)
);

BUFx2_ASAP7_75t_L g4880 ( 
.A(n_4288),
.Y(n_4880)
);

BUFx2_ASAP7_75t_SL g4881 ( 
.A(n_3895),
.Y(n_4881)
);

OAI22xp5_ASAP7_75t_SL g4882 ( 
.A1(n_4338),
.A2(n_3236),
.B1(n_3220),
.B2(n_3415),
.Y(n_4882)
);

INVxp67_ASAP7_75t_SL g4883 ( 
.A(n_4203),
.Y(n_4883)
);

HB1xp67_ASAP7_75t_L g4884 ( 
.A(n_4148),
.Y(n_4884)
);

INVx2_ASAP7_75t_SL g4885 ( 
.A(n_4320),
.Y(n_4885)
);

NAND2xp5_ASAP7_75t_L g4886 ( 
.A(n_4163),
.B(n_3019),
.Y(n_4886)
);

NOR2xp33_ASAP7_75t_SL g4887 ( 
.A(n_4022),
.B(n_3427),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_L g4888 ( 
.A(n_4163),
.B(n_3019),
.Y(n_4888)
);

CKINVDCx11_ASAP7_75t_R g4889 ( 
.A(n_3910),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_3859),
.Y(n_4890)
);

INVx2_ASAP7_75t_SL g4891 ( 
.A(n_4320),
.Y(n_4891)
);

NAND2xp5_ASAP7_75t_L g4892 ( 
.A(n_4164),
.B(n_3034),
.Y(n_4892)
);

NOR2xp33_ASAP7_75t_L g4893 ( 
.A(n_4338),
.B(n_3190),
.Y(n_4893)
);

CKINVDCx5p33_ASAP7_75t_R g4894 ( 
.A(n_4013),
.Y(n_4894)
);

A2O1A1Ixp33_ASAP7_75t_L g4895 ( 
.A1(n_4212),
.A2(n_3427),
.B(n_3443),
.C(n_3428),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_3859),
.Y(n_4896)
);

NOR2xp33_ASAP7_75t_L g4897 ( 
.A(n_4181),
.B(n_3190),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_3874),
.Y(n_4898)
);

INVx4_ASAP7_75t_L g4899 ( 
.A(n_4432),
.Y(n_4899)
);

CKINVDCx14_ASAP7_75t_R g4900 ( 
.A(n_3847),
.Y(n_4900)
);

INVx2_ASAP7_75t_SL g4901 ( 
.A(n_4320),
.Y(n_4901)
);

BUFx2_ASAP7_75t_L g4902 ( 
.A(n_4288),
.Y(n_4902)
);

NOR2xp67_ASAP7_75t_L g4903 ( 
.A(n_4324),
.B(n_3190),
.Y(n_4903)
);

AOI21xp5_ASAP7_75t_L g4904 ( 
.A1(n_4298),
.A2(n_3398),
.B(n_3350),
.Y(n_4904)
);

NOR2xp33_ASAP7_75t_L g4905 ( 
.A(n_4181),
.B(n_3195),
.Y(n_4905)
);

AND2x2_ASAP7_75t_L g4906 ( 
.A(n_4279),
.B(n_3679),
.Y(n_4906)
);

OAI22xp5_ASAP7_75t_L g4907 ( 
.A1(n_4015),
.A2(n_3213),
.B1(n_3224),
.B2(n_3195),
.Y(n_4907)
);

NOR2xp33_ASAP7_75t_L g4908 ( 
.A(n_4287),
.B(n_3195),
.Y(n_4908)
);

INVx1_ASAP7_75t_L g4909 ( 
.A(n_3874),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_3874),
.Y(n_4910)
);

INVxp67_ASAP7_75t_L g4911 ( 
.A(n_4164),
.Y(n_4911)
);

AOI222xp33_ASAP7_75t_L g4912 ( 
.A1(n_4032),
.A2(n_3461),
.B1(n_3417),
.B2(n_3425),
.C1(n_3371),
.C2(n_3333),
.Y(n_4912)
);

INVx3_ASAP7_75t_L g4913 ( 
.A(n_3858),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_L g4914 ( 
.A(n_3868),
.B(n_3887),
.Y(n_4914)
);

NOR2xp33_ASAP7_75t_L g4915 ( 
.A(n_4287),
.B(n_3195),
.Y(n_4915)
);

O2A1O1Ixp33_ASAP7_75t_L g4916 ( 
.A1(n_4028),
.A2(n_3213),
.B(n_3224),
.C(n_3208),
.Y(n_4916)
);

CKINVDCx5p33_ASAP7_75t_R g4917 ( 
.A(n_4013),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_3876),
.Y(n_4918)
);

NOR2xp33_ASAP7_75t_SL g4919 ( 
.A(n_4022),
.B(n_3394),
.Y(n_4919)
);

NOR2xp33_ASAP7_75t_L g4920 ( 
.A(n_4427),
.B(n_3213),
.Y(n_4920)
);

NOR2xp67_ASAP7_75t_SL g4921 ( 
.A(n_3913),
.B(n_3367),
.Y(n_4921)
);

AND2x2_ASAP7_75t_L g4922 ( 
.A(n_4291),
.B(n_3790),
.Y(n_4922)
);

INVx8_ASAP7_75t_L g4923 ( 
.A(n_4052),
.Y(n_4923)
);

A2O1A1Ixp33_ASAP7_75t_SL g4924 ( 
.A1(n_4544),
.A2(n_4456),
.B(n_4269),
.C(n_4564),
.Y(n_4924)
);

XOR2xp5_ASAP7_75t_L g4925 ( 
.A(n_3910),
.B(n_4142),
.Y(n_4925)
);

AOI22xp33_ASAP7_75t_L g4926 ( 
.A1(n_3936),
.A2(n_3236),
.B1(n_3220),
.B2(n_3415),
.Y(n_4926)
);

BUFx12f_ASAP7_75t_L g4927 ( 
.A(n_3931),
.Y(n_4927)
);

BUFx3_ASAP7_75t_L g4928 ( 
.A(n_4347),
.Y(n_4928)
);

AOI22xp33_ASAP7_75t_L g4929 ( 
.A1(n_3979),
.A2(n_3236),
.B1(n_3415),
.B2(n_3394),
.Y(n_4929)
);

HB1xp67_ASAP7_75t_L g4930 ( 
.A(n_3833),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_3876),
.Y(n_4931)
);

INVx1_ASAP7_75t_L g4932 ( 
.A(n_3876),
.Y(n_4932)
);

AOI21xp5_ASAP7_75t_L g4933 ( 
.A1(n_4298),
.A2(n_3398),
.B(n_3367),
.Y(n_4933)
);

OAI22xp5_ASAP7_75t_L g4934 ( 
.A1(n_4027),
.A2(n_3224),
.B1(n_3034),
.B2(n_3516),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_3878),
.Y(n_4935)
);

INVx1_ASAP7_75t_SL g4936 ( 
.A(n_3909),
.Y(n_4936)
);

OAI221xp5_ASAP7_75t_L g4937 ( 
.A1(n_3979),
.A2(n_3422),
.B1(n_3417),
.B2(n_3425),
.C(n_3236),
.Y(n_4937)
);

INVx3_ASAP7_75t_L g4938 ( 
.A(n_3858),
.Y(n_4938)
);

AOI22xp33_ASAP7_75t_L g4939 ( 
.A1(n_4032),
.A2(n_3415),
.B1(n_3750),
.B2(n_3743),
.Y(n_4939)
);

CKINVDCx20_ASAP7_75t_R g4940 ( 
.A(n_4142),
.Y(n_4940)
);

AOI21x1_ASAP7_75t_L g4941 ( 
.A1(n_4223),
.A2(n_3444),
.B(n_3455),
.Y(n_4941)
);

OAI22xp5_ASAP7_75t_SL g4942 ( 
.A1(n_4354),
.A2(n_4427),
.B1(n_4212),
.B2(n_4235),
.Y(n_4942)
);

INVx1_ASAP7_75t_L g4943 ( 
.A(n_3878),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_3878),
.Y(n_4944)
);

OR2x2_ASAP7_75t_L g4945 ( 
.A(n_4006),
.B(n_3790),
.Y(n_4945)
);

A2O1A1Ixp33_ASAP7_75t_SL g4946 ( 
.A1(n_4544),
.A2(n_3516),
.B(n_3661),
.C(n_3721),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_3884),
.Y(n_4947)
);

A2O1A1Ixp33_ASAP7_75t_L g4948 ( 
.A1(n_4235),
.A2(n_3371),
.B(n_3333),
.C(n_3222),
.Y(n_4948)
);

AOI21xp5_ASAP7_75t_L g4949 ( 
.A1(n_4223),
.A2(n_3367),
.B(n_3398),
.Y(n_4949)
);

AOI21xp5_ASAP7_75t_L g4950 ( 
.A1(n_4281),
.A2(n_3367),
.B(n_3398),
.Y(n_4950)
);

A2O1A1Ixp33_ASAP7_75t_L g4951 ( 
.A1(n_4073),
.A2(n_3371),
.B(n_3222),
.C(n_3270),
.Y(n_4951)
);

CKINVDCx14_ASAP7_75t_R g4952 ( 
.A(n_3847),
.Y(n_4952)
);

AOI22xp5_ASAP7_75t_L g4953 ( 
.A1(n_3908),
.A2(n_3415),
.B1(n_3371),
.B2(n_3372),
.Y(n_4953)
);

BUFx2_ASAP7_75t_L g4954 ( 
.A(n_4322),
.Y(n_4954)
);

AND2x4_ASAP7_75t_SL g4955 ( 
.A(n_3840),
.B(n_3367),
.Y(n_4955)
);

INVx2_ASAP7_75t_SL g4956 ( 
.A(n_4402),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_3884),
.Y(n_4957)
);

OAI22xp5_ASAP7_75t_L g4958 ( 
.A1(n_4027),
.A2(n_3661),
.B1(n_3721),
.B2(n_3398),
.Y(n_4958)
);

BUFx5_ASAP7_75t_L g4959 ( 
.A(n_4432),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_3884),
.Y(n_4960)
);

OAI22xp5_ASAP7_75t_L g4961 ( 
.A1(n_3881),
.A2(n_3367),
.B1(n_3398),
.B2(n_3372),
.Y(n_4961)
);

HB1xp67_ASAP7_75t_L g4962 ( 
.A(n_3833),
.Y(n_4962)
);

INVx4_ASAP7_75t_L g4963 ( 
.A(n_4451),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_3893),
.Y(n_4964)
);

OAI22xp5_ASAP7_75t_L g4965 ( 
.A1(n_3881),
.A2(n_3390),
.B1(n_3208),
.B2(n_3455),
.Y(n_4965)
);

BUFx2_ASAP7_75t_L g4966 ( 
.A(n_4322),
.Y(n_4966)
);

AOI21xp5_ASAP7_75t_L g4967 ( 
.A1(n_4281),
.A2(n_3390),
.B(n_3266),
.Y(n_4967)
);

INVx3_ASAP7_75t_L g4968 ( 
.A(n_3858),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_3893),
.Y(n_4969)
);

INVx5_ASAP7_75t_L g4970 ( 
.A(n_4178),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_3893),
.Y(n_4971)
);

HB1xp67_ASAP7_75t_L g4972 ( 
.A(n_3873),
.Y(n_4972)
);

INVx1_ASAP7_75t_SL g4973 ( 
.A(n_3909),
.Y(n_4973)
);

BUFx6f_ASAP7_75t_L g4974 ( 
.A(n_3835),
.Y(n_4974)
);

INVx5_ASAP7_75t_L g4975 ( 
.A(n_4178),
.Y(n_4975)
);

AND2x2_ASAP7_75t_L g4976 ( 
.A(n_4291),
.B(n_3790),
.Y(n_4976)
);

AOI222xp33_ASAP7_75t_L g4977 ( 
.A1(n_3922),
.A2(n_3750),
.B1(n_3743),
.B2(n_3714),
.C1(n_3709),
.C2(n_3270),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_L g4978 ( 
.A(n_3868),
.B(n_3750),
.Y(n_4978)
);

NOR2xp33_ASAP7_75t_L g4979 ( 
.A(n_4564),
.B(n_3743),
.Y(n_4979)
);

NOR2xp33_ASAP7_75t_L g4980 ( 
.A(n_4354),
.B(n_3714),
.Y(n_4980)
);

BUFx12f_ASAP7_75t_L g4981 ( 
.A(n_3931),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_L g4982 ( 
.A(n_3887),
.B(n_3714),
.Y(n_4982)
);

A2O1A1Ixp33_ASAP7_75t_SL g4983 ( 
.A1(n_4456),
.A2(n_3709),
.B(n_3256),
.C(n_3200),
.Y(n_4983)
);

AOI21xp5_ASAP7_75t_L g4984 ( 
.A1(n_4559),
.A2(n_3256),
.B(n_3327),
.Y(n_4984)
);

AOI21xp5_ASAP7_75t_L g4985 ( 
.A1(n_4559),
.A2(n_4137),
.B(n_4308),
.Y(n_4985)
);

AOI21xp5_ASAP7_75t_L g4986 ( 
.A1(n_4308),
.A2(n_3262),
.B(n_3327),
.Y(n_4986)
);

BUFx6f_ASAP7_75t_L g4987 ( 
.A(n_3835),
.Y(n_4987)
);

BUFx6f_ASAP7_75t_L g4988 ( 
.A(n_3835),
.Y(n_4988)
);

NAND2x1p5_ASAP7_75t_L g4989 ( 
.A(n_4672),
.B(n_3840),
.Y(n_4989)
);

INVxp67_ASAP7_75t_L g4990 ( 
.A(n_4009),
.Y(n_4990)
);

BUFx6f_ASAP7_75t_L g4991 ( 
.A(n_3835),
.Y(n_4991)
);

OAI22xp5_ASAP7_75t_SL g4992 ( 
.A1(n_3896),
.A2(n_3709),
.B1(n_3225),
.B2(n_3215),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_3897),
.Y(n_4993)
);

AOI22xp33_ASAP7_75t_L g4994 ( 
.A1(n_4149),
.A2(n_2881),
.B1(n_3245),
.B2(n_3201),
.Y(n_4994)
);

INVx2_ASAP7_75t_L g4995 ( 
.A(n_4037),
.Y(n_4995)
);

AOI21xp33_ASAP7_75t_L g4996 ( 
.A1(n_3834),
.A2(n_2881),
.B(n_3173),
.Y(n_4996)
);

INVx2_ASAP7_75t_L g4997 ( 
.A(n_4037),
.Y(n_4997)
);

AND2x4_ASAP7_75t_L g4998 ( 
.A(n_4178),
.B(n_3173),
.Y(n_4998)
);

INVx2_ASAP7_75t_L g4999 ( 
.A(n_4037),
.Y(n_4999)
);

A2O1A1Ixp33_ASAP7_75t_L g5000 ( 
.A1(n_4628),
.A2(n_3207),
.B(n_3210),
.C(n_3211),
.Y(n_5000)
);

AOI21xp5_ASAP7_75t_L g5001 ( 
.A1(n_4310),
.A2(n_3207),
.B(n_3210),
.Y(n_5001)
);

INVx2_ASAP7_75t_L g5002 ( 
.A(n_4045),
.Y(n_5002)
);

NAND2x1p5_ASAP7_75t_L g5003 ( 
.A(n_4672),
.B(n_3225),
.Y(n_5003)
);

BUFx6f_ASAP7_75t_L g5004 ( 
.A(n_3835),
.Y(n_5004)
);

CKINVDCx5p33_ASAP7_75t_R g5005 ( 
.A(n_4161),
.Y(n_5005)
);

BUFx3_ASAP7_75t_L g5006 ( 
.A(n_4347),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4009),
.B(n_3211),
.Y(n_5007)
);

AND2x2_ASAP7_75t_L g5008 ( 
.A(n_4311),
.B(n_3215),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_L g5009 ( 
.A(n_4174),
.B(n_3227),
.Y(n_5009)
);

OR2x2_ASAP7_75t_L g5010 ( 
.A(n_4006),
.B(n_3227),
.Y(n_5010)
);

INVx2_ASAP7_75t_L g5011 ( 
.A(n_4045),
.Y(n_5011)
);

NAND2xp5_ASAP7_75t_L g5012 ( 
.A(n_4174),
.B(n_3228),
.Y(n_5012)
);

AOI21xp5_ASAP7_75t_L g5013 ( 
.A1(n_4310),
.A2(n_3228),
.B(n_3233),
.Y(n_5013)
);

AOI21xp5_ASAP7_75t_L g5014 ( 
.A1(n_4319),
.A2(n_3233),
.B(n_3238),
.Y(n_5014)
);

A2O1A1Ixp33_ASAP7_75t_SL g5015 ( 
.A1(n_4269),
.A2(n_3238),
.B(n_3239),
.C(n_3242),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_3897),
.Y(n_5016)
);

INVx3_ASAP7_75t_L g5017 ( 
.A(n_3858),
.Y(n_5017)
);

INVx1_ASAP7_75t_SL g5018 ( 
.A(n_4018),
.Y(n_5018)
);

NAND2xp5_ASAP7_75t_L g5019 ( 
.A(n_4174),
.B(n_3855),
.Y(n_5019)
);

AOI21xp5_ASAP7_75t_L g5020 ( 
.A1(n_4319),
.A2(n_3239),
.B(n_3242),
.Y(n_5020)
);

BUFx12f_ASAP7_75t_L g5021 ( 
.A(n_4447),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_3897),
.Y(n_5022)
);

A2O1A1Ixp33_ASAP7_75t_L g5023 ( 
.A1(n_4628),
.A2(n_3243),
.B(n_3245),
.C(n_3249),
.Y(n_5023)
);

AND2x4_ASAP7_75t_L g5024 ( 
.A(n_4178),
.B(n_3243),
.Y(n_5024)
);

BUFx3_ASAP7_75t_L g5025 ( 
.A(n_4610),
.Y(n_5025)
);

BUFx2_ASAP7_75t_L g5026 ( 
.A(n_4328),
.Y(n_5026)
);

INVx2_ASAP7_75t_L g5027 ( 
.A(n_4045),
.Y(n_5027)
);

BUFx2_ASAP7_75t_L g5028 ( 
.A(n_4328),
.Y(n_5028)
);

AOI21xp5_ASAP7_75t_L g5029 ( 
.A1(n_4323),
.A2(n_3249),
.B(n_3264),
.Y(n_5029)
);

AO21x2_ASAP7_75t_L g5030 ( 
.A1(n_4346),
.A2(n_3264),
.B(n_3266),
.Y(n_5030)
);

INVx2_ASAP7_75t_L g5031 ( 
.A(n_4045),
.Y(n_5031)
);

BUFx6f_ASAP7_75t_L g5032 ( 
.A(n_3835),
.Y(n_5032)
);

INVx5_ASAP7_75t_L g5033 ( 
.A(n_4178),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_L g5034 ( 
.A(n_3855),
.B(n_3268),
.Y(n_5034)
);

NOR2xp33_ASAP7_75t_R g5035 ( 
.A(n_4393),
.B(n_3268),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_3898),
.Y(n_5036)
);

OAI22xp33_ASAP7_75t_L g5037 ( 
.A1(n_4057),
.A2(n_3285),
.B1(n_3286),
.B2(n_3291),
.Y(n_5037)
);

AND2x4_ASAP7_75t_L g5038 ( 
.A(n_3948),
.B(n_3285),
.Y(n_5038)
);

AND2x4_ASAP7_75t_L g5039 ( 
.A(n_3948),
.B(n_3286),
.Y(n_5039)
);

INVx2_ASAP7_75t_L g5040 ( 
.A(n_4046),
.Y(n_5040)
);

NAND2xp5_ASAP7_75t_SL g5041 ( 
.A(n_3899),
.B(n_3291),
.Y(n_5041)
);

BUFx3_ASAP7_75t_L g5042 ( 
.A(n_4610),
.Y(n_5042)
);

CKINVDCx6p67_ASAP7_75t_R g5043 ( 
.A(n_3839),
.Y(n_5043)
);

BUFx3_ASAP7_75t_L g5044 ( 
.A(n_4610),
.Y(n_5044)
);

BUFx6f_ASAP7_75t_L g5045 ( 
.A(n_3835),
.Y(n_5045)
);

AOI21xp5_ASAP7_75t_L g5046 ( 
.A1(n_4323),
.A2(n_3295),
.B(n_3299),
.Y(n_5046)
);

INVx2_ASAP7_75t_L g5047 ( 
.A(n_4046),
.Y(n_5047)
);

NOR2xp33_ASAP7_75t_L g5048 ( 
.A(n_4194),
.B(n_3299),
.Y(n_5048)
);

NAND2x1p5_ASAP7_75t_L g5049 ( 
.A(n_4672),
.B(n_3302),
.Y(n_5049)
);

INVx2_ASAP7_75t_L g5050 ( 
.A(n_4046),
.Y(n_5050)
);

NAND2xp5_ASAP7_75t_L g5051 ( 
.A(n_3837),
.B(n_3302),
.Y(n_5051)
);

AOI21xp5_ASAP7_75t_L g5052 ( 
.A1(n_4332),
.A2(n_4371),
.B(n_4345),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_3837),
.B(n_3307),
.Y(n_5053)
);

INVx2_ASAP7_75t_L g5054 ( 
.A(n_4046),
.Y(n_5054)
);

AOI21xp5_ASAP7_75t_L g5055 ( 
.A1(n_4332),
.A2(n_3309),
.B(n_3319),
.Y(n_5055)
);

AOI21xp5_ASAP7_75t_L g5056 ( 
.A1(n_4345),
.A2(n_3309),
.B(n_3319),
.Y(n_5056)
);

AOI22xp5_ASAP7_75t_L g5057 ( 
.A1(n_4057),
.A2(n_3322),
.B1(n_3323),
.B2(n_4081),
.Y(n_5057)
);

INVx5_ASAP7_75t_L g5058 ( 
.A(n_4052),
.Y(n_5058)
);

AND2x2_ASAP7_75t_L g5059 ( 
.A(n_4311),
.B(n_3322),
.Y(n_5059)
);

BUFx6f_ASAP7_75t_L g5060 ( 
.A(n_3835),
.Y(n_5060)
);

INVx2_ASAP7_75t_L g5061 ( 
.A(n_4053),
.Y(n_5061)
);

HB1xp67_ASAP7_75t_L g5062 ( 
.A(n_3873),
.Y(n_5062)
);

BUFx2_ASAP7_75t_L g5063 ( 
.A(n_4334),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_L g5064 ( 
.A(n_3838),
.B(n_3864),
.Y(n_5064)
);

AOI21xp5_ASAP7_75t_L g5065 ( 
.A1(n_4371),
.A2(n_4431),
.B(n_4375),
.Y(n_5065)
);

INVx2_ASAP7_75t_L g5066 ( 
.A(n_4053),
.Y(n_5066)
);

NAND2xp5_ASAP7_75t_L g5067 ( 
.A(n_3838),
.B(n_3864),
.Y(n_5067)
);

AND2x2_ASAP7_75t_L g5068 ( 
.A(n_4596),
.B(n_4601),
.Y(n_5068)
);

BUFx3_ASAP7_75t_L g5069 ( 
.A(n_4610),
.Y(n_5069)
);

INVx2_ASAP7_75t_L g5070 ( 
.A(n_4053),
.Y(n_5070)
);

O2A1O1Ixp33_ASAP7_75t_L g5071 ( 
.A1(n_4028),
.A2(n_3899),
.B(n_3885),
.C(n_4091),
.Y(n_5071)
);

AOI21xp5_ASAP7_75t_L g5072 ( 
.A1(n_4375),
.A2(n_4435),
.B(n_4431),
.Y(n_5072)
);

OAI22xp5_ASAP7_75t_SL g5073 ( 
.A1(n_3896),
.A2(n_4540),
.B1(n_3834),
.B2(n_4247),
.Y(n_5073)
);

INVx1_ASAP7_75t_SL g5074 ( 
.A(n_4018),
.Y(n_5074)
);

INVxp67_ASAP7_75t_SL g5075 ( 
.A(n_4203),
.Y(n_5075)
);

INVx2_ASAP7_75t_L g5076 ( 
.A(n_4053),
.Y(n_5076)
);

NOR2xp67_ASAP7_75t_L g5077 ( 
.A(n_4324),
.B(n_4325),
.Y(n_5077)
);

INVx2_ASAP7_75t_L g5078 ( 
.A(n_4062),
.Y(n_5078)
);

AOI21xp5_ASAP7_75t_L g5079 ( 
.A1(n_4435),
.A2(n_4459),
.B(n_4438),
.Y(n_5079)
);

INVx2_ASAP7_75t_L g5080 ( 
.A(n_4062),
.Y(n_5080)
);

OR2x6_ASAP7_75t_L g5081 ( 
.A(n_4090),
.B(n_3856),
.Y(n_5081)
);

HB1xp67_ASAP7_75t_L g5082 ( 
.A(n_3880),
.Y(n_5082)
);

A2O1A1Ixp33_ASAP7_75t_L g5083 ( 
.A1(n_4169),
.A2(n_3885),
.B(n_4466),
.C(n_4125),
.Y(n_5083)
);

NAND3xp33_ASAP7_75t_L g5084 ( 
.A(n_4466),
.B(n_4470),
.C(n_4504),
.Y(n_5084)
);

NOR2xp33_ASAP7_75t_SL g5085 ( 
.A(n_4102),
.B(n_3969),
.Y(n_5085)
);

INVxp67_ASAP7_75t_SL g5086 ( 
.A(n_4198),
.Y(n_5086)
);

AOI22xp33_ASAP7_75t_L g5087 ( 
.A1(n_4149),
.A2(n_3916),
.B1(n_3983),
.B2(n_3892),
.Y(n_5087)
);

INVx3_ASAP7_75t_L g5088 ( 
.A(n_3858),
.Y(n_5088)
);

AOI21xp5_ASAP7_75t_L g5089 ( 
.A1(n_4438),
.A2(n_4474),
.B(n_4459),
.Y(n_5089)
);

NAND2xp5_ASAP7_75t_L g5090 ( 
.A(n_3870),
.B(n_3872),
.Y(n_5090)
);

NAND2xp5_ASAP7_75t_SL g5091 ( 
.A(n_4169),
.B(n_4081),
.Y(n_5091)
);

INVx2_ASAP7_75t_L g5092 ( 
.A(n_4062),
.Y(n_5092)
);

AND2x4_ASAP7_75t_L g5093 ( 
.A(n_3948),
.B(n_3950),
.Y(n_5093)
);

CKINVDCx20_ASAP7_75t_R g5094 ( 
.A(n_4173),
.Y(n_5094)
);

CKINVDCx20_ASAP7_75t_R g5095 ( 
.A(n_4173),
.Y(n_5095)
);

BUFx3_ASAP7_75t_L g5096 ( 
.A(n_4625),
.Y(n_5096)
);

INVx3_ASAP7_75t_L g5097 ( 
.A(n_3889),
.Y(n_5097)
);

BUFx2_ASAP7_75t_L g5098 ( 
.A(n_4334),
.Y(n_5098)
);

NAND2x1_ASAP7_75t_SL g5099 ( 
.A(n_3959),
.B(n_4114),
.Y(n_5099)
);

AND2x2_ASAP7_75t_L g5100 ( 
.A(n_4596),
.B(n_4601),
.Y(n_5100)
);

O2A1O1Ixp33_ASAP7_75t_L g5101 ( 
.A1(n_4116),
.A2(n_3892),
.B(n_3983),
.C(n_3916),
.Y(n_5101)
);

AO32x2_ASAP7_75t_L g5102 ( 
.A1(n_4129),
.A2(n_4138),
.A3(n_4590),
.B1(n_4143),
.B2(n_4058),
.Y(n_5102)
);

NOR2xp33_ASAP7_75t_L g5103 ( 
.A(n_4194),
.B(n_3896),
.Y(n_5103)
);

A2O1A1Ixp33_ASAP7_75t_L g5104 ( 
.A1(n_4121),
.A2(n_4125),
.B(n_4602),
.C(n_4134),
.Y(n_5104)
);

INVx2_ASAP7_75t_L g5105 ( 
.A(n_4062),
.Y(n_5105)
);

AND2x4_ASAP7_75t_L g5106 ( 
.A(n_3948),
.B(n_3950),
.Y(n_5106)
);

NAND2xp5_ASAP7_75t_SL g5107 ( 
.A(n_4470),
.B(n_3959),
.Y(n_5107)
);

O2A1O1Ixp33_ASAP7_75t_L g5108 ( 
.A1(n_4116),
.A2(n_4021),
.B(n_4076),
.C(n_4134),
.Y(n_5108)
);

AND2x4_ASAP7_75t_L g5109 ( 
.A(n_3948),
.B(n_3950),
.Y(n_5109)
);

AOI22xp33_ASAP7_75t_L g5110 ( 
.A1(n_4021),
.A2(n_4076),
.B1(n_4095),
.B2(n_4504),
.Y(n_5110)
);

AOI22xp33_ASAP7_75t_L g5111 ( 
.A1(n_4095),
.A2(n_4093),
.B1(n_4274),
.B2(n_4635),
.Y(n_5111)
);

BUFx3_ASAP7_75t_L g5112 ( 
.A(n_4625),
.Y(n_5112)
);

INVx2_ASAP7_75t_L g5113 ( 
.A(n_4080),
.Y(n_5113)
);

INVx4_ASAP7_75t_L g5114 ( 
.A(n_4451),
.Y(n_5114)
);

BUFx2_ASAP7_75t_L g5115 ( 
.A(n_4337),
.Y(n_5115)
);

AOI21xp5_ASAP7_75t_L g5116 ( 
.A1(n_4474),
.A2(n_4502),
.B(n_4500),
.Y(n_5116)
);

AOI21x1_ASAP7_75t_L g5117 ( 
.A1(n_4586),
.A2(n_4607),
.B(n_4515),
.Y(n_5117)
);

AND2x4_ASAP7_75t_L g5118 ( 
.A(n_3948),
.B(n_3950),
.Y(n_5118)
);

INVx2_ASAP7_75t_L g5119 ( 
.A(n_4080),
.Y(n_5119)
);

A2O1A1Ixp33_ASAP7_75t_L g5120 ( 
.A1(n_4121),
.A2(n_4602),
.B(n_4612),
.C(n_4128),
.Y(n_5120)
);

AND2x4_ASAP7_75t_L g5121 ( 
.A(n_3950),
.B(n_4268),
.Y(n_5121)
);

BUFx6f_ASAP7_75t_L g5122 ( 
.A(n_3848),
.Y(n_5122)
);

A2O1A1Ixp33_ASAP7_75t_L g5123 ( 
.A1(n_4612),
.A2(n_4128),
.B(n_4119),
.C(n_4464),
.Y(n_5123)
);

BUFx2_ASAP7_75t_L g5124 ( 
.A(n_4337),
.Y(n_5124)
);

OR2x6_ASAP7_75t_SL g5125 ( 
.A(n_3860),
.B(n_3861),
.Y(n_5125)
);

NAND2xp5_ASAP7_75t_L g5126 ( 
.A(n_3870),
.B(n_3872),
.Y(n_5126)
);

AND2x2_ASAP7_75t_L g5127 ( 
.A(n_4601),
.B(n_4659),
.Y(n_5127)
);

BUFx2_ASAP7_75t_L g5128 ( 
.A(n_3974),
.Y(n_5128)
);

AOI21xp5_ASAP7_75t_L g5129 ( 
.A1(n_4500),
.A2(n_4511),
.B(n_4502),
.Y(n_5129)
);

OAI21xp5_ASAP7_75t_L g5130 ( 
.A1(n_4107),
.A2(n_4079),
.B(n_4162),
.Y(n_5130)
);

BUFx12f_ASAP7_75t_L g5131 ( 
.A(n_4447),
.Y(n_5131)
);

O2A1O1Ixp33_ASAP7_75t_L g5132 ( 
.A1(n_4107),
.A2(n_4119),
.B(n_4219),
.C(n_4210),
.Y(n_5132)
);

AND2x2_ASAP7_75t_L g5133 ( 
.A(n_4659),
.B(n_4224),
.Y(n_5133)
);

BUFx12f_ASAP7_75t_L g5134 ( 
.A(n_4576),
.Y(n_5134)
);

O2A1O1Ixp33_ASAP7_75t_L g5135 ( 
.A1(n_4210),
.A2(n_4172),
.B(n_4590),
.C(n_4245),
.Y(n_5135)
);

NOR2xp33_ASAP7_75t_L g5136 ( 
.A(n_4409),
.B(n_4247),
.Y(n_5136)
);

AND2x2_ASAP7_75t_L g5137 ( 
.A(n_4659),
.B(n_4224),
.Y(n_5137)
);

NAND2xp5_ASAP7_75t_SL g5138 ( 
.A(n_4114),
.B(n_4611),
.Y(n_5138)
);

OAI22xp5_ASAP7_75t_L g5139 ( 
.A1(n_4112),
.A2(n_4109),
.B1(n_4101),
.B2(n_4464),
.Y(n_5139)
);

NOR2xp67_ASAP7_75t_L g5140 ( 
.A(n_4325),
.B(n_4501),
.Y(n_5140)
);

INVxp67_ASAP7_75t_L g5141 ( 
.A(n_4198),
.Y(n_5141)
);

BUFx6f_ASAP7_75t_L g5142 ( 
.A(n_3848),
.Y(n_5142)
);

AOI21xp5_ASAP7_75t_L g5143 ( 
.A1(n_4511),
.A2(n_4543),
.B(n_4535),
.Y(n_5143)
);

BUFx2_ASAP7_75t_L g5144 ( 
.A(n_3974),
.Y(n_5144)
);

BUFx2_ASAP7_75t_L g5145 ( 
.A(n_3974),
.Y(n_5145)
);

HB1xp67_ASAP7_75t_L g5146 ( 
.A(n_3880),
.Y(n_5146)
);

BUFx2_ASAP7_75t_L g5147 ( 
.A(n_3994),
.Y(n_5147)
);

BUFx2_ASAP7_75t_L g5148 ( 
.A(n_3994),
.Y(n_5148)
);

INVx5_ASAP7_75t_L g5149 ( 
.A(n_4052),
.Y(n_5149)
);

AND2x2_ASAP7_75t_L g5150 ( 
.A(n_4224),
.B(n_4263),
.Y(n_5150)
);

NAND3xp33_ASAP7_75t_L g5151 ( 
.A(n_4101),
.B(n_4112),
.C(n_4109),
.Y(n_5151)
);

NAND2xp5_ASAP7_75t_L g5152 ( 
.A(n_3906),
.B(n_3911),
.Y(n_5152)
);

O2A1O1Ixp33_ASAP7_75t_L g5153 ( 
.A1(n_4172),
.A2(n_4245),
.B(n_4093),
.C(n_4471),
.Y(n_5153)
);

NAND2xp5_ASAP7_75t_L g5154 ( 
.A(n_3906),
.B(n_3911),
.Y(n_5154)
);

NAND2xp5_ASAP7_75t_L g5155 ( 
.A(n_3914),
.B(n_3923),
.Y(n_5155)
);

A2O1A1Ixp33_ASAP7_75t_L g5156 ( 
.A1(n_4162),
.A2(n_4471),
.B(n_4157),
.C(n_4362),
.Y(n_5156)
);

NOR2x1_ASAP7_75t_L g5157 ( 
.A(n_4227),
.B(n_4563),
.Y(n_5157)
);

CKINVDCx8_ASAP7_75t_R g5158 ( 
.A(n_4486),
.Y(n_5158)
);

NOR2xp33_ASAP7_75t_L g5159 ( 
.A(n_4409),
.B(n_4469),
.Y(n_5159)
);

A2O1A1Ixp33_ASAP7_75t_L g5160 ( 
.A1(n_4157),
.A2(n_4362),
.B(n_4208),
.C(n_4213),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_3914),
.B(n_3923),
.Y(n_5161)
);

A2O1A1Ixp33_ASAP7_75t_L g5162 ( 
.A1(n_4208),
.A2(n_4213),
.B(n_4329),
.C(n_4260),
.Y(n_5162)
);

NAND3xp33_ASAP7_75t_L g5163 ( 
.A(n_4579),
.B(n_4259),
.C(n_3929),
.Y(n_5163)
);

AOI21xp5_ASAP7_75t_L g5164 ( 
.A1(n_4535),
.A2(n_4546),
.B(n_4543),
.Y(n_5164)
);

OAI22xp5_ASAP7_75t_L g5165 ( 
.A1(n_4260),
.A2(n_4259),
.B1(n_4381),
.B2(n_4365),
.Y(n_5165)
);

AOI21xp5_ASAP7_75t_L g5166 ( 
.A1(n_4546),
.A2(n_4177),
.B(n_4048),
.Y(n_5166)
);

AOI22xp33_ASAP7_75t_L g5167 ( 
.A1(n_4274),
.A2(n_4635),
.B1(n_4329),
.B2(n_3913),
.Y(n_5167)
);

NOR2x1_ASAP7_75t_L g5168 ( 
.A(n_4563),
.B(n_4217),
.Y(n_5168)
);

INVxp67_ASAP7_75t_L g5169 ( 
.A(n_4200),
.Y(n_5169)
);

BUFx8_ASAP7_75t_SL g5170 ( 
.A(n_4547),
.Y(n_5170)
);

CKINVDCx5p33_ASAP7_75t_R g5171 ( 
.A(n_4161),
.Y(n_5171)
);

NAND2xp5_ASAP7_75t_L g5172 ( 
.A(n_3928),
.B(n_3934),
.Y(n_5172)
);

BUFx4f_ASAP7_75t_SL g5173 ( 
.A(n_4360),
.Y(n_5173)
);

AOI21xp5_ASAP7_75t_L g5174 ( 
.A1(n_4048),
.A2(n_4277),
.B(n_4177),
.Y(n_5174)
);

NOR2xp33_ASAP7_75t_L g5175 ( 
.A(n_4469),
.B(n_4477),
.Y(n_5175)
);

OAI21x1_ASAP7_75t_L g5176 ( 
.A1(n_4277),
.A2(n_3966),
.B(n_4201),
.Y(n_5176)
);

BUFx2_ASAP7_75t_L g5177 ( 
.A(n_3994),
.Y(n_5177)
);

AND2x2_ASAP7_75t_SL g5178 ( 
.A(n_4102),
.B(n_4011),
.Y(n_5178)
);

CKINVDCx5p33_ASAP7_75t_R g5179 ( 
.A(n_4294),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_4519),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_3928),
.B(n_3934),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_SL g5182 ( 
.A(n_4318),
.B(n_4217),
.Y(n_5182)
);

OAI22xp5_ASAP7_75t_L g5183 ( 
.A1(n_4365),
.A2(n_4381),
.B1(n_4528),
.B2(n_4387),
.Y(n_5183)
);

INVxp67_ASAP7_75t_SL g5184 ( 
.A(n_4501),
.Y(n_5184)
);

AOI21xp5_ASAP7_75t_L g5185 ( 
.A1(n_4433),
.A2(n_3966),
.B(n_3929),
.Y(n_5185)
);

INVxp67_ASAP7_75t_L g5186 ( 
.A(n_4200),
.Y(n_5186)
);

OAI21xp33_ASAP7_75t_SL g5187 ( 
.A1(n_4632),
.A2(n_3939),
.B(n_3935),
.Y(n_5187)
);

INVx4_ASAP7_75t_L g5188 ( 
.A(n_4451),
.Y(n_5188)
);

AOI21xp5_ASAP7_75t_L g5189 ( 
.A1(n_4433),
.A2(n_3966),
.B(n_3929),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_4519),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_4533),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_4533),
.Y(n_5192)
);

A2O1A1Ixp33_ASAP7_75t_L g5193 ( 
.A1(n_4579),
.A2(n_4648),
.B(n_4593),
.C(n_4191),
.Y(n_5193)
);

AND2x2_ASAP7_75t_L g5194 ( 
.A(n_4263),
.B(n_4661),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_3846),
.Y(n_5195)
);

OAI21x1_ASAP7_75t_SL g5196 ( 
.A1(n_4629),
.A2(n_4528),
.B(n_4573),
.Y(n_5196)
);

INVx5_ASAP7_75t_L g5197 ( 
.A(n_4052),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_3846),
.Y(n_5198)
);

AND2x2_ASAP7_75t_L g5199 ( 
.A(n_4263),
.B(n_4661),
.Y(n_5199)
);

NOR2xp33_ASAP7_75t_SL g5200 ( 
.A(n_4102),
.B(n_3969),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_3915),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_3915),
.Y(n_5202)
);

BUFx8_ASAP7_75t_L g5203 ( 
.A(n_4231),
.Y(n_5203)
);

HB1xp67_ASAP7_75t_L g5204 ( 
.A(n_4411),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_3917),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_3917),
.Y(n_5206)
);

OAI22xp5_ASAP7_75t_L g5207 ( 
.A1(n_4372),
.A2(n_4387),
.B1(n_3844),
.B2(n_3849),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_L g5208 ( 
.A(n_3935),
.B(n_3939),
.Y(n_5208)
);

BUFx2_ASAP7_75t_L g5209 ( 
.A(n_4016),
.Y(n_5209)
);

BUFx4f_ASAP7_75t_L g5210 ( 
.A(n_4451),
.Y(n_5210)
);

INVx1_ASAP7_75t_SL g5211 ( 
.A(n_4055),
.Y(n_5211)
);

OAI22xp5_ASAP7_75t_L g5212 ( 
.A1(n_4372),
.A2(n_3844),
.B1(n_3849),
.B2(n_4540),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_3919),
.Y(n_5213)
);

AOI22xp33_ASAP7_75t_L g5214 ( 
.A1(n_4274),
.A2(n_4593),
.B1(n_4664),
.B2(n_4477),
.Y(n_5214)
);

NAND2xp5_ASAP7_75t_L g5215 ( 
.A(n_3940),
.B(n_3945),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_3919),
.Y(n_5216)
);

BUFx2_ASAP7_75t_L g5217 ( 
.A(n_4016),
.Y(n_5217)
);

INVx3_ASAP7_75t_L g5218 ( 
.A(n_3921),
.Y(n_5218)
);

OAI22xp5_ASAP7_75t_L g5219 ( 
.A1(n_3965),
.A2(n_4207),
.B1(n_4406),
.B2(n_4274),
.Y(n_5219)
);

NAND2xp5_ASAP7_75t_L g5220 ( 
.A(n_3940),
.B(n_3945),
.Y(n_5220)
);

NOR2x1_ASAP7_75t_L g5221 ( 
.A(n_4560),
.B(n_4636),
.Y(n_5221)
);

AOI21xp5_ASAP7_75t_L g5222 ( 
.A1(n_3922),
.A2(n_4530),
.B(n_4495),
.Y(n_5222)
);

BUFx2_ASAP7_75t_L g5223 ( 
.A(n_4016),
.Y(n_5223)
);

BUFx6f_ASAP7_75t_SL g5224 ( 
.A(n_4102),
.Y(n_5224)
);

AND2x6_ASAP7_75t_L g5225 ( 
.A(n_4568),
.B(n_4487),
.Y(n_5225)
);

NOR2xp33_ASAP7_75t_L g5226 ( 
.A(n_3922),
.B(n_4638),
.Y(n_5226)
);

OAI22xp5_ASAP7_75t_SL g5227 ( 
.A1(n_4294),
.A2(n_4196),
.B1(n_3904),
.B2(n_3965),
.Y(n_5227)
);

INVx3_ASAP7_75t_L g5228 ( 
.A(n_3921),
.Y(n_5228)
);

INVx1_ASAP7_75t_L g5229 ( 
.A(n_3920),
.Y(n_5229)
);

INVx3_ASAP7_75t_L g5230 ( 
.A(n_3921),
.Y(n_5230)
);

OAI22xp5_ASAP7_75t_L g5231 ( 
.A1(n_4207),
.A2(n_4406),
.B1(n_4327),
.B2(n_4182),
.Y(n_5231)
);

OAI22xp5_ASAP7_75t_L g5232 ( 
.A1(n_4182),
.A2(n_4327),
.B1(n_3857),
.B2(n_3904),
.Y(n_5232)
);

OAI22xp5_ASAP7_75t_L g5233 ( 
.A1(n_4182),
.A2(n_4327),
.B1(n_3857),
.B2(n_4239),
.Y(n_5233)
);

INVx1_ASAP7_75t_L g5234 ( 
.A(n_3920),
.Y(n_5234)
);

INVxp67_ASAP7_75t_SL g5235 ( 
.A(n_4495),
.Y(n_5235)
);

NOR2xp33_ASAP7_75t_L g5236 ( 
.A(n_4636),
.B(n_3951),
.Y(n_5236)
);

BUFx2_ASAP7_75t_L g5237 ( 
.A(n_4017),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_3926),
.Y(n_5238)
);

INVx3_ASAP7_75t_L g5239 ( 
.A(n_3921),
.Y(n_5239)
);

NAND2xp5_ASAP7_75t_SL g5240 ( 
.A(n_4318),
.B(n_4632),
.Y(n_5240)
);

CKINVDCx5p33_ASAP7_75t_R g5241 ( 
.A(n_3995),
.Y(n_5241)
);

NAND2xp5_ASAP7_75t_L g5242 ( 
.A(n_3951),
.B(n_3956),
.Y(n_5242)
);

HB1xp67_ASAP7_75t_L g5243 ( 
.A(n_4411),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_3926),
.Y(n_5244)
);

INVx3_ASAP7_75t_L g5245 ( 
.A(n_3924),
.Y(n_5245)
);

INVx1_ASAP7_75t_SL g5246 ( 
.A(n_4055),
.Y(n_5246)
);

NOR2xp33_ASAP7_75t_L g5247 ( 
.A(n_3956),
.B(n_3962),
.Y(n_5247)
);

AOI22xp33_ASAP7_75t_L g5248 ( 
.A1(n_4664),
.A2(n_4503),
.B1(n_4499),
.B2(n_4346),
.Y(n_5248)
);

OA22x2_ASAP7_75t_L g5249 ( 
.A1(n_4565),
.A2(n_4641),
.B1(n_4626),
.B2(n_4549),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_3927),
.Y(n_5250)
);

NAND2x1p5_ASAP7_75t_L g5251 ( 
.A(n_4672),
.B(n_3882),
.Y(n_5251)
);

BUFx2_ASAP7_75t_L g5252 ( 
.A(n_4017),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_SL g5253 ( 
.A(n_4570),
.B(n_4191),
.Y(n_5253)
);

AOI222xp33_ASAP7_75t_L g5254 ( 
.A1(n_4400),
.A2(n_4499),
.B1(n_4503),
.B2(n_4570),
.C1(n_3860),
.C2(n_3861),
.Y(n_5254)
);

CKINVDCx5p33_ASAP7_75t_R g5255 ( 
.A(n_3995),
.Y(n_5255)
);

INVx1_ASAP7_75t_L g5256 ( 
.A(n_3927),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_3947),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_3947),
.Y(n_5258)
);

NAND2xp5_ASAP7_75t_SL g5259 ( 
.A(n_4140),
.B(n_4145),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_L g5260 ( 
.A(n_3962),
.B(n_3968),
.Y(n_5260)
);

OAI22xp5_ASAP7_75t_L g5261 ( 
.A1(n_4236),
.A2(n_4249),
.B1(n_4251),
.B2(n_4239),
.Y(n_5261)
);

AND2x4_ASAP7_75t_L g5262 ( 
.A(n_4268),
.B(n_4206),
.Y(n_5262)
);

A2O1A1Ixp33_ASAP7_75t_SL g5263 ( 
.A1(n_4269),
.A2(n_4403),
.B(n_4457),
.C(n_4383),
.Y(n_5263)
);

OAI21xp33_ASAP7_75t_L g5264 ( 
.A1(n_3862),
.A2(n_3977),
.B(n_3968),
.Y(n_5264)
);

INVxp67_ASAP7_75t_L g5265 ( 
.A(n_4216),
.Y(n_5265)
);

OR2x6_ASAP7_75t_L g5266 ( 
.A(n_4090),
.B(n_3856),
.Y(n_5266)
);

AOI21xp5_ASAP7_75t_L g5267 ( 
.A1(n_4530),
.A2(n_4201),
.B(n_4408),
.Y(n_5267)
);

BUFx2_ASAP7_75t_L g5268 ( 
.A(n_4017),
.Y(n_5268)
);

NOR2xp33_ASAP7_75t_L g5269 ( 
.A(n_3977),
.B(n_3978),
.Y(n_5269)
);

AOI21xp5_ASAP7_75t_L g5270 ( 
.A1(n_4408),
.A2(n_3862),
.B(n_4315),
.Y(n_5270)
);

AOI22xp5_ASAP7_75t_L g5271 ( 
.A1(n_3875),
.A2(n_4624),
.B1(n_4626),
.B2(n_4674),
.Y(n_5271)
);

AND2x2_ASAP7_75t_L g5272 ( 
.A(n_4663),
.B(n_4352),
.Y(n_5272)
);

NAND2xp5_ASAP7_75t_L g5273 ( 
.A(n_3978),
.B(n_3987),
.Y(n_5273)
);

NAND2xp5_ASAP7_75t_SL g5274 ( 
.A(n_4140),
.B(n_4145),
.Y(n_5274)
);

NAND2xp5_ASAP7_75t_L g5275 ( 
.A(n_3987),
.B(n_3991),
.Y(n_5275)
);

INVx3_ASAP7_75t_L g5276 ( 
.A(n_3924),
.Y(n_5276)
);

OAI22xp5_ASAP7_75t_L g5277 ( 
.A1(n_4236),
.A2(n_4251),
.B1(n_4256),
.B2(n_4249),
.Y(n_5277)
);

AO32x2_ASAP7_75t_L g5278 ( 
.A1(n_4129),
.A2(n_4138),
.A3(n_4143),
.B1(n_4058),
.B2(n_4012),
.Y(n_5278)
);

O2A1O1Ixp33_ASAP7_75t_L g5279 ( 
.A1(n_4560),
.A2(n_4674),
.B(n_4591),
.C(n_4665),
.Y(n_5279)
);

AOI21xp5_ASAP7_75t_L g5280 ( 
.A1(n_4315),
.A2(n_4079),
.B(n_4333),
.Y(n_5280)
);

A2O1A1Ixp33_ASAP7_75t_L g5281 ( 
.A1(n_4648),
.A2(n_4400),
.B(n_4641),
.C(n_4573),
.Y(n_5281)
);

BUFx2_ASAP7_75t_L g5282 ( 
.A(n_4030),
.Y(n_5282)
);

INVx8_ASAP7_75t_L g5283 ( 
.A(n_4052),
.Y(n_5283)
);

NAND2xp5_ASAP7_75t_L g5284 ( 
.A(n_3991),
.B(n_3992),
.Y(n_5284)
);

O2A1O1Ixp5_ASAP7_75t_SL g5285 ( 
.A1(n_4479),
.A2(n_4515),
.B(n_4607),
.C(n_4586),
.Y(n_5285)
);

A2O1A1Ixp33_ASAP7_75t_L g5286 ( 
.A1(n_4665),
.A2(n_4551),
.B(n_4204),
.C(n_4594),
.Y(n_5286)
);

AND2x2_ASAP7_75t_L g5287 ( 
.A(n_4663),
.B(n_4352),
.Y(n_5287)
);

INVx1_ASAP7_75t_L g5288 ( 
.A(n_3949),
.Y(n_5288)
);

O2A1O1Ixp5_ASAP7_75t_SL g5289 ( 
.A1(n_4591),
.A2(n_4633),
.B(n_4160),
.C(n_4403),
.Y(n_5289)
);

HB1xp67_ASAP7_75t_L g5290 ( 
.A(n_4434),
.Y(n_5290)
);

AOI21xp5_ASAP7_75t_L g5291 ( 
.A1(n_4079),
.A2(n_4336),
.B(n_4333),
.Y(n_5291)
);

AOI21xp5_ASAP7_75t_L g5292 ( 
.A1(n_4336),
.A2(n_4341),
.B(n_3996),
.Y(n_5292)
);

NAND2xp5_ASAP7_75t_SL g5293 ( 
.A(n_4282),
.B(n_4314),
.Y(n_5293)
);

HB1xp67_ASAP7_75t_L g5294 ( 
.A(n_4434),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_3992),
.B(n_3996),
.Y(n_5295)
);

AOI22xp5_ASAP7_75t_L g5296 ( 
.A1(n_3875),
.A2(n_4624),
.B1(n_4571),
.B2(n_4205),
.Y(n_5296)
);

NAND2xp5_ASAP7_75t_L g5297 ( 
.A(n_4004),
.B(n_4019),
.Y(n_5297)
);

AOI22xp33_ASAP7_75t_L g5298 ( 
.A1(n_4576),
.A2(n_4565),
.B1(n_4571),
.B2(n_4569),
.Y(n_5298)
);

AOI21xp5_ASAP7_75t_L g5299 ( 
.A1(n_4341),
.A2(n_4019),
.B(n_4004),
.Y(n_5299)
);

NAND2xp5_ASAP7_75t_L g5300 ( 
.A(n_4023),
.B(n_4029),
.Y(n_5300)
);

AND2x6_ASAP7_75t_SL g5301 ( 
.A(n_4285),
.B(n_3941),
.Y(n_5301)
);

NOR2xp33_ASAP7_75t_L g5302 ( 
.A(n_4023),
.B(n_4029),
.Y(n_5302)
);

OAI22xp5_ASAP7_75t_L g5303 ( 
.A1(n_4256),
.A2(n_4270),
.B1(n_4296),
.B2(n_4267),
.Y(n_5303)
);

HB1xp67_ASAP7_75t_L g5304 ( 
.A(n_3943),
.Y(n_5304)
);

NAND2xp5_ASAP7_75t_L g5305 ( 
.A(n_4035),
.B(n_4041),
.Y(n_5305)
);

OAI22xp5_ASAP7_75t_L g5306 ( 
.A1(n_4267),
.A2(n_4296),
.B1(n_4297),
.B2(n_4270),
.Y(n_5306)
);

INVx3_ASAP7_75t_L g5307 ( 
.A(n_3924),
.Y(n_5307)
);

BUFx2_ASAP7_75t_L g5308 ( 
.A(n_4030),
.Y(n_5308)
);

AOI21xp5_ASAP7_75t_L g5309 ( 
.A1(n_4035),
.A2(n_4042),
.B(n_4041),
.Y(n_5309)
);

NOR2x1_ASAP7_75t_SL g5310 ( 
.A(n_4486),
.B(n_4629),
.Y(n_5310)
);

AOI21x1_ASAP7_75t_L g5311 ( 
.A1(n_4150),
.A2(n_4603),
.B(n_4594),
.Y(n_5311)
);

INVx3_ASAP7_75t_L g5312 ( 
.A(n_3924),
.Y(n_5312)
);

NAND2xp5_ASAP7_75t_L g5313 ( 
.A(n_4042),
.B(n_4050),
.Y(n_5313)
);

O2A1O1Ixp33_ASAP7_75t_L g5314 ( 
.A1(n_4204),
.A2(n_4569),
.B(n_4457),
.C(n_4383),
.Y(n_5314)
);

O2A1O1Ixp33_ASAP7_75t_L g5315 ( 
.A1(n_4050),
.A2(n_4065),
.B(n_4067),
.C(n_4051),
.Y(n_5315)
);

NOR2xp33_ASAP7_75t_R g5316 ( 
.A(n_4393),
.B(n_4454),
.Y(n_5316)
);

INVx6_ASAP7_75t_L g5317 ( 
.A(n_4002),
.Y(n_5317)
);

AND2x6_ASAP7_75t_L g5318 ( 
.A(n_4568),
.B(n_4487),
.Y(n_5318)
);

OAI22xp5_ASAP7_75t_L g5319 ( 
.A1(n_4297),
.A2(n_4313),
.B1(n_4065),
.B2(n_4067),
.Y(n_5319)
);

OAI22xp5_ASAP7_75t_L g5320 ( 
.A1(n_4313),
.A2(n_4072),
.B1(n_4082),
.B2(n_4051),
.Y(n_5320)
);

INVx1_ASAP7_75t_L g5321 ( 
.A(n_3949),
.Y(n_5321)
);

BUFx2_ASAP7_75t_L g5322 ( 
.A(n_4030),
.Y(n_5322)
);

INVx1_ASAP7_75t_L g5323 ( 
.A(n_3952),
.Y(n_5323)
);

CKINVDCx5p33_ASAP7_75t_R g5324 ( 
.A(n_4285),
.Y(n_5324)
);

OAI22xp5_ASAP7_75t_L g5325 ( 
.A1(n_4072),
.A2(n_4084),
.B1(n_4085),
.B2(n_4082),
.Y(n_5325)
);

BUFx2_ASAP7_75t_L g5326 ( 
.A(n_4063),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_3952),
.Y(n_5327)
);

AOI22xp5_ASAP7_75t_L g5328 ( 
.A1(n_4205),
.A2(n_4578),
.B1(n_4011),
.B2(n_3971),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_L g5329 ( 
.A(n_4084),
.B(n_4085),
.Y(n_5329)
);

AOI221xp5_ASAP7_75t_L g5330 ( 
.A1(n_4099),
.A2(n_4104),
.B1(n_4127),
.B2(n_4118),
.C(n_4115),
.Y(n_5330)
);

NAND2xp5_ASAP7_75t_L g5331 ( 
.A(n_4099),
.B(n_4104),
.Y(n_5331)
);

AOI21xp5_ASAP7_75t_L g5332 ( 
.A1(n_4115),
.A2(n_4127),
.B(n_4118),
.Y(n_5332)
);

NAND2xp5_ASAP7_75t_SL g5333 ( 
.A(n_4282),
.B(n_4314),
.Y(n_5333)
);

AOI21xp5_ASAP7_75t_L g5334 ( 
.A1(n_4130),
.A2(n_4139),
.B(n_4136),
.Y(n_5334)
);

INVx1_ASAP7_75t_SL g5335 ( 
.A(n_3971),
.Y(n_5335)
);

BUFx4f_ASAP7_75t_SL g5336 ( 
.A(n_4360),
.Y(n_5336)
);

AOI22xp33_ASAP7_75t_L g5337 ( 
.A1(n_4565),
.A2(n_4597),
.B1(n_4350),
.B2(n_4527),
.Y(n_5337)
);

BUFx12f_ASAP7_75t_L g5338 ( 
.A(n_4547),
.Y(n_5338)
);

O2A1O1Ixp33_ASAP7_75t_L g5339 ( 
.A1(n_4130),
.A2(n_4139),
.B(n_4141),
.C(n_4136),
.Y(n_5339)
);

BUFx12f_ASAP7_75t_L g5340 ( 
.A(n_4587),
.Y(n_5340)
);

NAND2xp5_ASAP7_75t_L g5341 ( 
.A(n_4141),
.B(n_4144),
.Y(n_5341)
);

NAND2xp5_ASAP7_75t_SL g5342 ( 
.A(n_4144),
.B(n_4147),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_3954),
.Y(n_5343)
);

OAI22x1_ASAP7_75t_L g5344 ( 
.A1(n_4551),
.A2(n_4153),
.B1(n_3903),
.B2(n_4290),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_3954),
.Y(n_5345)
);

NAND2xp5_ASAP7_75t_L g5346 ( 
.A(n_4147),
.B(n_4170),
.Y(n_5346)
);

NAND2xp5_ASAP7_75t_L g5347 ( 
.A(n_4170),
.B(n_4175),
.Y(n_5347)
);

AOI22xp33_ASAP7_75t_L g5348 ( 
.A1(n_4597),
.A2(n_4350),
.B1(n_4527),
.B2(n_4011),
.Y(n_5348)
);

INVx2_ASAP7_75t_SL g5349 ( 
.A(n_4492),
.Y(n_5349)
);

INVx1_ASAP7_75t_SL g5350 ( 
.A(n_3854),
.Y(n_5350)
);

NAND2xp5_ASAP7_75t_L g5351 ( 
.A(n_4175),
.B(n_4179),
.Y(n_5351)
);

AND2x4_ASAP7_75t_L g5352 ( 
.A(n_4268),
.B(n_4206),
.Y(n_5352)
);

NAND2x2_ASAP7_75t_L g5353 ( 
.A(n_3933),
.B(n_4202),
.Y(n_5353)
);

O2A1O1Ixp33_ASAP7_75t_L g5354 ( 
.A1(n_4179),
.A2(n_4388),
.B(n_4368),
.C(n_4603),
.Y(n_5354)
);

BUFx2_ASAP7_75t_L g5355 ( 
.A(n_4063),
.Y(n_5355)
);

BUFx12f_ASAP7_75t_L g5356 ( 
.A(n_4587),
.Y(n_5356)
);

BUFx2_ASAP7_75t_L g5357 ( 
.A(n_4063),
.Y(n_5357)
);

AOI21xp5_ASAP7_75t_L g5358 ( 
.A1(n_4631),
.A2(n_4673),
.B(n_4523),
.Y(n_5358)
);

NOR2xp33_ASAP7_75t_L g5359 ( 
.A(n_4606),
.B(n_4407),
.Y(n_5359)
);

INVx4_ASAP7_75t_L g5360 ( 
.A(n_4442),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_3955),
.Y(n_5361)
);

AOI22xp33_ASAP7_75t_L g5362 ( 
.A1(n_4011),
.A2(n_3980),
.B1(n_3882),
.B2(n_4578),
.Y(n_5362)
);

INVx4_ASAP7_75t_L g5363 ( 
.A(n_4442),
.Y(n_5363)
);

A2O1A1Ixp33_ASAP7_75t_L g5364 ( 
.A1(n_4551),
.A2(n_4668),
.B(n_4588),
.C(n_4031),
.Y(n_5364)
);

INVx1_ASAP7_75t_L g5365 ( 
.A(n_3955),
.Y(n_5365)
);

AOI22xp33_ASAP7_75t_L g5366 ( 
.A1(n_3882),
.A2(n_3980),
.B1(n_4388),
.B2(n_4368),
.Y(n_5366)
);

A2O1A1Ixp33_ASAP7_75t_L g5367 ( 
.A1(n_4668),
.A2(n_4588),
.B(n_4031),
.C(n_4096),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_3957),
.Y(n_5368)
);

NAND2xp5_ASAP7_75t_SL g5369 ( 
.A(n_3981),
.B(n_4031),
.Y(n_5369)
);

BUFx2_ASAP7_75t_L g5370 ( 
.A(n_4074),
.Y(n_5370)
);

O2A1O1Ixp33_ASAP7_75t_L g5371 ( 
.A1(n_4647),
.A2(n_4523),
.B(n_4189),
.C(n_4190),
.Y(n_5371)
);

HB1xp67_ASAP7_75t_L g5372 ( 
.A(n_3943),
.Y(n_5372)
);

AOI21xp5_ASAP7_75t_L g5373 ( 
.A1(n_4631),
.A2(n_4673),
.B(n_4031),
.Y(n_5373)
);

INVx1_ASAP7_75t_L g5374 ( 
.A(n_3957),
.Y(n_5374)
);

BUFx3_ASAP7_75t_L g5375 ( 
.A(n_4658),
.Y(n_5375)
);

NAND2x1p5_ASAP7_75t_L g5376 ( 
.A(n_4672),
.B(n_3882),
.Y(n_5376)
);

INVx1_ASAP7_75t_L g5377 ( 
.A(n_3960),
.Y(n_5377)
);

OAI22xp5_ASAP7_75t_L g5378 ( 
.A1(n_4606),
.A2(n_4426),
.B1(n_4407),
.B2(n_4031),
.Y(n_5378)
);

OAI22xp5_ASAP7_75t_L g5379 ( 
.A1(n_4407),
.A2(n_4426),
.B1(n_4096),
.B2(n_3981),
.Y(n_5379)
);

OAI21xp5_ASAP7_75t_L g5380 ( 
.A1(n_4647),
.A2(n_4584),
.B(n_4160),
.Y(n_5380)
);

OAI22xp5_ASAP7_75t_L g5381 ( 
.A1(n_4426),
.A2(n_4096),
.B1(n_3981),
.B2(n_4644),
.Y(n_5381)
);

BUFx3_ASAP7_75t_L g5382 ( 
.A(n_4002),
.Y(n_5382)
);

INVx1_ASAP7_75t_L g5383 ( 
.A(n_3960),
.Y(n_5383)
);

OAI22xp33_ASAP7_75t_L g5384 ( 
.A1(n_4498),
.A2(n_3953),
.B1(n_4096),
.B2(n_3981),
.Y(n_5384)
);

OAI22xp5_ASAP7_75t_L g5385 ( 
.A1(n_3981),
.A2(n_4096),
.B1(n_4657),
.B2(n_4644),
.Y(n_5385)
);

NOR2xp33_ASAP7_75t_L g5386 ( 
.A(n_3829),
.B(n_3894),
.Y(n_5386)
);

INVx1_ASAP7_75t_L g5387 ( 
.A(n_3961),
.Y(n_5387)
);

AOI21xp33_ASAP7_75t_L g5388 ( 
.A1(n_4633),
.A2(n_4190),
.B(n_4189),
.Y(n_5388)
);

O2A1O1Ixp33_ASAP7_75t_L g5389 ( 
.A1(n_3829),
.A2(n_3894),
.B(n_4580),
.C(n_4216),
.Y(n_5389)
);

INVx8_ASAP7_75t_L g5390 ( 
.A(n_4052),
.Y(n_5390)
);

NAND2xp5_ASAP7_75t_L g5391 ( 
.A(n_4452),
.B(n_4524),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_3961),
.Y(n_5392)
);

AND2x4_ASAP7_75t_L g5393 ( 
.A(n_4268),
.B(n_4206),
.Y(n_5393)
);

NAND2xp5_ASAP7_75t_L g5394 ( 
.A(n_4452),
.B(n_4524),
.Y(n_5394)
);

NAND2xp5_ASAP7_75t_SL g5395 ( 
.A(n_4584),
.B(n_4662),
.Y(n_5395)
);

OAI22xp33_ASAP7_75t_L g5396 ( 
.A1(n_4498),
.A2(n_3953),
.B1(n_4454),
.B2(n_4644),
.Y(n_5396)
);

INVx1_ASAP7_75t_L g5397 ( 
.A(n_3963),
.Y(n_5397)
);

A2O1A1Ixp33_ASAP7_75t_SL g5398 ( 
.A1(n_3972),
.A2(n_4033),
.B(n_4026),
.C(n_4614),
.Y(n_5398)
);

HB1xp67_ASAP7_75t_L g5399 ( 
.A(n_4639),
.Y(n_5399)
);

AOI21xp5_ASAP7_75t_L g5400 ( 
.A1(n_4349),
.A2(n_4657),
.B(n_4644),
.Y(n_5400)
);

NOR2xp33_ASAP7_75t_L g5401 ( 
.A(n_4437),
.B(n_4448),
.Y(n_5401)
);

A2O1A1Ixp33_ASAP7_75t_SL g5402 ( 
.A1(n_3972),
.A2(n_4033),
.B(n_4026),
.C(n_4614),
.Y(n_5402)
);

O2A1O1Ixp33_ASAP7_75t_SL g5403 ( 
.A1(n_4188),
.A2(n_4366),
.B(n_3970),
.C(n_4003),
.Y(n_5403)
);

AOI21xp5_ASAP7_75t_L g5404 ( 
.A1(n_4349),
.A2(n_4657),
.B(n_4644),
.Y(n_5404)
);

NAND2xp5_ASAP7_75t_L g5405 ( 
.A(n_4452),
.B(n_4529),
.Y(n_5405)
);

OAI22xp5_ASAP7_75t_L g5406 ( 
.A1(n_4657),
.A2(n_3980),
.B1(n_3882),
.B2(n_4222),
.Y(n_5406)
);

AND2x2_ASAP7_75t_L g5407 ( 
.A(n_4663),
.B(n_4355),
.Y(n_5407)
);

CKINVDCx16_ASAP7_75t_R g5408 ( 
.A(n_3839),
.Y(n_5408)
);

AOI21xp5_ASAP7_75t_L g5409 ( 
.A1(n_4657),
.A2(n_4075),
.B(n_4074),
.Y(n_5409)
);

AND2x6_ASAP7_75t_L g5410 ( 
.A(n_4568),
.B(n_4487),
.Y(n_5410)
);

NOR2xp33_ASAP7_75t_L g5411 ( 
.A(n_4437),
.B(n_4448),
.Y(n_5411)
);

NAND2xp5_ASAP7_75t_L g5412 ( 
.A(n_4529),
.B(n_4539),
.Y(n_5412)
);

O2A1O1Ixp33_ASAP7_75t_L g5413 ( 
.A1(n_4580),
.A2(n_4153),
.B(n_3903),
.C(n_4188),
.Y(n_5413)
);

OAI22xp5_ASAP7_75t_SL g5414 ( 
.A1(n_4538),
.A2(n_3839),
.B1(n_4094),
.B2(n_3958),
.Y(n_5414)
);

NAND2xp5_ASAP7_75t_L g5415 ( 
.A(n_4539),
.B(n_4542),
.Y(n_5415)
);

NOR2xp33_ASAP7_75t_L g5416 ( 
.A(n_4437),
.B(n_4448),
.Y(n_5416)
);

AOI21xp5_ASAP7_75t_L g5417 ( 
.A1(n_4074),
.A2(n_4075),
.B(n_3990),
.Y(n_5417)
);

AO32x1_ASAP7_75t_L g5418 ( 
.A1(n_3970),
.A2(n_4003),
.A3(n_3990),
.B1(n_3932),
.B2(n_3946),
.Y(n_5418)
);

INVx1_ASAP7_75t_SL g5419 ( 
.A(n_3854),
.Y(n_5419)
);

BUFx2_ASAP7_75t_L g5420 ( 
.A(n_4075),
.Y(n_5420)
);

OR2x2_ASAP7_75t_L g5421 ( 
.A(n_4006),
.B(n_3854),
.Y(n_5421)
);

CKINVDCx14_ASAP7_75t_R g5422 ( 
.A(n_4360),
.Y(n_5422)
);

AOI21xp5_ASAP7_75t_L g5423 ( 
.A1(n_3970),
.A2(n_4003),
.B(n_3990),
.Y(n_5423)
);

AOI221xp5_ASAP7_75t_L g5424 ( 
.A1(n_4510),
.A2(n_4526),
.B1(n_4531),
.B2(n_4525),
.C(n_4521),
.Y(n_5424)
);

AND2x4_ASAP7_75t_L g5425 ( 
.A(n_4206),
.B(n_3973),
.Y(n_5425)
);

AOI21x1_ASAP7_75t_L g5426 ( 
.A1(n_4150),
.A2(n_3998),
.B(n_4633),
.Y(n_5426)
);

BUFx2_ASAP7_75t_L g5427 ( 
.A(n_3843),
.Y(n_5427)
);

CKINVDCx5p33_ASAP7_75t_R g5428 ( 
.A(n_4538),
.Y(n_5428)
);

BUFx2_ASAP7_75t_L g5429 ( 
.A(n_3843),
.Y(n_5429)
);

OAI22xp33_ASAP7_75t_L g5430 ( 
.A1(n_3980),
.A2(n_4662),
.B1(n_3958),
.B2(n_4094),
.Y(n_5430)
);

INVx2_ASAP7_75t_SL g5431 ( 
.A(n_4517),
.Y(n_5431)
);

NOR2xp33_ASAP7_75t_L g5432 ( 
.A(n_4061),
.B(n_4100),
.Y(n_5432)
);

NAND2xp5_ASAP7_75t_L g5433 ( 
.A(n_4542),
.B(n_4550),
.Y(n_5433)
);

BUFx2_ASAP7_75t_SL g5434 ( 
.A(n_4672),
.Y(n_5434)
);

INVxp67_ASAP7_75t_L g5435 ( 
.A(n_4639),
.Y(n_5435)
);

AND2x4_ASAP7_75t_L g5436 ( 
.A(n_4206),
.B(n_3973),
.Y(n_5436)
);

AOI22xp33_ASAP7_75t_L g5437 ( 
.A1(n_3980),
.A2(n_3839),
.B1(n_4094),
.B2(n_3958),
.Y(n_5437)
);

INVx4_ASAP7_75t_L g5438 ( 
.A(n_4442),
.Y(n_5438)
);

NOR2xp67_ASAP7_75t_SL g5439 ( 
.A(n_3958),
.B(n_4094),
.Y(n_5439)
);

INVx1_ASAP7_75t_SL g5440 ( 
.A(n_3989),
.Y(n_5440)
);

CKINVDCx20_ASAP7_75t_R g5441 ( 
.A(n_4397),
.Y(n_5441)
);

AOI22xp5_ASAP7_75t_L g5442 ( 
.A1(n_4615),
.A2(n_4627),
.B1(n_4621),
.B2(n_4623),
.Y(n_5442)
);

NAND2xp5_ASAP7_75t_L g5443 ( 
.A(n_4550),
.B(n_4554),
.Y(n_5443)
);

NAND2xp5_ASAP7_75t_L g5444 ( 
.A(n_4554),
.B(n_4555),
.Y(n_5444)
);

INVxp67_ASAP7_75t_SL g5445 ( 
.A(n_4645),
.Y(n_5445)
);

AND2x4_ASAP7_75t_L g5446 ( 
.A(n_4206),
.B(n_3973),
.Y(n_5446)
);

NAND2xp33_ASAP7_75t_L g5447 ( 
.A(n_4234),
.B(n_4258),
.Y(n_5447)
);

O2A1O1Ixp33_ASAP7_75t_L g5448 ( 
.A1(n_4316),
.A2(n_4351),
.B(n_4353),
.C(n_4321),
.Y(n_5448)
);

BUFx3_ASAP7_75t_L g5449 ( 
.A(n_4002),
.Y(n_5449)
);

AND2x2_ASAP7_75t_L g5450 ( 
.A(n_4355),
.B(n_3841),
.Y(n_5450)
);

OAI21xp5_ASAP7_75t_L g5451 ( 
.A1(n_4061),
.A2(n_4100),
.B(n_4555),
.Y(n_5451)
);

O2A1O1Ixp33_ASAP7_75t_L g5452 ( 
.A1(n_4316),
.A2(n_4351),
.B(n_4353),
.C(n_4321),
.Y(n_5452)
);

INVx1_ASAP7_75t_SL g5453 ( 
.A(n_3989),
.Y(n_5453)
);

NAND2xp5_ASAP7_75t_L g5454 ( 
.A(n_4561),
.B(n_4510),
.Y(n_5454)
);

NOR2xp33_ASAP7_75t_L g5455 ( 
.A(n_4356),
.B(n_4357),
.Y(n_5455)
);

AOI21xp5_ASAP7_75t_L g5456 ( 
.A1(n_3938),
.A2(n_4001),
.B(n_3944),
.Y(n_5456)
);

INVx4_ASAP7_75t_L g5457 ( 
.A(n_4517),
.Y(n_5457)
);

NAND2xp5_ASAP7_75t_L g5458 ( 
.A(n_4561),
.B(n_4521),
.Y(n_5458)
);

AND2x2_ASAP7_75t_L g5459 ( 
.A(n_3841),
.B(n_3845),
.Y(n_5459)
);

NOR2xp33_ASAP7_75t_L g5460 ( 
.A(n_4356),
.B(n_4357),
.Y(n_5460)
);

AND2x4_ASAP7_75t_L g5461 ( 
.A(n_3973),
.B(n_4005),
.Y(n_5461)
);

O2A1O1Ixp5_ASAP7_75t_SL g5462 ( 
.A1(n_4645),
.A2(n_4654),
.B(n_4667),
.C(n_4651),
.Y(n_5462)
);

OAI22xp5_ASAP7_75t_L g5463 ( 
.A1(n_4222),
.A2(n_4302),
.B1(n_4397),
.B2(n_4106),
.Y(n_5463)
);

OAI22xp5_ASAP7_75t_L g5464 ( 
.A1(n_4302),
.A2(n_4397),
.B1(n_4106),
.B2(n_4621),
.Y(n_5464)
);

NAND2x1p5_ASAP7_75t_L g5465 ( 
.A(n_3865),
.B(n_3937),
.Y(n_5465)
);

NOR2x1_ASAP7_75t_R g5466 ( 
.A(n_4122),
.B(n_4234),
.Y(n_5466)
);

AOI21xp5_ASAP7_75t_L g5467 ( 
.A1(n_3938),
.A2(n_4001),
.B(n_3944),
.Y(n_5467)
);

BUFx2_ASAP7_75t_L g5468 ( 
.A(n_3843),
.Y(n_5468)
);

BUFx12f_ASAP7_75t_L g5469 ( 
.A(n_4122),
.Y(n_5469)
);

BUFx2_ASAP7_75t_L g5470 ( 
.A(n_3866),
.Y(n_5470)
);

NAND2xp5_ASAP7_75t_L g5471 ( 
.A(n_4525),
.B(n_4526),
.Y(n_5471)
);

A2O1A1Ixp33_ASAP7_75t_L g5472 ( 
.A1(n_4588),
.A2(n_4605),
.B(n_4293),
.C(n_4290),
.Y(n_5472)
);

AND2x4_ASAP7_75t_L g5473 ( 
.A(n_3973),
.B(n_4005),
.Y(n_5473)
);

NAND2x1p5_ASAP7_75t_L g5474 ( 
.A(n_3865),
.B(n_3937),
.Y(n_5474)
);

HB1xp67_ASAP7_75t_L g5475 ( 
.A(n_4639),
.Y(n_5475)
);

AND2x2_ASAP7_75t_SL g5476 ( 
.A(n_4211),
.B(n_4214),
.Y(n_5476)
);

BUFx12f_ASAP7_75t_L g5477 ( 
.A(n_4122),
.Y(n_5477)
);

NOR4xp25_ASAP7_75t_L g5478 ( 
.A(n_4619),
.B(n_3989),
.C(n_4650),
.D(n_4367),
.Y(n_5478)
);

AND2x4_ASAP7_75t_L g5479 ( 
.A(n_3973),
.B(n_4005),
.Y(n_5479)
);

AOI21xp5_ASAP7_75t_L g5480 ( 
.A1(n_3938),
.A2(n_4001),
.B(n_3944),
.Y(n_5480)
);

AOI21xp5_ASAP7_75t_L g5481 ( 
.A1(n_3938),
.A2(n_4001),
.B(n_3944),
.Y(n_5481)
);

AND2x2_ASAP7_75t_L g5482 ( 
.A(n_3841),
.B(n_3845),
.Y(n_5482)
);

AOI22xp5_ASAP7_75t_L g5483 ( 
.A1(n_4615),
.A2(n_4627),
.B1(n_4623),
.B2(n_4122),
.Y(n_5483)
);

OR2x6_ASAP7_75t_L g5484 ( 
.A(n_4090),
.B(n_3856),
.Y(n_5484)
);

AOI21xp5_ASAP7_75t_L g5485 ( 
.A1(n_3938),
.A2(n_4001),
.B(n_3944),
.Y(n_5485)
);

HB1xp67_ASAP7_75t_L g5486 ( 
.A(n_4643),
.Y(n_5486)
);

BUFx2_ASAP7_75t_L g5487 ( 
.A(n_3866),
.Y(n_5487)
);

AND2x4_ASAP7_75t_L g5488 ( 
.A(n_4005),
.B(n_4020),
.Y(n_5488)
);

OR2x6_ASAP7_75t_L g5489 ( 
.A(n_3856),
.B(n_3886),
.Y(n_5489)
);

AOI22xp33_ASAP7_75t_L g5490 ( 
.A1(n_4052),
.A2(n_4485),
.B1(n_4238),
.B2(n_4367),
.Y(n_5490)
);

AOI21xp5_ASAP7_75t_L g5491 ( 
.A1(n_4038),
.A2(n_4117),
.B(n_4097),
.Y(n_5491)
);

AOI21xp5_ASAP7_75t_L g5492 ( 
.A1(n_4038),
.A2(n_4117),
.B(n_4097),
.Y(n_5492)
);

AND2x4_ASAP7_75t_L g5493 ( 
.A(n_4005),
.B(n_4020),
.Y(n_5493)
);

NOR2xp33_ASAP7_75t_L g5494 ( 
.A(n_4359),
.B(n_4361),
.Y(n_5494)
);

AOI21xp5_ASAP7_75t_L g5495 ( 
.A1(n_4038),
.A2(n_4117),
.B(n_4097),
.Y(n_5495)
);

NOR2xp33_ASAP7_75t_L g5496 ( 
.A(n_4359),
.B(n_4361),
.Y(n_5496)
);

O2A1O1Ixp33_ASAP7_75t_L g5497 ( 
.A1(n_4364),
.A2(n_4370),
.B(n_4373),
.C(n_4369),
.Y(n_5497)
);

NAND2x1p5_ASAP7_75t_L g5498 ( 
.A(n_3865),
.B(n_3937),
.Y(n_5498)
);

AND2x2_ASAP7_75t_L g5499 ( 
.A(n_3845),
.B(n_3867),
.Y(n_5499)
);

O2A1O1Ixp33_ASAP7_75t_L g5500 ( 
.A1(n_4364),
.A2(n_4370),
.B(n_4373),
.C(n_4369),
.Y(n_5500)
);

NAND2x2_ASAP7_75t_L g5501 ( 
.A(n_3933),
.B(n_4202),
.Y(n_5501)
);

NAND2xp5_ASAP7_75t_L g5502 ( 
.A(n_4531),
.B(n_4536),
.Y(n_5502)
);

AND2x2_ASAP7_75t_L g5503 ( 
.A(n_3867),
.B(n_3902),
.Y(n_5503)
);

BUFx2_ASAP7_75t_L g5504 ( 
.A(n_3866),
.Y(n_5504)
);

A2O1A1Ixp33_ASAP7_75t_L g5505 ( 
.A1(n_4588),
.A2(n_4605),
.B(n_4293),
.C(n_4290),
.Y(n_5505)
);

OA21x2_ASAP7_75t_L g5506 ( 
.A1(n_4651),
.A2(n_4667),
.B(n_4582),
.Y(n_5506)
);

AOI21xp5_ASAP7_75t_L g5507 ( 
.A1(n_4038),
.A2(n_4117),
.B(n_4097),
.Y(n_5507)
);

BUFx3_ASAP7_75t_L g5508 ( 
.A(n_4002),
.Y(n_5508)
);

BUFx2_ASAP7_75t_L g5509 ( 
.A(n_3901),
.Y(n_5509)
);

AOI21xp5_ASAP7_75t_L g5510 ( 
.A1(n_4038),
.A2(n_4117),
.B(n_4097),
.Y(n_5510)
);

HB1xp67_ASAP7_75t_L g5511 ( 
.A(n_4643),
.Y(n_5511)
);

BUFx2_ASAP7_75t_L g5512 ( 
.A(n_3901),
.Y(n_5512)
);

HB1xp67_ASAP7_75t_L g5513 ( 
.A(n_4643),
.Y(n_5513)
);

A2O1A1Ixp33_ASAP7_75t_L g5514 ( 
.A1(n_4605),
.A2(n_4293),
.B(n_4290),
.C(n_4491),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_3982),
.Y(n_5515)
);

AOI222xp33_ASAP7_75t_L g5516 ( 
.A1(n_3941),
.A2(n_4619),
.B1(n_4150),
.B2(n_4618),
.C1(n_4640),
.C2(n_4630),
.Y(n_5516)
);

A2O1A1Ixp33_ASAP7_75t_L g5517 ( 
.A1(n_4605),
.A2(n_4293),
.B(n_4290),
.C(n_4491),
.Y(n_5517)
);

INVx2_ASAP7_75t_SL g5518 ( 
.A(n_4088),
.Y(n_5518)
);

INVx1_ASAP7_75t_L g5519 ( 
.A(n_3984),
.Y(n_5519)
);

AOI22xp33_ASAP7_75t_L g5520 ( 
.A1(n_4052),
.A2(n_4485),
.B1(n_4238),
.B2(n_4367),
.Y(n_5520)
);

HB1xp67_ASAP7_75t_L g5521 ( 
.A(n_4649),
.Y(n_5521)
);

OAI22xp5_ASAP7_75t_L g5522 ( 
.A1(n_4650),
.A2(n_4185),
.B1(n_4158),
.B2(n_4151),
.Y(n_5522)
);

AND2x2_ASAP7_75t_L g5523 ( 
.A(n_3867),
.B(n_3902),
.Y(n_5523)
);

AOI22xp5_ASAP7_75t_L g5524 ( 
.A1(n_4343),
.A2(n_4566),
.B1(n_4238),
.B2(n_4485),
.Y(n_5524)
);

NOR2xp33_ASAP7_75t_SL g5525 ( 
.A(n_4002),
.B(n_4232),
.Y(n_5525)
);

AND2x4_ASAP7_75t_L g5526 ( 
.A(n_4005),
.B(n_4020),
.Y(n_5526)
);

BUFx12f_ASAP7_75t_L g5527 ( 
.A(n_4258),
.Y(n_5527)
);

INVx5_ASAP7_75t_L g5528 ( 
.A(n_4052),
.Y(n_5528)
);

O2A1O1Ixp33_ASAP7_75t_L g5529 ( 
.A1(n_4374),
.A2(n_4377),
.B(n_4380),
.C(n_4378),
.Y(n_5529)
);

AND2x2_ASAP7_75t_L g5530 ( 
.A(n_3902),
.B(n_4059),
.Y(n_5530)
);

NOR2xp33_ASAP7_75t_SL g5531 ( 
.A(n_4232),
.B(n_4326),
.Y(n_5531)
);

A2O1A1Ixp33_ASAP7_75t_L g5532 ( 
.A1(n_4290),
.A2(n_4293),
.B(n_4343),
.C(n_3937),
.Y(n_5532)
);

OAI22xp5_ASAP7_75t_L g5533 ( 
.A1(n_4185),
.A2(n_4158),
.B1(n_4309),
.B2(n_4151),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_3984),
.Y(n_5534)
);

AOI21xp5_ASAP7_75t_L g5535 ( 
.A1(n_4151),
.A2(n_4309),
.B(n_4158),
.Y(n_5535)
);

O2A1O1Ixp33_ASAP7_75t_L g5536 ( 
.A1(n_4374),
.A2(n_4377),
.B(n_4380),
.C(n_4378),
.Y(n_5536)
);

NAND2xp5_ASAP7_75t_L g5537 ( 
.A(n_4536),
.B(n_4537),
.Y(n_5537)
);

NAND2xp5_ASAP7_75t_SL g5538 ( 
.A(n_4653),
.B(n_4068),
.Y(n_5538)
);

INVx1_ASAP7_75t_L g5539 ( 
.A(n_3985),
.Y(n_5539)
);

BUFx2_ASAP7_75t_L g5540 ( 
.A(n_3901),
.Y(n_5540)
);

CKINVDCx8_ASAP7_75t_R g5541 ( 
.A(n_4486),
.Y(n_5541)
);

AOI22xp33_ASAP7_75t_L g5542 ( 
.A1(n_4052),
.A2(n_4485),
.B1(n_4238),
.B2(n_4343),
.Y(n_5542)
);

NOR2x1_ASAP7_75t_SL g5543 ( 
.A(n_5434),
.B(n_4549),
.Y(n_5543)
);

NAND2xp5_ASAP7_75t_L g5544 ( 
.A(n_5299),
.B(n_4537),
.Y(n_5544)
);

AND2x4_ASAP7_75t_L g5545 ( 
.A(n_4970),
.B(n_4293),
.Y(n_5545)
);

AND2x4_ASAP7_75t_L g5546 ( 
.A(n_4970),
.B(n_4020),
.Y(n_5546)
);

NAND2xp5_ASAP7_75t_SL g5547 ( 
.A(n_5226),
.B(n_4184),
.Y(n_5547)
);

BUFx12f_ASAP7_75t_L g5548 ( 
.A(n_5301),
.Y(n_5548)
);

BUFx2_ASAP7_75t_L g5549 ( 
.A(n_5278),
.Y(n_5549)
);

NAND2x1p5_ASAP7_75t_L g5550 ( 
.A(n_5210),
.B(n_3865),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_5204),
.Y(n_5551)
);

OAI21x1_ASAP7_75t_L g5552 ( 
.A1(n_4746),
.A2(n_4575),
.B(n_4278),
.Y(n_5552)
);

INVx2_ASAP7_75t_L g5553 ( 
.A(n_4690),
.Y(n_5553)
);

AOI22xp5_ASAP7_75t_L g5554 ( 
.A1(n_5103),
.A2(n_4238),
.B1(n_4485),
.B2(n_4052),
.Y(n_5554)
);

INVx2_ASAP7_75t_L g5555 ( 
.A(n_4690),
.Y(n_5555)
);

AO21x2_ASAP7_75t_L g5556 ( 
.A1(n_4984),
.A2(n_4654),
.B(n_4582),
.Y(n_5556)
);

NAND2xp5_ASAP7_75t_L g5557 ( 
.A(n_5299),
.B(n_4548),
.Y(n_5557)
);

INVx3_ASAP7_75t_L g5558 ( 
.A(n_5121),
.Y(n_5558)
);

AOI22xp33_ASAP7_75t_L g5559 ( 
.A1(n_5103),
.A2(n_4485),
.B1(n_4238),
.B2(n_4549),
.Y(n_5559)
);

NAND2xp5_ASAP7_75t_L g5560 ( 
.A(n_5309),
.B(n_5332),
.Y(n_5560)
);

INVx3_ASAP7_75t_L g5561 ( 
.A(n_5121),
.Y(n_5561)
);

INVx2_ASAP7_75t_L g5562 ( 
.A(n_4690),
.Y(n_5562)
);

A2O1A1Ixp33_ASAP7_75t_L g5563 ( 
.A1(n_4871),
.A2(n_4214),
.B(n_4211),
.C(n_3937),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_5204),
.Y(n_5564)
);

INVx3_ASAP7_75t_L g5565 ( 
.A(n_5121),
.Y(n_5565)
);

BUFx4_ASAP7_75t_SL g5566 ( 
.A(n_5301),
.Y(n_5566)
);

INVx2_ASAP7_75t_L g5567 ( 
.A(n_4716),
.Y(n_5567)
);

INVxp67_ASAP7_75t_SL g5568 ( 
.A(n_5077),
.Y(n_5568)
);

BUFx2_ASAP7_75t_L g5569 ( 
.A(n_5278),
.Y(n_5569)
);

OR2x2_ASAP7_75t_SL g5570 ( 
.A(n_5163),
.B(n_4669),
.Y(n_5570)
);

BUFx6f_ASAP7_75t_L g5571 ( 
.A(n_4974),
.Y(n_5571)
);

AOI21x1_ASAP7_75t_L g5572 ( 
.A1(n_5117),
.A2(n_3998),
.B(n_4589),
.Y(n_5572)
);

AND2x6_ASAP7_75t_L g5573 ( 
.A(n_4758),
.B(n_4568),
.Y(n_5573)
);

HB1xp67_ASAP7_75t_L g5574 ( 
.A(n_4822),
.Y(n_5574)
);

INVxp67_ASAP7_75t_L g5575 ( 
.A(n_5125),
.Y(n_5575)
);

INVx2_ASAP7_75t_SL g5576 ( 
.A(n_4970),
.Y(n_5576)
);

AOI21xp33_ASAP7_75t_L g5577 ( 
.A1(n_4871),
.A2(n_4598),
.B(n_4548),
.Y(n_5577)
);

AOI21xp5_ASAP7_75t_L g5578 ( 
.A1(n_5185),
.A2(n_4572),
.B(n_4567),
.Y(n_5578)
);

AOI21xp5_ASAP7_75t_L g5579 ( 
.A1(n_5185),
.A2(n_5189),
.B(n_5174),
.Y(n_5579)
);

INVx3_ASAP7_75t_L g5580 ( 
.A(n_5121),
.Y(n_5580)
);

AOI21xp5_ASAP7_75t_L g5581 ( 
.A1(n_5189),
.A2(n_4572),
.B(n_4567),
.Y(n_5581)
);

INVx4_ASAP7_75t_L g5582 ( 
.A(n_5210),
.Y(n_5582)
);

CKINVDCx20_ASAP7_75t_R g5583 ( 
.A(n_4753),
.Y(n_5583)
);

CKINVDCx8_ASAP7_75t_R g5584 ( 
.A(n_5434),
.Y(n_5584)
);

NAND2xp5_ASAP7_75t_L g5585 ( 
.A(n_5309),
.B(n_4225),
.Y(n_5585)
);

AND2x2_ASAP7_75t_L g5586 ( 
.A(n_5150),
.B(n_3907),
.Y(n_5586)
);

HB1xp67_ASAP7_75t_L g5587 ( 
.A(n_4822),
.Y(n_5587)
);

AOI22xp33_ASAP7_75t_L g5588 ( 
.A1(n_5073),
.A2(n_4485),
.B1(n_4238),
.B2(n_4549),
.Y(n_5588)
);

CKINVDCx16_ASAP7_75t_R g5589 ( 
.A(n_5134),
.Y(n_5589)
);

INVx2_ASAP7_75t_L g5590 ( 
.A(n_4716),
.Y(n_5590)
);

BUFx6f_ASAP7_75t_L g5591 ( 
.A(n_4974),
.Y(n_5591)
);

NOR2x1_ASAP7_75t_SL g5592 ( 
.A(n_4739),
.B(n_4549),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_5243),
.Y(n_5593)
);

INVx2_ASAP7_75t_L g5594 ( 
.A(n_4716),
.Y(n_5594)
);

NOR2xp33_ASAP7_75t_L g5595 ( 
.A(n_4732),
.B(n_4598),
.Y(n_5595)
);

AND2x4_ASAP7_75t_L g5596 ( 
.A(n_4970),
.B(n_4020),
.Y(n_5596)
);

AOI22xp33_ASAP7_75t_L g5597 ( 
.A1(n_5073),
.A2(n_4485),
.B1(n_4238),
.B2(n_4549),
.Y(n_5597)
);

INVx5_ASAP7_75t_L g5598 ( 
.A(n_5058),
.Y(n_5598)
);

AND2x2_ASAP7_75t_SL g5599 ( 
.A(n_5178),
.B(n_4211),
.Y(n_5599)
);

NOR2xp33_ASAP7_75t_L g5600 ( 
.A(n_4732),
.B(n_4669),
.Y(n_5600)
);

INVx2_ASAP7_75t_L g5601 ( 
.A(n_4718),
.Y(n_5601)
);

INVx1_ASAP7_75t_SL g5602 ( 
.A(n_4881),
.Y(n_5602)
);

NAND2xp5_ASAP7_75t_SL g5603 ( 
.A(n_5226),
.B(n_4184),
.Y(n_5603)
);

BUFx6f_ASAP7_75t_L g5604 ( 
.A(n_4974),
.Y(n_5604)
);

INVx2_ASAP7_75t_L g5605 ( 
.A(n_4718),
.Y(n_5605)
);

AND2x4_ASAP7_75t_L g5606 ( 
.A(n_4970),
.B(n_4044),
.Y(n_5606)
);

INVx2_ASAP7_75t_L g5607 ( 
.A(n_4718),
.Y(n_5607)
);

OAI22xp5_ASAP7_75t_L g5608 ( 
.A1(n_4814),
.A2(n_4656),
.B1(n_4231),
.B2(n_4253),
.Y(n_5608)
);

BUFx6f_ASAP7_75t_L g5609 ( 
.A(n_4974),
.Y(n_5609)
);

OAI22xp5_ASAP7_75t_L g5610 ( 
.A1(n_4814),
.A2(n_4656),
.B1(n_4231),
.B2(n_4253),
.Y(n_5610)
);

CKINVDCx5p33_ASAP7_75t_R g5611 ( 
.A(n_4889),
.Y(n_5611)
);

BUFx2_ASAP7_75t_L g5612 ( 
.A(n_5278),
.Y(n_5612)
);

A2O1A1Ixp33_ASAP7_75t_L g5613 ( 
.A1(n_5123),
.A2(n_4214),
.B(n_3937),
.C(n_3964),
.Y(n_5613)
);

BUFx6f_ASAP7_75t_L g5614 ( 
.A(n_4974),
.Y(n_5614)
);

CKINVDCx5p33_ASAP7_75t_R g5615 ( 
.A(n_4889),
.Y(n_5615)
);

NAND2xp5_ASAP7_75t_L g5616 ( 
.A(n_5332),
.B(n_4225),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_5243),
.Y(n_5617)
);

INVx2_ASAP7_75t_L g5618 ( 
.A(n_4726),
.Y(n_5618)
);

BUFx4_ASAP7_75t_SL g5619 ( 
.A(n_4753),
.Y(n_5619)
);

OAI21x1_ASAP7_75t_L g5620 ( 
.A1(n_4746),
.A2(n_4575),
.B(n_4278),
.Y(n_5620)
);

INVx1_ASAP7_75t_L g5621 ( 
.A(n_5290),
.Y(n_5621)
);

BUFx4f_ASAP7_75t_L g5622 ( 
.A(n_4862),
.Y(n_5622)
);

BUFx2_ASAP7_75t_L g5623 ( 
.A(n_5278),
.Y(n_5623)
);

A2O1A1Ixp33_ASAP7_75t_L g5624 ( 
.A1(n_5123),
.A2(n_3937),
.B(n_3964),
.C(n_3865),
.Y(n_5624)
);

AND2x2_ASAP7_75t_L g5625 ( 
.A(n_5150),
.B(n_3907),
.Y(n_5625)
);

OAI21xp33_ASAP7_75t_L g5626 ( 
.A1(n_5163),
.A2(n_4646),
.B(n_4642),
.Y(n_5626)
);

OAI22xp5_ASAP7_75t_SL g5627 ( 
.A1(n_5227),
.A2(n_4414),
.B1(n_4382),
.B2(n_4566),
.Y(n_5627)
);

BUFx12f_ASAP7_75t_L g5628 ( 
.A(n_5134),
.Y(n_5628)
);

CKINVDCx8_ASAP7_75t_R g5629 ( 
.A(n_4881),
.Y(n_5629)
);

INVx2_ASAP7_75t_SL g5630 ( 
.A(n_4975),
.Y(n_5630)
);

AOI22xp33_ASAP7_75t_L g5631 ( 
.A1(n_4942),
.A2(n_4485),
.B1(n_4238),
.B2(n_4549),
.Y(n_5631)
);

NOR2xp33_ASAP7_75t_L g5632 ( 
.A(n_4839),
.B(n_5136),
.Y(n_5632)
);

INVx1_ASAP7_75t_L g5633 ( 
.A(n_5290),
.Y(n_5633)
);

HB1xp67_ASAP7_75t_L g5634 ( 
.A(n_4846),
.Y(n_5634)
);

BUFx6f_ASAP7_75t_L g5635 ( 
.A(n_4974),
.Y(n_5635)
);

AND2x4_ASAP7_75t_L g5636 ( 
.A(n_4975),
.B(n_5033),
.Y(n_5636)
);

BUFx2_ASAP7_75t_L g5637 ( 
.A(n_5278),
.Y(n_5637)
);

NAND2x2_ASAP7_75t_L g5638 ( 
.A(n_4686),
.B(n_4505),
.Y(n_5638)
);

BUFx6f_ASAP7_75t_L g5639 ( 
.A(n_4974),
.Y(n_5639)
);

NAND2xp5_ASAP7_75t_L g5640 ( 
.A(n_5334),
.B(n_4225),
.Y(n_5640)
);

BUFx3_ASAP7_75t_L g5641 ( 
.A(n_4975),
.Y(n_5641)
);

BUFx3_ASAP7_75t_L g5642 ( 
.A(n_4975),
.Y(n_5642)
);

NAND2xp5_ASAP7_75t_L g5643 ( 
.A(n_5334),
.B(n_4228),
.Y(n_5643)
);

INVx1_ASAP7_75t_L g5644 ( 
.A(n_5294),
.Y(n_5644)
);

OAI22xp5_ASAP7_75t_L g5645 ( 
.A1(n_4942),
.A2(n_4241),
.B1(n_4257),
.B2(n_4253),
.Y(n_5645)
);

BUFx2_ASAP7_75t_L g5646 ( 
.A(n_5278),
.Y(n_5646)
);

AND2x2_ASAP7_75t_L g5647 ( 
.A(n_5133),
.B(n_3942),
.Y(n_5647)
);

A2O1A1Ixp33_ASAP7_75t_L g5648 ( 
.A1(n_5135),
.A2(n_3937),
.B(n_3964),
.C(n_3865),
.Y(n_5648)
);

AOI21xp5_ASAP7_75t_L g5649 ( 
.A1(n_4985),
.A2(n_4583),
.B(n_4577),
.Y(n_5649)
);

BUFx3_ASAP7_75t_L g5650 ( 
.A(n_4975),
.Y(n_5650)
);

OAI221xp5_ASAP7_75t_L g5651 ( 
.A1(n_5193),
.A2(n_4653),
.B1(n_4652),
.B2(n_4649),
.C(n_4642),
.Y(n_5651)
);

INVx2_ASAP7_75t_L g5652 ( 
.A(n_4726),
.Y(n_5652)
);

INVx2_ASAP7_75t_L g5653 ( 
.A(n_4726),
.Y(n_5653)
);

OR2x2_ASAP7_75t_L g5654 ( 
.A(n_5233),
.B(n_4646),
.Y(n_5654)
);

INVx1_ASAP7_75t_L g5655 ( 
.A(n_5294),
.Y(n_5655)
);

OAI22xp5_ASAP7_75t_L g5656 ( 
.A1(n_5087),
.A2(n_4241),
.B1(n_4342),
.B2(n_4257),
.Y(n_5656)
);

INVx2_ASAP7_75t_SL g5657 ( 
.A(n_4975),
.Y(n_5657)
);

AOI22xp33_ASAP7_75t_L g5658 ( 
.A1(n_5139),
.A2(n_4485),
.B1(n_4238),
.B2(n_4630),
.Y(n_5658)
);

BUFx4_ASAP7_75t_SL g5659 ( 
.A(n_4866),
.Y(n_5659)
);

OAI22xp33_ASAP7_75t_L g5660 ( 
.A1(n_5139),
.A2(n_4123),
.B1(n_4455),
.B2(n_4098),
.Y(n_5660)
);

INVx1_ASAP7_75t_L g5661 ( 
.A(n_5399),
.Y(n_5661)
);

OR2x2_ASAP7_75t_L g5662 ( 
.A(n_5233),
.B(n_4154),
.Y(n_5662)
);

BUFx2_ASAP7_75t_L g5663 ( 
.A(n_5278),
.Y(n_5663)
);

OAI22xp5_ASAP7_75t_L g5664 ( 
.A1(n_5087),
.A2(n_5110),
.B1(n_5159),
.B2(n_5136),
.Y(n_5664)
);

NAND2xp5_ASAP7_75t_L g5665 ( 
.A(n_5086),
.B(n_4228),
.Y(n_5665)
);

BUFx3_ASAP7_75t_L g5666 ( 
.A(n_5033),
.Y(n_5666)
);

BUFx6f_ASAP7_75t_L g5667 ( 
.A(n_4974),
.Y(n_5667)
);

AOI22xp33_ASAP7_75t_L g5668 ( 
.A1(n_5151),
.A2(n_4485),
.B1(n_4238),
.B2(n_4640),
.Y(n_5668)
);

INVx1_ASAP7_75t_L g5669 ( 
.A(n_5399),
.Y(n_5669)
);

AND2x4_ASAP7_75t_L g5670 ( 
.A(n_5033),
.B(n_5262),
.Y(n_5670)
);

NOR2xp67_ASAP7_75t_SL g5671 ( 
.A(n_5084),
.B(n_4098),
.Y(n_5671)
);

AO21x1_ASAP7_75t_L g5672 ( 
.A1(n_5130),
.A2(n_4385),
.B(n_4384),
.Y(n_5672)
);

INVx1_ASAP7_75t_SL g5673 ( 
.A(n_4710),
.Y(n_5673)
);

AOI22xp33_ASAP7_75t_L g5674 ( 
.A1(n_5151),
.A2(n_3856),
.B1(n_4168),
.B2(n_3886),
.Y(n_5674)
);

HB1xp67_ASAP7_75t_L g5675 ( 
.A(n_4846),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5475),
.Y(n_5676)
);

AND2x6_ASAP7_75t_L g5677 ( 
.A(n_4758),
.B(n_4568),
.Y(n_5677)
);

NAND2xp5_ASAP7_75t_L g5678 ( 
.A(n_5086),
.B(n_4228),
.Y(n_5678)
);

NOR2xp33_ASAP7_75t_L g5679 ( 
.A(n_4839),
.B(n_4384),
.Y(n_5679)
);

INVx1_ASAP7_75t_SL g5680 ( 
.A(n_4710),
.Y(n_5680)
);

NAND2xp5_ASAP7_75t_L g5681 ( 
.A(n_5264),
.B(n_4199),
.Y(n_5681)
);

OAI22xp5_ASAP7_75t_L g5682 ( 
.A1(n_5110),
.A2(n_5159),
.B1(n_5156),
.B2(n_5084),
.Y(n_5682)
);

INVx3_ASAP7_75t_L g5683 ( 
.A(n_4987),
.Y(n_5683)
);

AOI21xp5_ASAP7_75t_L g5684 ( 
.A1(n_4985),
.A2(n_4557),
.B(n_4404),
.Y(n_5684)
);

NAND2xp5_ASAP7_75t_L g5685 ( 
.A(n_5264),
.B(n_4199),
.Y(n_5685)
);

INVx3_ASAP7_75t_L g5686 ( 
.A(n_4987),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5475),
.Y(n_5687)
);

AOI22xp33_ASAP7_75t_L g5688 ( 
.A1(n_5165),
.A2(n_3856),
.B1(n_4168),
.B2(n_3886),
.Y(n_5688)
);

NAND2xp5_ASAP7_75t_L g5689 ( 
.A(n_5231),
.B(n_4199),
.Y(n_5689)
);

NAND2xp5_ASAP7_75t_L g5690 ( 
.A(n_5231),
.B(n_4215),
.Y(n_5690)
);

BUFx6f_ASAP7_75t_L g5691 ( 
.A(n_4987),
.Y(n_5691)
);

BUFx2_ASAP7_75t_L g5692 ( 
.A(n_5278),
.Y(n_5692)
);

NOR2xp33_ASAP7_75t_L g5693 ( 
.A(n_5104),
.B(n_4385),
.Y(n_5693)
);

INVx4_ASAP7_75t_L g5694 ( 
.A(n_5210),
.Y(n_5694)
);

AOI22xp5_ASAP7_75t_L g5695 ( 
.A1(n_5167),
.A2(n_4568),
.B1(n_4534),
.B2(n_4487),
.Y(n_5695)
);

INVx2_ASAP7_75t_L g5696 ( 
.A(n_4747),
.Y(n_5696)
);

HB1xp67_ASAP7_75t_L g5697 ( 
.A(n_4868),
.Y(n_5697)
);

CKINVDCx16_ASAP7_75t_R g5698 ( 
.A(n_5134),
.Y(n_5698)
);

BUFx3_ASAP7_75t_L g5699 ( 
.A(n_5033),
.Y(n_5699)
);

INVx2_ASAP7_75t_L g5700 ( 
.A(n_4747),
.Y(n_5700)
);

INVx3_ASAP7_75t_L g5701 ( 
.A(n_4987),
.Y(n_5701)
);

NAND2xp5_ASAP7_75t_L g5702 ( 
.A(n_5141),
.B(n_4215),
.Y(n_5702)
);

AOI21xp5_ASAP7_75t_L g5703 ( 
.A1(n_5135),
.A2(n_4557),
.B(n_4404),
.Y(n_5703)
);

AND2x4_ASAP7_75t_L g5704 ( 
.A(n_5033),
.B(n_4443),
.Y(n_5704)
);

NOR2xp33_ASAP7_75t_L g5705 ( 
.A(n_5104),
.B(n_5120),
.Y(n_5705)
);

BUFx3_ASAP7_75t_L g5706 ( 
.A(n_5058),
.Y(n_5706)
);

AND2x2_ASAP7_75t_L g5707 ( 
.A(n_5137),
.B(n_4059),
.Y(n_5707)
);

NAND2xp5_ASAP7_75t_SL g5708 ( 
.A(n_5210),
.B(n_5153),
.Y(n_5708)
);

INVx1_ASAP7_75t_L g5709 ( 
.A(n_5486),
.Y(n_5709)
);

OAI22xp5_ASAP7_75t_L g5710 ( 
.A1(n_5156),
.A2(n_4241),
.B1(n_4342),
.B2(n_4257),
.Y(n_5710)
);

AOI21xp5_ASAP7_75t_L g5711 ( 
.A1(n_5166),
.A2(n_4562),
.B(n_4391),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_5486),
.Y(n_5712)
);

BUFx2_ASAP7_75t_L g5713 ( 
.A(n_5102),
.Y(n_5713)
);

AOI22xp33_ASAP7_75t_L g5714 ( 
.A1(n_5165),
.A2(n_3856),
.B1(n_4168),
.B2(n_3886),
.Y(n_5714)
);

INVx2_ASAP7_75t_SL g5715 ( 
.A(n_5058),
.Y(n_5715)
);

CKINVDCx14_ASAP7_75t_R g5716 ( 
.A(n_4784),
.Y(n_5716)
);

AND2x4_ASAP7_75t_L g5717 ( 
.A(n_5262),
.B(n_4064),
.Y(n_5717)
);

AND2x2_ASAP7_75t_L g5718 ( 
.A(n_5137),
.B(n_4059),
.Y(n_5718)
);

OR2x6_ASAP7_75t_L g5719 ( 
.A(n_4923),
.B(n_4152),
.Y(n_5719)
);

INVx6_ASAP7_75t_SL g5720 ( 
.A(n_5489),
.Y(n_5720)
);

INVx1_ASAP7_75t_SL g5721 ( 
.A(n_4936),
.Y(n_5721)
);

NAND2xp5_ASAP7_75t_L g5722 ( 
.A(n_5141),
.B(n_4215),
.Y(n_5722)
);

NOR2xp33_ASAP7_75t_SL g5723 ( 
.A(n_5071),
.B(n_4232),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_5511),
.Y(n_5724)
);

NAND2xp5_ASAP7_75t_L g5725 ( 
.A(n_5207),
.B(n_4389),
.Y(n_5725)
);

HB1xp67_ASAP7_75t_L g5726 ( 
.A(n_4868),
.Y(n_5726)
);

INVx3_ASAP7_75t_L g5727 ( 
.A(n_4987),
.Y(n_5727)
);

INVx3_ASAP7_75t_L g5728 ( 
.A(n_4987),
.Y(n_5728)
);

INVx4_ASAP7_75t_L g5729 ( 
.A(n_5210),
.Y(n_5729)
);

BUFx2_ASAP7_75t_L g5730 ( 
.A(n_5102),
.Y(n_5730)
);

INVx2_ASAP7_75t_L g5731 ( 
.A(n_4747),
.Y(n_5731)
);

NAND2xp5_ASAP7_75t_SL g5732 ( 
.A(n_5153),
.B(n_4184),
.Y(n_5732)
);

AND2x2_ASAP7_75t_L g5733 ( 
.A(n_5137),
.B(n_4066),
.Y(n_5733)
);

INVx1_ASAP7_75t_L g5734 ( 
.A(n_5511),
.Y(n_5734)
);

NAND2xp5_ASAP7_75t_L g5735 ( 
.A(n_5207),
.B(n_4389),
.Y(n_5735)
);

OAI22xp5_ASAP7_75t_SL g5736 ( 
.A1(n_5227),
.A2(n_4382),
.B1(n_4414),
.B2(n_4342),
.Y(n_5736)
);

INVx2_ASAP7_75t_L g5737 ( 
.A(n_4759),
.Y(n_5737)
);

OAI22x1_ASAP7_75t_L g5738 ( 
.A1(n_5175),
.A2(n_4575),
.B1(n_4449),
.B2(n_4450),
.Y(n_5738)
);

INVxp67_ASAP7_75t_L g5739 ( 
.A(n_5125),
.Y(n_5739)
);

BUFx6f_ASAP7_75t_L g5740 ( 
.A(n_4987),
.Y(n_5740)
);

AOI22xp33_ASAP7_75t_L g5741 ( 
.A1(n_5167),
.A2(n_4168),
.B1(n_3886),
.B2(n_4487),
.Y(n_5741)
);

INVxp67_ASAP7_75t_L g5742 ( 
.A(n_5125),
.Y(n_5742)
);

INVx2_ASAP7_75t_L g5743 ( 
.A(n_4759),
.Y(n_5743)
);

INVx2_ASAP7_75t_L g5744 ( 
.A(n_4759),
.Y(n_5744)
);

NAND2xp5_ASAP7_75t_L g5745 ( 
.A(n_4691),
.B(n_4391),
.Y(n_5745)
);

BUFx4_ASAP7_75t_SL g5746 ( 
.A(n_4866),
.Y(n_5746)
);

BUFx3_ASAP7_75t_L g5747 ( 
.A(n_5058),
.Y(n_5747)
);

CKINVDCx11_ASAP7_75t_R g5748 ( 
.A(n_4940),
.Y(n_5748)
);

INVx2_ASAP7_75t_L g5749 ( 
.A(n_4768),
.Y(n_5749)
);

AOI22xp5_ASAP7_75t_L g5750 ( 
.A1(n_5091),
.A2(n_4534),
.B1(n_4487),
.B2(n_4478),
.Y(n_5750)
);

AOI22xp5_ASAP7_75t_L g5751 ( 
.A1(n_5091),
.A2(n_4534),
.B1(n_4478),
.B2(n_4453),
.Y(n_5751)
);

BUFx3_ASAP7_75t_L g5752 ( 
.A(n_5058),
.Y(n_5752)
);

BUFx3_ASAP7_75t_L g5753 ( 
.A(n_5058),
.Y(n_5753)
);

NOR2xp33_ASAP7_75t_R g5754 ( 
.A(n_4784),
.B(n_4232),
.Y(n_5754)
);

HB1xp67_ASAP7_75t_L g5755 ( 
.A(n_4879),
.Y(n_5755)
);

CKINVDCx11_ASAP7_75t_R g5756 ( 
.A(n_4940),
.Y(n_5756)
);

INVx1_ASAP7_75t_SL g5757 ( 
.A(n_4936),
.Y(n_5757)
);

CKINVDCx5p33_ASAP7_75t_R g5758 ( 
.A(n_5094),
.Y(n_5758)
);

INVxp67_ASAP7_75t_L g5759 ( 
.A(n_4684),
.Y(n_5759)
);

AND3x1_ASAP7_75t_L g5760 ( 
.A(n_5120),
.B(n_4505),
.C(n_4453),
.Y(n_5760)
);

INVx1_ASAP7_75t_L g5761 ( 
.A(n_5513),
.Y(n_5761)
);

BUFx3_ASAP7_75t_L g5762 ( 
.A(n_5058),
.Y(n_5762)
);

INVx2_ASAP7_75t_L g5763 ( 
.A(n_4768),
.Y(n_5763)
);

BUFx3_ASAP7_75t_L g5764 ( 
.A(n_5058),
.Y(n_5764)
);

INVx6_ASAP7_75t_SL g5765 ( 
.A(n_5489),
.Y(n_5765)
);

NAND2xp5_ASAP7_75t_L g5766 ( 
.A(n_4691),
.B(n_4395),
.Y(n_5766)
);

INVx2_ASAP7_75t_L g5767 ( 
.A(n_4768),
.Y(n_5767)
);

AOI21xp33_ASAP7_75t_L g5768 ( 
.A1(n_5132),
.A2(n_4652),
.B(n_4649),
.Y(n_5768)
);

AND2x2_ASAP7_75t_L g5769 ( 
.A(n_5194),
.B(n_4066),
.Y(n_5769)
);

AOI21xp5_ASAP7_75t_L g5770 ( 
.A1(n_5166),
.A2(n_4984),
.B(n_5222),
.Y(n_5770)
);

BUFx3_ASAP7_75t_L g5771 ( 
.A(n_5149),
.Y(n_5771)
);

AND2x2_ASAP7_75t_L g5772 ( 
.A(n_5194),
.B(n_4066),
.Y(n_5772)
);

INVx1_ASAP7_75t_L g5773 ( 
.A(n_5513),
.Y(n_5773)
);

AND2x2_ASAP7_75t_L g5774 ( 
.A(n_5194),
.B(n_4126),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_5521),
.Y(n_5775)
);

INVx5_ASAP7_75t_L g5776 ( 
.A(n_5149),
.Y(n_5776)
);

OAI21x1_ASAP7_75t_L g5777 ( 
.A1(n_4746),
.A2(n_4575),
.B(n_4278),
.Y(n_5777)
);

BUFx2_ASAP7_75t_L g5778 ( 
.A(n_5102),
.Y(n_5778)
);

NAND2xp5_ASAP7_75t_L g5779 ( 
.A(n_4760),
.B(n_4395),
.Y(n_5779)
);

AND2x2_ASAP7_75t_L g5780 ( 
.A(n_5199),
.B(n_4126),
.Y(n_5780)
);

OR2x6_ASAP7_75t_L g5781 ( 
.A(n_4923),
.B(n_5283),
.Y(n_5781)
);

INVx2_ASAP7_75t_L g5782 ( 
.A(n_4799),
.Y(n_5782)
);

NAND3xp33_ASAP7_75t_L g5783 ( 
.A(n_5132),
.B(n_4652),
.C(n_4398),
.Y(n_5783)
);

NAND2xp5_ASAP7_75t_L g5784 ( 
.A(n_4760),
.B(n_4396),
.Y(n_5784)
);

AOI22xp33_ASAP7_75t_L g5785 ( 
.A1(n_5111),
.A2(n_4168),
.B1(n_3886),
.B2(n_4534),
.Y(n_5785)
);

INVx1_ASAP7_75t_L g5786 ( 
.A(n_5521),
.Y(n_5786)
);

OAI22xp5_ASAP7_75t_L g5787 ( 
.A1(n_5175),
.A2(n_4226),
.B1(n_4158),
.B2(n_4151),
.Y(n_5787)
);

BUFx2_ASAP7_75t_L g5788 ( 
.A(n_5102),
.Y(n_5788)
);

BUFx2_ASAP7_75t_L g5789 ( 
.A(n_5102),
.Y(n_5789)
);

INVxp67_ASAP7_75t_L g5790 ( 
.A(n_4684),
.Y(n_5790)
);

AOI22xp33_ASAP7_75t_L g5791 ( 
.A1(n_5111),
.A2(n_4168),
.B1(n_3886),
.B2(n_4534),
.Y(n_5791)
);

INVx8_ASAP7_75t_L g5792 ( 
.A(n_4923),
.Y(n_5792)
);

HB1xp67_ASAP7_75t_L g5793 ( 
.A(n_4879),
.Y(n_5793)
);

BUFx3_ASAP7_75t_L g5794 ( 
.A(n_5149),
.Y(n_5794)
);

INVx1_ASAP7_75t_L g5795 ( 
.A(n_4884),
.Y(n_5795)
);

INVx2_ASAP7_75t_L g5796 ( 
.A(n_4799),
.Y(n_5796)
);

INVx2_ASAP7_75t_SL g5797 ( 
.A(n_5149),
.Y(n_5797)
);

OR2x6_ASAP7_75t_L g5798 ( 
.A(n_4923),
.B(n_4152),
.Y(n_5798)
);

NAND2xp5_ASAP7_75t_L g5799 ( 
.A(n_5247),
.B(n_4396),
.Y(n_5799)
);

NAND2xp5_ASAP7_75t_L g5800 ( 
.A(n_5247),
.B(n_4398),
.Y(n_5800)
);

CKINVDCx8_ASAP7_75t_R g5801 ( 
.A(n_4852),
.Y(n_5801)
);

BUFx2_ASAP7_75t_L g5802 ( 
.A(n_5102),
.Y(n_5802)
);

INVx1_ASAP7_75t_L g5803 ( 
.A(n_4884),
.Y(n_5803)
);

AOI22xp5_ASAP7_75t_L g5804 ( 
.A1(n_5214),
.A2(n_4534),
.B1(n_4478),
.B2(n_4195),
.Y(n_5804)
);

AND2x2_ASAP7_75t_L g5805 ( 
.A(n_5199),
.B(n_4126),
.Y(n_5805)
);

NOR2xp33_ASAP7_75t_L g5806 ( 
.A(n_5183),
.B(n_4401),
.Y(n_5806)
);

NAND2xp5_ASAP7_75t_L g5807 ( 
.A(n_5269),
.B(n_4401),
.Y(n_5807)
);

NAND2xp5_ASAP7_75t_L g5808 ( 
.A(n_5269),
.B(n_4410),
.Y(n_5808)
);

AOI22xp33_ASAP7_75t_L g5809 ( 
.A1(n_5214),
.A2(n_5219),
.B1(n_5183),
.B2(n_4765),
.Y(n_5809)
);

CKINVDCx5p33_ASAP7_75t_R g5810 ( 
.A(n_5094),
.Y(n_5810)
);

INVx3_ASAP7_75t_L g5811 ( 
.A(n_4988),
.Y(n_5811)
);

HB1xp67_ASAP7_75t_L g5812 ( 
.A(n_4687),
.Y(n_5812)
);

INVx1_ASAP7_75t_L g5813 ( 
.A(n_5180),
.Y(n_5813)
);

CKINVDCx8_ASAP7_75t_R g5814 ( 
.A(n_4852),
.Y(n_5814)
);

BUFx2_ASAP7_75t_L g5815 ( 
.A(n_5102),
.Y(n_5815)
);

HB1xp67_ASAP7_75t_L g5816 ( 
.A(n_4687),
.Y(n_5816)
);

INVx2_ASAP7_75t_SL g5817 ( 
.A(n_5149),
.Y(n_5817)
);

OAI22xp33_ASAP7_75t_L g5818 ( 
.A1(n_5271),
.A2(n_4123),
.B1(n_4455),
.B2(n_4098),
.Y(n_5818)
);

INVx3_ASAP7_75t_L g5819 ( 
.A(n_4988),
.Y(n_5819)
);

BUFx3_ASAP7_75t_L g5820 ( 
.A(n_5149),
.Y(n_5820)
);

AND2x2_ASAP7_75t_L g5821 ( 
.A(n_5199),
.B(n_5272),
.Y(n_5821)
);

INVx4_ASAP7_75t_SL g5822 ( 
.A(n_5225),
.Y(n_5822)
);

BUFx12f_ASAP7_75t_L g5823 ( 
.A(n_4730),
.Y(n_5823)
);

NAND2xp5_ASAP7_75t_L g5824 ( 
.A(n_5302),
.B(n_4410),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_5180),
.Y(n_5825)
);

INVx3_ASAP7_75t_L g5826 ( 
.A(n_4988),
.Y(n_5826)
);

BUFx3_ASAP7_75t_L g5827 ( 
.A(n_5149),
.Y(n_5827)
);

NAND2xp5_ASAP7_75t_L g5828 ( 
.A(n_5302),
.B(n_4413),
.Y(n_5828)
);

INVx1_ASAP7_75t_L g5829 ( 
.A(n_5190),
.Y(n_5829)
);

NOR2xp33_ASAP7_75t_L g5830 ( 
.A(n_5236),
.B(n_4413),
.Y(n_5830)
);

BUFx8_ASAP7_75t_SL g5831 ( 
.A(n_5095),
.Y(n_5831)
);

NAND2xp5_ASAP7_75t_L g5832 ( 
.A(n_5019),
.B(n_4415),
.Y(n_5832)
);

CKINVDCx5p33_ASAP7_75t_R g5833 ( 
.A(n_5095),
.Y(n_5833)
);

INVx4_ASAP7_75t_L g5834 ( 
.A(n_4739),
.Y(n_5834)
);

NAND2x1p5_ASAP7_75t_L g5835 ( 
.A(n_4921),
.B(n_3865),
.Y(n_5835)
);

NOR2xp33_ASAP7_75t_L g5836 ( 
.A(n_5236),
.B(n_4415),
.Y(n_5836)
);

BUFx2_ASAP7_75t_L g5837 ( 
.A(n_5102),
.Y(n_5837)
);

INVx1_ASAP7_75t_L g5838 ( 
.A(n_5190),
.Y(n_5838)
);

AOI21xp5_ASAP7_75t_L g5839 ( 
.A1(n_5222),
.A2(n_4562),
.B(n_4417),
.Y(n_5839)
);

INVx3_ASAP7_75t_L g5840 ( 
.A(n_4988),
.Y(n_5840)
);

NAND2xp5_ASAP7_75t_L g5841 ( 
.A(n_5019),
.B(n_4416),
.Y(n_5841)
);

AOI21xp5_ASAP7_75t_L g5842 ( 
.A1(n_4861),
.A2(n_4417),
.B(n_4416),
.Y(n_5842)
);

NOR2xp67_ASAP7_75t_L g5843 ( 
.A(n_5417),
.B(n_4243),
.Y(n_5843)
);

BUFx3_ASAP7_75t_L g5844 ( 
.A(n_5149),
.Y(n_5844)
);

CKINVDCx5p33_ASAP7_75t_R g5845 ( 
.A(n_5170),
.Y(n_5845)
);

BUFx4_ASAP7_75t_SL g5846 ( 
.A(n_5441),
.Y(n_5846)
);

O2A1O1Ixp33_ASAP7_75t_L g5847 ( 
.A1(n_4712),
.A2(n_4421),
.B(n_4422),
.C(n_4419),
.Y(n_5847)
);

HB1xp67_ASAP7_75t_L g5848 ( 
.A(n_4703),
.Y(n_5848)
);

INVx2_ASAP7_75t_SL g5849 ( 
.A(n_5197),
.Y(n_5849)
);

INVx1_ASAP7_75t_SL g5850 ( 
.A(n_4973),
.Y(n_5850)
);

AND2x2_ASAP7_75t_L g5851 ( 
.A(n_5287),
.B(n_4088),
.Y(n_5851)
);

INVx4_ASAP7_75t_L g5852 ( 
.A(n_4739),
.Y(n_5852)
);

AOI21xp5_ASAP7_75t_L g5853 ( 
.A1(n_4861),
.A2(n_4421),
.B(n_4419),
.Y(n_5853)
);

INVx1_ASAP7_75t_L g5854 ( 
.A(n_5191),
.Y(n_5854)
);

INVx4_ASAP7_75t_L g5855 ( 
.A(n_4787),
.Y(n_5855)
);

AND2x2_ASAP7_75t_L g5856 ( 
.A(n_5287),
.B(n_4088),
.Y(n_5856)
);

O2A1O1Ixp33_ASAP7_75t_L g5857 ( 
.A1(n_4712),
.A2(n_4429),
.B(n_4436),
.C(n_4422),
.Y(n_5857)
);

AND2x4_ASAP7_75t_L g5858 ( 
.A(n_5352),
.B(n_5393),
.Y(n_5858)
);

CKINVDCx8_ASAP7_75t_R g5859 ( 
.A(n_5408),
.Y(n_5859)
);

BUFx3_ASAP7_75t_L g5860 ( 
.A(n_5197),
.Y(n_5860)
);

AND2x2_ASAP7_75t_SL g5861 ( 
.A(n_5178),
.B(n_3831),
.Y(n_5861)
);

AOI21xp5_ASAP7_75t_SL g5862 ( 
.A1(n_5193),
.A2(n_4243),
.B(n_4429),
.Y(n_5862)
);

OR2x6_ASAP7_75t_L g5863 ( 
.A(n_4923),
.B(n_4152),
.Y(n_5863)
);

AOI22xp33_ASAP7_75t_SL g5864 ( 
.A1(n_5219),
.A2(n_3937),
.B1(n_3964),
.B2(n_3865),
.Y(n_5864)
);

BUFx6f_ASAP7_75t_L g5865 ( 
.A(n_4988),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_5191),
.Y(n_5866)
);

CKINVDCx20_ASAP7_75t_R g5867 ( 
.A(n_5170),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5192),
.Y(n_5868)
);

BUFx3_ASAP7_75t_L g5869 ( 
.A(n_5197),
.Y(n_5869)
);

NOR2x1_ASAP7_75t_SL g5870 ( 
.A(n_4787),
.B(n_4152),
.Y(n_5870)
);

INVx3_ASAP7_75t_L g5871 ( 
.A(n_4991),
.Y(n_5871)
);

BUFx3_ASAP7_75t_L g5872 ( 
.A(n_5197),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5192),
.Y(n_5873)
);

AOI21xp5_ASAP7_75t_L g5874 ( 
.A1(n_4794),
.A2(n_4440),
.B(n_4436),
.Y(n_5874)
);

INVx8_ASAP7_75t_L g5875 ( 
.A(n_4923),
.Y(n_5875)
);

CKINVDCx8_ASAP7_75t_R g5876 ( 
.A(n_5408),
.Y(n_5876)
);

INVx1_ASAP7_75t_L g5877 ( 
.A(n_4679),
.Y(n_5877)
);

INVx5_ASAP7_75t_L g5878 ( 
.A(n_5197),
.Y(n_5878)
);

INVxp67_ASAP7_75t_SL g5879 ( 
.A(n_5077),
.Y(n_5879)
);

INVx5_ASAP7_75t_L g5880 ( 
.A(n_5197),
.Y(n_5880)
);

INVx1_ASAP7_75t_L g5881 ( 
.A(n_4679),
.Y(n_5881)
);

INVx5_ASAP7_75t_L g5882 ( 
.A(n_5197),
.Y(n_5882)
);

AOI22xp33_ASAP7_75t_L g5883 ( 
.A1(n_4765),
.A2(n_4168),
.B1(n_4449),
.B2(n_4443),
.Y(n_5883)
);

INVx5_ASAP7_75t_L g5884 ( 
.A(n_5197),
.Y(n_5884)
);

BUFx3_ASAP7_75t_L g5885 ( 
.A(n_5528),
.Y(n_5885)
);

BUFx3_ASAP7_75t_L g5886 ( 
.A(n_5528),
.Y(n_5886)
);

INVx1_ASAP7_75t_L g5887 ( 
.A(n_4682),
.Y(n_5887)
);

AOI22xp5_ASAP7_75t_L g5888 ( 
.A1(n_4887),
.A2(n_4209),
.B1(n_4254),
.B2(n_4195),
.Y(n_5888)
);

INVx2_ASAP7_75t_SL g5889 ( 
.A(n_5528),
.Y(n_5889)
);

HB1xp67_ASAP7_75t_L g5890 ( 
.A(n_4703),
.Y(n_5890)
);

BUFx4f_ASAP7_75t_L g5891 ( 
.A(n_4862),
.Y(n_5891)
);

OR2x2_ASAP7_75t_L g5892 ( 
.A(n_5478),
.B(n_4154),
.Y(n_5892)
);

INVx3_ASAP7_75t_L g5893 ( 
.A(n_4991),
.Y(n_5893)
);

AOI21xp5_ASAP7_75t_L g5894 ( 
.A1(n_4794),
.A2(n_4924),
.B(n_5291),
.Y(n_5894)
);

AOI22xp33_ASAP7_75t_L g5895 ( 
.A1(n_5130),
.A2(n_4449),
.B1(n_4450),
.B2(n_4443),
.Y(n_5895)
);

NAND2xp5_ASAP7_75t_L g5896 ( 
.A(n_5325),
.B(n_4440),
.Y(n_5896)
);

CKINVDCx5p33_ASAP7_75t_R g5897 ( 
.A(n_5338),
.Y(n_5897)
);

INVx1_ASAP7_75t_L g5898 ( 
.A(n_4682),
.Y(n_5898)
);

BUFx4_ASAP7_75t_SL g5899 ( 
.A(n_5441),
.Y(n_5899)
);

BUFx2_ASAP7_75t_L g5900 ( 
.A(n_5393),
.Y(n_5900)
);

INVx1_ASAP7_75t_L g5901 ( 
.A(n_4683),
.Y(n_5901)
);

BUFx2_ASAP7_75t_L g5902 ( 
.A(n_5393),
.Y(n_5902)
);

NAND2xp5_ASAP7_75t_L g5903 ( 
.A(n_5325),
.B(n_4445),
.Y(n_5903)
);

NAND2xp5_ASAP7_75t_L g5904 ( 
.A(n_5168),
.B(n_4445),
.Y(n_5904)
);

HB1xp67_ASAP7_75t_L g5905 ( 
.A(n_4770),
.Y(n_5905)
);

INVx1_ASAP7_75t_SL g5906 ( 
.A(n_4973),
.Y(n_5906)
);

BUFx12f_ASAP7_75t_L g5907 ( 
.A(n_4751),
.Y(n_5907)
);

NAND2xp5_ASAP7_75t_L g5908 ( 
.A(n_5168),
.B(n_4446),
.Y(n_5908)
);

BUFx2_ASAP7_75t_L g5909 ( 
.A(n_5393),
.Y(n_5909)
);

INVx4_ASAP7_75t_L g5910 ( 
.A(n_4787),
.Y(n_5910)
);

AND2x6_ASAP7_75t_L g5911 ( 
.A(n_4748),
.B(n_4195),
.Y(n_5911)
);

NAND2xp5_ASAP7_75t_L g5912 ( 
.A(n_5292),
.B(n_4446),
.Y(n_5912)
);

BUFx2_ASAP7_75t_L g5913 ( 
.A(n_4684),
.Y(n_5913)
);

CKINVDCx11_ASAP7_75t_R g5914 ( 
.A(n_5338),
.Y(n_5914)
);

INVx2_ASAP7_75t_SL g5915 ( 
.A(n_5528),
.Y(n_5915)
);

NAND2x2_ASAP7_75t_L g5916 ( 
.A(n_4686),
.B(n_4366),
.Y(n_5916)
);

AOI22xp5_ASAP7_75t_L g5917 ( 
.A1(n_4887),
.A2(n_4209),
.B1(n_4254),
.B2(n_4195),
.Y(n_5917)
);

NAND2xp5_ASAP7_75t_L g5918 ( 
.A(n_5292),
.B(n_4458),
.Y(n_5918)
);

BUFx2_ASAP7_75t_L g5919 ( 
.A(n_4731),
.Y(n_5919)
);

AO21x2_ASAP7_75t_L g5920 ( 
.A1(n_4996),
.A2(n_4675),
.B(n_4671),
.Y(n_5920)
);

INVx2_ASAP7_75t_SL g5921 ( 
.A(n_5528),
.Y(n_5921)
);

NAND2xp5_ASAP7_75t_L g5922 ( 
.A(n_5157),
.B(n_4458),
.Y(n_5922)
);

INVx1_ASAP7_75t_L g5923 ( 
.A(n_4683),
.Y(n_5923)
);

INVx5_ASAP7_75t_L g5924 ( 
.A(n_5528),
.Y(n_5924)
);

BUFx2_ASAP7_75t_L g5925 ( 
.A(n_4731),
.Y(n_5925)
);

INVx5_ASAP7_75t_L g5926 ( 
.A(n_5528),
.Y(n_5926)
);

AND2x4_ASAP7_75t_L g5927 ( 
.A(n_5528),
.B(n_4443),
.Y(n_5927)
);

INVx8_ASAP7_75t_L g5928 ( 
.A(n_4923),
.Y(n_5928)
);

INVx1_ASAP7_75t_L g5929 ( 
.A(n_4685),
.Y(n_5929)
);

AOI22xp5_ASAP7_75t_L g5930 ( 
.A1(n_5271),
.A2(n_4254),
.B1(n_4255),
.B2(n_4209),
.Y(n_5930)
);

OAI22xp5_ASAP7_75t_L g5931 ( 
.A1(n_5071),
.A2(n_4226),
.B1(n_4158),
.B2(n_4151),
.Y(n_5931)
);

INVx2_ASAP7_75t_SL g5932 ( 
.A(n_5093),
.Y(n_5932)
);

AND2x4_ASAP7_75t_L g5933 ( 
.A(n_5093),
.B(n_5106),
.Y(n_5933)
);

INVxp67_ASAP7_75t_L g5934 ( 
.A(n_4731),
.Y(n_5934)
);

INVx3_ASAP7_75t_L g5935 ( 
.A(n_4991),
.Y(n_5935)
);

BUFx12f_ASAP7_75t_L g5936 ( 
.A(n_5324),
.Y(n_5936)
);

INVx3_ASAP7_75t_L g5937 ( 
.A(n_5004),
.Y(n_5937)
);

NOR2xp33_ASAP7_75t_L g5938 ( 
.A(n_5108),
.B(n_4460),
.Y(n_5938)
);

HB1xp67_ASAP7_75t_L g5939 ( 
.A(n_4770),
.Y(n_5939)
);

NOR2xp33_ASAP7_75t_L g5940 ( 
.A(n_5108),
.B(n_4460),
.Y(n_5940)
);

OR2x2_ASAP7_75t_L g5941 ( 
.A(n_5478),
.B(n_4156),
.Y(n_5941)
);

BUFx12f_ASAP7_75t_L g5942 ( 
.A(n_5338),
.Y(n_5942)
);

INVx1_ASAP7_75t_L g5943 ( 
.A(n_4685),
.Y(n_5943)
);

INVx1_ASAP7_75t_L g5944 ( 
.A(n_4689),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_4689),
.Y(n_5945)
);

AND2x6_ASAP7_75t_L g5946 ( 
.A(n_4748),
.B(n_4209),
.Y(n_5946)
);

NAND2xp5_ASAP7_75t_L g5947 ( 
.A(n_5330),
.B(n_4462),
.Y(n_5947)
);

O2A1O1Ixp33_ASAP7_75t_L g5948 ( 
.A1(n_5083),
.A2(n_4463),
.B(n_4465),
.C(n_4462),
.Y(n_5948)
);

INVx3_ASAP7_75t_L g5949 ( 
.A(n_5004),
.Y(n_5949)
);

INVx5_ASAP7_75t_L g5950 ( 
.A(n_5283),
.Y(n_5950)
);

A2O1A1Ixp33_ASAP7_75t_L g5951 ( 
.A1(n_5083),
.A2(n_5364),
.B(n_5279),
.C(n_5281),
.Y(n_5951)
);

CKINVDCx5p33_ASAP7_75t_R g5952 ( 
.A(n_5340),
.Y(n_5952)
);

OAI221xp5_ASAP7_75t_L g5953 ( 
.A1(n_5281),
.A2(n_4575),
.B1(n_4514),
.B2(n_4467),
.C(n_4473),
.Y(n_5953)
);

INVxp67_ASAP7_75t_L g5954 ( 
.A(n_4806),
.Y(n_5954)
);

INVx2_ASAP7_75t_SL g5955 ( 
.A(n_5093),
.Y(n_5955)
);

INVx3_ASAP7_75t_L g5956 ( 
.A(n_5004),
.Y(n_5956)
);

INVx3_ASAP7_75t_SL g5957 ( 
.A(n_4781),
.Y(n_5957)
);

BUFx4f_ASAP7_75t_L g5958 ( 
.A(n_4862),
.Y(n_5958)
);

INVxp67_ASAP7_75t_SL g5959 ( 
.A(n_4806),
.Y(n_5959)
);

AND2x6_ASAP7_75t_L g5960 ( 
.A(n_4715),
.B(n_4254),
.Y(n_5960)
);

AOI22xp33_ASAP7_75t_L g5961 ( 
.A1(n_5248),
.A2(n_4450),
.B1(n_4472),
.B2(n_4449),
.Y(n_5961)
);

OAI22xp5_ASAP7_75t_L g5962 ( 
.A1(n_5101),
.A2(n_4425),
.B1(n_4309),
.B2(n_4123),
.Y(n_5962)
);

INVx1_ASAP7_75t_L g5963 ( 
.A(n_4695),
.Y(n_5963)
);

NOR2xp33_ASAP7_75t_SL g5964 ( 
.A(n_5101),
.B(n_4232),
.Y(n_5964)
);

INVx1_ASAP7_75t_SL g5965 ( 
.A(n_5018),
.Y(n_5965)
);

INVx1_ASAP7_75t_L g5966 ( 
.A(n_4695),
.Y(n_5966)
);

INVx1_ASAP7_75t_L g5967 ( 
.A(n_4707),
.Y(n_5967)
);

CKINVDCx5p33_ASAP7_75t_R g5968 ( 
.A(n_5340),
.Y(n_5968)
);

OAI21x1_ASAP7_75t_L g5969 ( 
.A1(n_5176),
.A2(n_4278),
.B(n_4166),
.Y(n_5969)
);

BUFx2_ASAP7_75t_L g5970 ( 
.A(n_4806),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_4707),
.Y(n_5971)
);

INVx1_ASAP7_75t_L g5972 ( 
.A(n_4719),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_4719),
.Y(n_5973)
);

NAND2xp5_ASAP7_75t_L g5974 ( 
.A(n_5330),
.B(n_4463),
.Y(n_5974)
);

O2A1O1Ixp33_ASAP7_75t_L g5975 ( 
.A1(n_4924),
.A2(n_5107),
.B(n_5162),
.C(n_5253),
.Y(n_5975)
);

AOI22xp33_ASAP7_75t_L g5976 ( 
.A1(n_5248),
.A2(n_4450),
.B1(n_4472),
.B2(n_4449),
.Y(n_5976)
);

NAND2xp5_ASAP7_75t_L g5977 ( 
.A(n_5315),
.B(n_4465),
.Y(n_5977)
);

HB1xp67_ASAP7_75t_L g5978 ( 
.A(n_4820),
.Y(n_5978)
);

NAND2xp5_ASAP7_75t_L g5979 ( 
.A(n_5315),
.B(n_4467),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_4728),
.Y(n_5980)
);

OR2x6_ASAP7_75t_L g5981 ( 
.A(n_5283),
.B(n_4152),
.Y(n_5981)
);

INVx4_ASAP7_75t_L g5982 ( 
.A(n_4787),
.Y(n_5982)
);

INVx3_ASAP7_75t_L g5983 ( 
.A(n_5004),
.Y(n_5983)
);

AOI21xp5_ASAP7_75t_L g5984 ( 
.A1(n_5291),
.A2(n_4475),
.B(n_4473),
.Y(n_5984)
);

INVx1_ASAP7_75t_L g5985 ( 
.A(n_4728),
.Y(n_5985)
);

AOI21xp5_ASAP7_75t_L g5986 ( 
.A1(n_5280),
.A2(n_4476),
.B(n_4475),
.Y(n_5986)
);

OR2x2_ASAP7_75t_L g5987 ( 
.A(n_4810),
.B(n_4156),
.Y(n_5987)
);

AOI22xp5_ASAP7_75t_L g5988 ( 
.A1(n_4919),
.A2(n_4262),
.B1(n_4289),
.B2(n_4255),
.Y(n_5988)
);

INVx3_ASAP7_75t_L g5989 ( 
.A(n_5004),
.Y(n_5989)
);

OAI22xp5_ASAP7_75t_L g5990 ( 
.A1(n_5162),
.A2(n_4309),
.B1(n_4425),
.B2(n_4455),
.Y(n_5990)
);

BUFx12f_ASAP7_75t_L g5991 ( 
.A(n_5340),
.Y(n_5991)
);

AOI22xp33_ASAP7_75t_L g5992 ( 
.A1(n_5048),
.A2(n_4472),
.B1(n_4450),
.B2(n_4262),
.Y(n_5992)
);

O2A1O1Ixp33_ASAP7_75t_L g5993 ( 
.A1(n_5107),
.A2(n_4480),
.B(n_4481),
.C(n_4476),
.Y(n_5993)
);

INVx3_ASAP7_75t_L g5994 ( 
.A(n_5004),
.Y(n_5994)
);

INVx8_ASAP7_75t_L g5995 ( 
.A(n_5283),
.Y(n_5995)
);

BUFx3_ASAP7_75t_L g5996 ( 
.A(n_5225),
.Y(n_5996)
);

BUFx3_ASAP7_75t_L g5997 ( 
.A(n_5225),
.Y(n_5997)
);

INVx5_ASAP7_75t_L g5998 ( 
.A(n_5283),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_4738),
.Y(n_5999)
);

INVx3_ASAP7_75t_L g6000 ( 
.A(n_5032),
.Y(n_6000)
);

BUFx2_ASAP7_75t_R g6001 ( 
.A(n_5428),
.Y(n_6001)
);

INVx2_ASAP7_75t_SL g6002 ( 
.A(n_5106),
.Y(n_6002)
);

INVx5_ASAP7_75t_L g6003 ( 
.A(n_5283),
.Y(n_6003)
);

AND2x4_ASAP7_75t_L g6004 ( 
.A(n_5106),
.B(n_5109),
.Y(n_6004)
);

OAI22xp5_ASAP7_75t_L g6005 ( 
.A1(n_5232),
.A2(n_5212),
.B1(n_4819),
.B2(n_4858),
.Y(n_6005)
);

AOI22xp33_ASAP7_75t_L g6006 ( 
.A1(n_5048),
.A2(n_5254),
.B1(n_5041),
.B2(n_4980),
.Y(n_6006)
);

OAI22xp5_ASAP7_75t_L g6007 ( 
.A1(n_5232),
.A2(n_4309),
.B1(n_4425),
.B2(n_3831),
.Y(n_6007)
);

OAI22xp5_ASAP7_75t_L g6008 ( 
.A1(n_5212),
.A2(n_4425),
.B1(n_3831),
.B2(n_4480),
.Y(n_6008)
);

HB1xp67_ASAP7_75t_L g6009 ( 
.A(n_4820),
.Y(n_6009)
);

BUFx2_ASAP7_75t_L g6010 ( 
.A(n_4810),
.Y(n_6010)
);

NAND2x2_ASAP7_75t_L g6011 ( 
.A(n_4686),
.B(n_3830),
.Y(n_6011)
);

AND2x2_ASAP7_75t_L g6012 ( 
.A(n_5407),
.B(n_4867),
.Y(n_6012)
);

AOI22xp5_ASAP7_75t_L g6013 ( 
.A1(n_4919),
.A2(n_4262),
.B1(n_4289),
.B2(n_4255),
.Y(n_6013)
);

AOI22xp5_ASAP7_75t_L g6014 ( 
.A1(n_5085),
.A2(n_5200),
.B1(n_4980),
.B2(n_5254),
.Y(n_6014)
);

AOI21xp5_ASAP7_75t_L g6015 ( 
.A1(n_5280),
.A2(n_4496),
.B(n_4481),
.Y(n_6015)
);

INVx3_ASAP7_75t_L g6016 ( 
.A(n_5032),
.Y(n_6016)
);

OAI22xp5_ASAP7_75t_L g6017 ( 
.A1(n_4816),
.A2(n_4425),
.B1(n_4508),
.B2(n_4496),
.Y(n_6017)
);

INVx6_ASAP7_75t_L g6018 ( 
.A(n_4853),
.Y(n_6018)
);

INVx3_ASAP7_75t_L g6019 ( 
.A(n_5032),
.Y(n_6019)
);

CKINVDCx20_ASAP7_75t_R g6020 ( 
.A(n_4925),
.Y(n_6020)
);

INVx3_ASAP7_75t_L g6021 ( 
.A(n_5032),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_4738),
.Y(n_6022)
);

NAND2xp5_ASAP7_75t_L g6023 ( 
.A(n_5339),
.B(n_5342),
.Y(n_6023)
);

NAND2xp33_ASAP7_75t_SL g6024 ( 
.A(n_4781),
.B(n_4634),
.Y(n_6024)
);

INVx6_ASAP7_75t_L g6025 ( 
.A(n_4853),
.Y(n_6025)
);

INVx2_ASAP7_75t_SL g6026 ( 
.A(n_5109),
.Y(n_6026)
);

INVx1_ASAP7_75t_SL g6027 ( 
.A(n_5018),
.Y(n_6027)
);

OAI21xp33_ASAP7_75t_L g6028 ( 
.A1(n_5187),
.A2(n_4509),
.B(n_4508),
.Y(n_6028)
);

BUFx6f_ASAP7_75t_L g6029 ( 
.A(n_5032),
.Y(n_6029)
);

OR2x2_ASAP7_75t_L g6030 ( 
.A(n_4810),
.B(n_4159),
.Y(n_6030)
);

OAI22xp5_ASAP7_75t_L g6031 ( 
.A1(n_4816),
.A2(n_4512),
.B1(n_4513),
.B2(n_4509),
.Y(n_6031)
);

NAND2xp5_ASAP7_75t_L g6032 ( 
.A(n_5339),
.B(n_5342),
.Y(n_6032)
);

BUFx12f_ASAP7_75t_L g6033 ( 
.A(n_5356),
.Y(n_6033)
);

OR2x2_ASAP7_75t_L g6034 ( 
.A(n_4828),
.B(n_4159),
.Y(n_6034)
);

INVx2_ASAP7_75t_SL g6035 ( 
.A(n_5109),
.Y(n_6035)
);

INVx4_ASAP7_75t_L g6036 ( 
.A(n_4787),
.Y(n_6036)
);

BUFx3_ASAP7_75t_L g6037 ( 
.A(n_5225),
.Y(n_6037)
);

OAI22xp5_ASAP7_75t_L g6038 ( 
.A1(n_4819),
.A2(n_4512),
.B1(n_4516),
.B2(n_4513),
.Y(n_6038)
);

OAI22xp5_ASAP7_75t_L g6039 ( 
.A1(n_4858),
.A2(n_4516),
.B1(n_4522),
.B2(n_4138),
.Y(n_6039)
);

INVx3_ASAP7_75t_L g6040 ( 
.A(n_5032),
.Y(n_6040)
);

INVx3_ASAP7_75t_L g6041 ( 
.A(n_5032),
.Y(n_6041)
);

NAND3xp33_ASAP7_75t_L g6042 ( 
.A(n_5160),
.B(n_4522),
.C(n_4618),
.Y(n_6042)
);

INVx2_ASAP7_75t_SL g6043 ( 
.A(n_5118),
.Y(n_6043)
);

NAND2xp5_ASAP7_75t_L g6044 ( 
.A(n_5187),
.B(n_4039),
.Y(n_6044)
);

INVxp67_ASAP7_75t_L g6045 ( 
.A(n_4828),
.Y(n_6045)
);

NAND2xp5_ASAP7_75t_L g6046 ( 
.A(n_5320),
.B(n_4039),
.Y(n_6046)
);

NAND2xp5_ASAP7_75t_L g6047 ( 
.A(n_5320),
.B(n_4047),
.Y(n_6047)
);

NAND2xp5_ASAP7_75t_L g6048 ( 
.A(n_4883),
.B(n_4047),
.Y(n_6048)
);

AOI22xp5_ASAP7_75t_L g6049 ( 
.A1(n_5085),
.A2(n_4262),
.B1(n_4289),
.B2(n_4255),
.Y(n_6049)
);

CKINVDCx5p33_ASAP7_75t_R g6050 ( 
.A(n_5356),
.Y(n_6050)
);

NOR2x1_ASAP7_75t_SL g6051 ( 
.A(n_4899),
.B(n_4152),
.Y(n_6051)
);

INVx2_ASAP7_75t_SL g6052 ( 
.A(n_5118),
.Y(n_6052)
);

O2A1O1Ixp5_ASAP7_75t_L g6053 ( 
.A1(n_5138),
.A2(n_4026),
.B(n_4033),
.C(n_3972),
.Y(n_6053)
);

INVxp67_ASAP7_75t_L g6054 ( 
.A(n_4828),
.Y(n_6054)
);

A2O1A1Ixp33_ASAP7_75t_L g6055 ( 
.A1(n_5364),
.A2(n_3964),
.B(n_4069),
.C(n_3865),
.Y(n_6055)
);

AO21x2_ASAP7_75t_L g6056 ( 
.A1(n_4996),
.A2(n_4675),
.B(n_4671),
.Y(n_6056)
);

NAND2xp5_ASAP7_75t_L g6057 ( 
.A(n_4883),
.B(n_4049),
.Y(n_6057)
);

INVx2_ASAP7_75t_SL g6058 ( 
.A(n_5118),
.Y(n_6058)
);

AOI22xp33_ASAP7_75t_L g6059 ( 
.A1(n_5041),
.A2(n_4292),
.B1(n_4331),
.B2(n_4289),
.Y(n_6059)
);

NAND2xp5_ASAP7_75t_L g6060 ( 
.A(n_5075),
.B(n_4049),
.Y(n_6060)
);

INVx1_ASAP7_75t_L g6061 ( 
.A(n_4743),
.Y(n_6061)
);

HB1xp67_ASAP7_75t_L g6062 ( 
.A(n_4990),
.Y(n_6062)
);

INVx4_ASAP7_75t_L g6063 ( 
.A(n_4899),
.Y(n_6063)
);

NAND2xp5_ASAP7_75t_L g6064 ( 
.A(n_5075),
.B(n_5455),
.Y(n_6064)
);

NAND2xp5_ASAP7_75t_L g6065 ( 
.A(n_5455),
.B(n_4060),
.Y(n_6065)
);

INVx3_ASAP7_75t_L g6066 ( 
.A(n_5045),
.Y(n_6066)
);

AOI21xp5_ASAP7_75t_L g6067 ( 
.A1(n_5235),
.A2(n_4468),
.B(n_4461),
.Y(n_6067)
);

INVx1_ASAP7_75t_L g6068 ( 
.A(n_4743),
.Y(n_6068)
);

CKINVDCx5p33_ASAP7_75t_R g6069 ( 
.A(n_5356),
.Y(n_6069)
);

AOI22xp5_ASAP7_75t_L g6070 ( 
.A1(n_5200),
.A2(n_4331),
.B1(n_4340),
.B2(n_4292),
.Y(n_6070)
);

AOI21xp5_ASAP7_75t_L g6071 ( 
.A1(n_5235),
.A2(n_4468),
.B(n_4461),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_4749),
.Y(n_6072)
);

O2A1O1Ixp33_ASAP7_75t_L g6073 ( 
.A1(n_5253),
.A2(n_4392),
.B(n_4399),
.C(n_4266),
.Y(n_6073)
);

NAND2xp5_ASAP7_75t_SL g6074 ( 
.A(n_4781),
.B(n_4243),
.Y(n_6074)
);

NAND2xp5_ASAP7_75t_L g6075 ( 
.A(n_5460),
.B(n_4060),
.Y(n_6075)
);

AND2x2_ASAP7_75t_L g6076 ( 
.A(n_4867),
.B(n_4670),
.Y(n_6076)
);

BUFx12f_ASAP7_75t_L g6077 ( 
.A(n_5021),
.Y(n_6077)
);

NAND2xp5_ASAP7_75t_L g6078 ( 
.A(n_5460),
.B(n_4233),
.Y(n_6078)
);

AOI22xp5_ASAP7_75t_L g6079 ( 
.A1(n_4680),
.A2(n_4331),
.B1(n_4340),
.B2(n_4292),
.Y(n_6079)
);

OAI21x1_ASAP7_75t_L g6080 ( 
.A1(n_5176),
.A2(n_4278),
.B(n_4166),
.Y(n_6080)
);

AOI21xp5_ASAP7_75t_SL g6081 ( 
.A1(n_5279),
.A2(n_3879),
.B(n_3836),
.Y(n_6081)
);

AOI21xp5_ASAP7_75t_L g6082 ( 
.A1(n_4986),
.A2(n_4468),
.B(n_4461),
.Y(n_6082)
);

AOI22xp5_ASAP7_75t_L g6083 ( 
.A1(n_4680),
.A2(n_4331),
.B1(n_4340),
.B2(n_4292),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_4749),
.Y(n_6084)
);

INVx4_ASAP7_75t_L g6085 ( 
.A(n_4899),
.Y(n_6085)
);

HB1xp67_ASAP7_75t_L g6086 ( 
.A(n_4990),
.Y(n_6086)
);

INVx8_ASAP7_75t_L g6087 ( 
.A(n_5283),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_4764),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_4764),
.Y(n_6089)
);

AOI21xp5_ASAP7_75t_L g6090 ( 
.A1(n_4986),
.A2(n_4585),
.B(n_4489),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_4771),
.Y(n_6091)
);

NAND2xp5_ASAP7_75t_L g6092 ( 
.A(n_5494),
.B(n_4233),
.Y(n_6092)
);

AND2x2_ASAP7_75t_L g6093 ( 
.A(n_4867),
.B(n_4670),
.Y(n_6093)
);

AND2x2_ASAP7_75t_L g6094 ( 
.A(n_5068),
.B(n_4589),
.Y(n_6094)
);

INVx4_ASAP7_75t_L g6095 ( 
.A(n_4899),
.Y(n_6095)
);

NAND2xp5_ASAP7_75t_L g6096 ( 
.A(n_5494),
.B(n_4233),
.Y(n_6096)
);

AOI21x1_ASAP7_75t_L g6097 ( 
.A1(n_5117),
.A2(n_4589),
.B(n_4237),
.Y(n_6097)
);

CKINVDCx5p33_ASAP7_75t_R g6098 ( 
.A(n_4754),
.Y(n_6098)
);

AOI22xp5_ASAP7_75t_L g6099 ( 
.A1(n_5296),
.A2(n_4774),
.B1(n_5249),
.B2(n_5057),
.Y(n_6099)
);

AOI21xp5_ASAP7_75t_L g6100 ( 
.A1(n_5001),
.A2(n_4585),
.B(n_4489),
.Y(n_6100)
);

NAND2x1p5_ASAP7_75t_L g6101 ( 
.A(n_4921),
.B(n_3964),
.Y(n_6101)
);

INVx3_ASAP7_75t_L g6102 ( 
.A(n_5045),
.Y(n_6102)
);

AND2x2_ASAP7_75t_L g6103 ( 
.A(n_5068),
.B(n_4335),
.Y(n_6103)
);

AND2x4_ASAP7_75t_L g6104 ( 
.A(n_5425),
.B(n_5436),
.Y(n_6104)
);

HB1xp67_ASAP7_75t_L g6105 ( 
.A(n_4914),
.Y(n_6105)
);

INVx1_ASAP7_75t_L g6106 ( 
.A(n_4771),
.Y(n_6106)
);

AOI21xp5_ASAP7_75t_L g6107 ( 
.A1(n_5001),
.A2(n_4585),
.B(n_4489),
.Y(n_6107)
);

NAND2xp5_ASAP7_75t_L g6108 ( 
.A(n_5496),
.B(n_4252),
.Y(n_6108)
);

INVx1_ASAP7_75t_SL g6109 ( 
.A(n_5074),
.Y(n_6109)
);

INVx1_ASAP7_75t_SL g6110 ( 
.A(n_5074),
.Y(n_6110)
);

AOI21xp5_ASAP7_75t_L g6111 ( 
.A1(n_5013),
.A2(n_4600),
.B(n_4599),
.Y(n_6111)
);

BUFx2_ASAP7_75t_L g6112 ( 
.A(n_4857),
.Y(n_6112)
);

INVx4_ASAP7_75t_L g6113 ( 
.A(n_4899),
.Y(n_6113)
);

INVx1_ASAP7_75t_SL g6114 ( 
.A(n_5211),
.Y(n_6114)
);

NAND2xp5_ASAP7_75t_L g6115 ( 
.A(n_5496),
.B(n_4252),
.Y(n_6115)
);

OAI22xp5_ASAP7_75t_L g6116 ( 
.A1(n_4700),
.A2(n_4741),
.B1(n_5160),
.B2(n_4735),
.Y(n_6116)
);

AOI221x1_ASAP7_75t_L g6117 ( 
.A1(n_4733),
.A2(n_4735),
.B1(n_4992),
.B2(n_5286),
.C(n_4965),
.Y(n_6117)
);

AND2x2_ASAP7_75t_L g6118 ( 
.A(n_5068),
.B(n_4335),
.Y(n_6118)
);

AOI21xp5_ASAP7_75t_L g6119 ( 
.A1(n_5013),
.A2(n_4600),
.B(n_4599),
.Y(n_6119)
);

AOI21xp5_ASAP7_75t_L g6120 ( 
.A1(n_5014),
.A2(n_4600),
.B(n_4599),
.Y(n_6120)
);

AND2x2_ASAP7_75t_SL g6121 ( 
.A(n_5178),
.B(n_4335),
.Y(n_6121)
);

INVx2_ASAP7_75t_SL g6122 ( 
.A(n_5425),
.Y(n_6122)
);

NAND2xp5_ASAP7_75t_L g6123 ( 
.A(n_4811),
.B(n_4911),
.Y(n_6123)
);

NAND2x1p5_ASAP7_75t_L g6124 ( 
.A(n_5178),
.B(n_3964),
.Y(n_6124)
);

INVx1_ASAP7_75t_L g6125 ( 
.A(n_4779),
.Y(n_6125)
);

BUFx3_ASAP7_75t_L g6126 ( 
.A(n_5225),
.Y(n_6126)
);

INVx1_ASAP7_75t_L g6127 ( 
.A(n_4779),
.Y(n_6127)
);

OR2x2_ASAP7_75t_SL g6128 ( 
.A(n_4733),
.B(n_4068),
.Y(n_6128)
);

O2A1O1Ixp33_ASAP7_75t_L g6129 ( 
.A1(n_5138),
.A2(n_4266),
.B(n_4399),
.C(n_4392),
.Y(n_6129)
);

INVx2_ASAP7_75t_SL g6130 ( 
.A(n_5425),
.Y(n_6130)
);

BUFx2_ASAP7_75t_L g6131 ( 
.A(n_4857),
.Y(n_6131)
);

AND2x2_ASAP7_75t_L g6132 ( 
.A(n_5100),
.B(n_4335),
.Y(n_6132)
);

INVx1_ASAP7_75t_SL g6133 ( 
.A(n_5211),
.Y(n_6133)
);

INVx1_ASAP7_75t_L g6134 ( 
.A(n_4783),
.Y(n_6134)
);

NAND2xp5_ASAP7_75t_L g6135 ( 
.A(n_4811),
.B(n_4252),
.Y(n_6135)
);

AND2x2_ASAP7_75t_L g6136 ( 
.A(n_5100),
.B(n_4335),
.Y(n_6136)
);

BUFx3_ASAP7_75t_L g6137 ( 
.A(n_5225),
.Y(n_6137)
);

BUFx3_ASAP7_75t_L g6138 ( 
.A(n_5225),
.Y(n_6138)
);

INVx1_ASAP7_75t_L g6139 ( 
.A(n_4783),
.Y(n_6139)
);

INVx2_ASAP7_75t_SL g6140 ( 
.A(n_5425),
.Y(n_6140)
);

AND2x2_ASAP7_75t_L g6141 ( 
.A(n_5100),
.B(n_4335),
.Y(n_6141)
);

BUFx3_ASAP7_75t_L g6142 ( 
.A(n_5225),
.Y(n_6142)
);

AND3x1_ASAP7_75t_SL g6143 ( 
.A(n_4900),
.B(n_4176),
.C(n_4171),
.Y(n_6143)
);

INVx1_ASAP7_75t_L g6144 ( 
.A(n_4785),
.Y(n_6144)
);

AOI22xp33_ASAP7_75t_L g6145 ( 
.A1(n_5249),
.A2(n_4386),
.B1(n_4405),
.B2(n_4340),
.Y(n_6145)
);

HB1xp67_ASAP7_75t_L g6146 ( 
.A(n_4914),
.Y(n_6146)
);

AND2x2_ASAP7_75t_L g6147 ( 
.A(n_5127),
.B(n_4423),
.Y(n_6147)
);

NOR2xp33_ASAP7_75t_L g6148 ( 
.A(n_4755),
.B(n_4266),
.Y(n_6148)
);

NAND2xp5_ASAP7_75t_L g6149 ( 
.A(n_4911),
.B(n_4444),
.Y(n_6149)
);

AND2x2_ASAP7_75t_L g6150 ( 
.A(n_5127),
.B(n_4423),
.Y(n_6150)
);

BUFx2_ASAP7_75t_L g6151 ( 
.A(n_4857),
.Y(n_6151)
);

CKINVDCx5p33_ASAP7_75t_R g6152 ( 
.A(n_4754),
.Y(n_6152)
);

NOR2xp33_ASAP7_75t_L g6153 ( 
.A(n_4755),
.B(n_4392),
.Y(n_6153)
);

INVx1_ASAP7_75t_L g6154 ( 
.A(n_4785),
.Y(n_6154)
);

NOR2xp33_ASAP7_75t_SL g6155 ( 
.A(n_5367),
.B(n_5396),
.Y(n_6155)
);

INVx2_ASAP7_75t_SL g6156 ( 
.A(n_5436),
.Y(n_6156)
);

INVx1_ASAP7_75t_L g6157 ( 
.A(n_4790),
.Y(n_6157)
);

NAND2xp5_ASAP7_75t_SL g6158 ( 
.A(n_4781),
.B(n_4399),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_4790),
.Y(n_6159)
);

INVx1_ASAP7_75t_SL g6160 ( 
.A(n_5246),
.Y(n_6160)
);

NOR2xp33_ASAP7_75t_SL g6161 ( 
.A(n_5367),
.B(n_4232),
.Y(n_6161)
);

NOR2xp33_ASAP7_75t_L g6162 ( 
.A(n_4803),
.B(n_4418),
.Y(n_6162)
);

OAI22xp5_ASAP7_75t_L g6163 ( 
.A1(n_4700),
.A2(n_4092),
.B1(n_4103),
.B2(n_4089),
.Y(n_6163)
);

INVxp67_ASAP7_75t_L g6164 ( 
.A(n_4880),
.Y(n_6164)
);

BUFx2_ASAP7_75t_SL g6165 ( 
.A(n_5541),
.Y(n_6165)
);

OAI22xp5_ASAP7_75t_L g6166 ( 
.A1(n_4741),
.A2(n_4092),
.B1(n_4103),
.B2(n_4089),
.Y(n_6166)
);

BUFx3_ASAP7_75t_L g6167 ( 
.A(n_5225),
.Y(n_6167)
);

INVx3_ASAP7_75t_L g6168 ( 
.A(n_5060),
.Y(n_6168)
);

CKINVDCx5p33_ASAP7_75t_R g6169 ( 
.A(n_4754),
.Y(n_6169)
);

AOI21x1_ASAP7_75t_L g6170 ( 
.A1(n_5267),
.A2(n_4237),
.B(n_4221),
.Y(n_6170)
);

CKINVDCx5p33_ASAP7_75t_R g6171 ( 
.A(n_4818),
.Y(n_6171)
);

AND2x2_ASAP7_75t_L g6172 ( 
.A(n_5127),
.B(n_4423),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_4793),
.Y(n_6173)
);

AOI22xp5_ASAP7_75t_SL g6174 ( 
.A1(n_5249),
.A2(n_5344),
.B1(n_4928),
.B2(n_5006),
.Y(n_6174)
);

NAND2xp5_ASAP7_75t_L g6175 ( 
.A(n_5371),
.B(n_4444),
.Y(n_6175)
);

AOI22xp33_ASAP7_75t_L g6176 ( 
.A1(n_5249),
.A2(n_4405),
.B1(n_4424),
.B2(n_4386),
.Y(n_6176)
);

BUFx2_ASAP7_75t_L g6177 ( 
.A(n_4880),
.Y(n_6177)
);

A2O1A1Ixp33_ASAP7_75t_L g6178 ( 
.A1(n_5472),
.A2(n_4069),
.B(n_3964),
.C(n_3836),
.Y(n_6178)
);

BUFx4_ASAP7_75t_SL g6179 ( 
.A(n_5179),
.Y(n_6179)
);

NAND2xp5_ASAP7_75t_L g6180 ( 
.A(n_5371),
.B(n_4444),
.Y(n_6180)
);

BUFx10_ASAP7_75t_L g6181 ( 
.A(n_4708),
.Y(n_6181)
);

CKINVDCx5p33_ASAP7_75t_R g6182 ( 
.A(n_4818),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_4793),
.Y(n_6183)
);

INVx1_ASAP7_75t_L g6184 ( 
.A(n_4796),
.Y(n_6184)
);

CKINVDCx5p33_ASAP7_75t_R g6185 ( 
.A(n_4818),
.Y(n_6185)
);

A2O1A1Ixp33_ASAP7_75t_L g6186 ( 
.A1(n_5472),
.A2(n_4069),
.B(n_3964),
.C(n_3836),
.Y(n_6186)
);

INVx1_ASAP7_75t_L g6187 ( 
.A(n_4796),
.Y(n_6187)
);

BUFx8_ASAP7_75t_SL g6188 ( 
.A(n_4927),
.Y(n_6188)
);

INVx1_ASAP7_75t_L g6189 ( 
.A(n_4804),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_4804),
.Y(n_6190)
);

INVx2_ASAP7_75t_SL g6191 ( 
.A(n_5446),
.Y(n_6191)
);

OR2x6_ASAP7_75t_L g6192 ( 
.A(n_5390),
.B(n_4152),
.Y(n_6192)
);

BUFx3_ASAP7_75t_L g6193 ( 
.A(n_5225),
.Y(n_6193)
);

BUFx2_ASAP7_75t_L g6194 ( 
.A(n_4880),
.Y(n_6194)
);

OR2x6_ASAP7_75t_SL g6195 ( 
.A(n_5378),
.B(n_4171),
.Y(n_6195)
);

INVx1_ASAP7_75t_L g6196 ( 
.A(n_4805),
.Y(n_6196)
);

OAI22xp33_ASAP7_75t_L g6197 ( 
.A1(n_5296),
.A2(n_4069),
.B1(n_4394),
.B2(n_4304),
.Y(n_6197)
);

BUFx12f_ASAP7_75t_L g6198 ( 
.A(n_5021),
.Y(n_6198)
);

INVx2_ASAP7_75t_SL g6199 ( 
.A(n_5446),
.Y(n_6199)
);

NAND2xp5_ASAP7_75t_L g6200 ( 
.A(n_5090),
.B(n_4552),
.Y(n_6200)
);

INVx1_ASAP7_75t_L g6201 ( 
.A(n_4805),
.Y(n_6201)
);

INVxp67_ASAP7_75t_SL g6202 ( 
.A(n_4902),
.Y(n_6202)
);

INVx1_ASAP7_75t_L g6203 ( 
.A(n_4836),
.Y(n_6203)
);

INVx3_ASAP7_75t_L g6204 ( 
.A(n_5060),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_4836),
.Y(n_6205)
);

HB1xp67_ASAP7_75t_L g6206 ( 
.A(n_4930),
.Y(n_6206)
);

NAND2xp5_ASAP7_75t_L g6207 ( 
.A(n_5090),
.B(n_4552),
.Y(n_6207)
);

INVx1_ASAP7_75t_L g6208 ( 
.A(n_4847),
.Y(n_6208)
);

OR2x2_ASAP7_75t_L g6209 ( 
.A(n_4902),
.B(n_4176),
.Y(n_6209)
);

OAI22xp5_ASAP7_75t_L g6210 ( 
.A1(n_5221),
.A2(n_4843),
.B1(n_5286),
.B2(n_4803),
.Y(n_6210)
);

AO32x2_ASAP7_75t_L g6211 ( 
.A1(n_5319),
.A2(n_5303),
.A3(n_5306),
.B1(n_5277),
.B2(n_5261),
.Y(n_6211)
);

BUFx4f_ASAP7_75t_L g6212 ( 
.A(n_4862),
.Y(n_6212)
);

OAI221xp5_ASAP7_75t_L g6213 ( 
.A1(n_5221),
.A2(n_4514),
.B1(n_4394),
.B2(n_4304),
.C(n_4613),
.Y(n_6213)
);

NOR2xp33_ASAP7_75t_L g6214 ( 
.A(n_5126),
.B(n_4418),
.Y(n_6214)
);

INVx3_ASAP7_75t_L g6215 ( 
.A(n_5122),
.Y(n_6215)
);

NAND2xp5_ASAP7_75t_SL g6216 ( 
.A(n_5516),
.B(n_4418),
.Y(n_6216)
);

NAND2xp5_ASAP7_75t_L g6217 ( 
.A(n_5126),
.B(n_4556),
.Y(n_6217)
);

BUFx2_ASAP7_75t_L g6218 ( 
.A(n_4902),
.Y(n_6218)
);

NAND2x1p5_ASAP7_75t_L g6219 ( 
.A(n_5293),
.B(n_5333),
.Y(n_6219)
);

OR2x2_ASAP7_75t_L g6220 ( 
.A(n_4954),
.B(n_4180),
.Y(n_6220)
);

NAND2xp5_ASAP7_75t_SL g6221 ( 
.A(n_5516),
.B(n_4086),
.Y(n_6221)
);

NAND2xp5_ASAP7_75t_SL g6222 ( 
.A(n_5182),
.B(n_5158),
.Y(n_6222)
);

INVx3_ASAP7_75t_L g6223 ( 
.A(n_5122),
.Y(n_6223)
);

NAND2xp5_ASAP7_75t_L g6224 ( 
.A(n_5152),
.B(n_4556),
.Y(n_6224)
);

BUFx3_ASAP7_75t_L g6225 ( 
.A(n_5318),
.Y(n_6225)
);

NAND2xp5_ASAP7_75t_L g6226 ( 
.A(n_5152),
.B(n_4574),
.Y(n_6226)
);

OR2x2_ASAP7_75t_L g6227 ( 
.A(n_4954),
.B(n_4180),
.Y(n_6227)
);

INVx6_ASAP7_75t_L g6228 ( 
.A(n_4853),
.Y(n_6228)
);

AOI22xp33_ASAP7_75t_L g6229 ( 
.A1(n_5057),
.A2(n_4386),
.B1(n_4424),
.B2(n_4405),
.Y(n_6229)
);

AOI22xp5_ASAP7_75t_L g6230 ( 
.A1(n_4774),
.A2(n_4405),
.B1(n_4424),
.B2(n_4386),
.Y(n_6230)
);

AOI222xp33_ASAP7_75t_L g6231 ( 
.A1(n_5395),
.A2(n_5240),
.B1(n_4843),
.B2(n_5505),
.C1(n_4869),
.C2(n_4821),
.Y(n_6231)
);

AOI21xp5_ASAP7_75t_L g6232 ( 
.A1(n_5014),
.A2(n_4655),
.B(n_4604),
.Y(n_6232)
);

NAND2xp5_ASAP7_75t_SL g6233 ( 
.A(n_5182),
.B(n_4086),
.Y(n_6233)
);

AOI22xp33_ASAP7_75t_L g6234 ( 
.A1(n_5395),
.A2(n_4424),
.B1(n_4532),
.B2(n_4441),
.Y(n_6234)
);

BUFx3_ASAP7_75t_L g6235 ( 
.A(n_5318),
.Y(n_6235)
);

NAND2x1p5_ASAP7_75t_L g6236 ( 
.A(n_5293),
.B(n_4069),
.Y(n_6236)
);

AOI22xp33_ASAP7_75t_L g6237 ( 
.A1(n_5240),
.A2(n_4441),
.B1(n_4553),
.B2(n_4532),
.Y(n_6237)
);

AND2x4_ASAP7_75t_L g6238 ( 
.A(n_5461),
.B(n_5473),
.Y(n_6238)
);

NAND2xp33_ASAP7_75t_L g6239 ( 
.A(n_4959),
.B(n_4634),
.Y(n_6239)
);

NAND2xp5_ASAP7_75t_L g6240 ( 
.A(n_5154),
.B(n_4574),
.Y(n_6240)
);

AOI22xp5_ASAP7_75t_L g6241 ( 
.A1(n_4772),
.A2(n_4532),
.B1(n_4553),
.B2(n_4441),
.Y(n_6241)
);

OR2x6_ASAP7_75t_L g6242 ( 
.A(n_5081),
.B(n_4514),
.Y(n_6242)
);

NAND2xp5_ASAP7_75t_SL g6243 ( 
.A(n_5158),
.B(n_4086),
.Y(n_6243)
);

OR2x6_ASAP7_75t_L g6244 ( 
.A(n_5081),
.B(n_5266),
.Y(n_6244)
);

INVx1_ASAP7_75t_SL g6245 ( 
.A(n_5246),
.Y(n_6245)
);

INVx5_ASAP7_75t_L g6246 ( 
.A(n_5318),
.Y(n_6246)
);

OAI22xp33_ASAP7_75t_L g6247 ( 
.A1(n_4778),
.A2(n_4069),
.B1(n_4394),
.B2(n_4304),
.Y(n_6247)
);

INVx1_ASAP7_75t_L g6248 ( 
.A(n_4847),
.Y(n_6248)
);

INVx1_ASAP7_75t_L g6249 ( 
.A(n_4854),
.Y(n_6249)
);

INVx1_ASAP7_75t_L g6250 ( 
.A(n_4854),
.Y(n_6250)
);

AOI22xp5_ASAP7_75t_L g6251 ( 
.A1(n_4772),
.A2(n_4532),
.B1(n_4553),
.B2(n_4441),
.Y(n_6251)
);

INVx3_ASAP7_75t_L g6252 ( 
.A(n_5122),
.Y(n_6252)
);

NAND2xp5_ASAP7_75t_L g6253 ( 
.A(n_5154),
.B(n_4574),
.Y(n_6253)
);

A2O1A1Ixp33_ASAP7_75t_L g6254 ( 
.A1(n_5505),
.A2(n_4069),
.B(n_3836),
.C(n_3976),
.Y(n_6254)
);

BUFx2_ASAP7_75t_L g6255 ( 
.A(n_4954),
.Y(n_6255)
);

INVx2_ASAP7_75t_SL g6256 ( 
.A(n_5461),
.Y(n_6256)
);

INVx5_ASAP7_75t_L g6257 ( 
.A(n_5318),
.Y(n_6257)
);

NAND2xp5_ASAP7_75t_L g6258 ( 
.A(n_5155),
.B(n_5161),
.Y(n_6258)
);

AND2x2_ASAP7_75t_L g6259 ( 
.A(n_5450),
.B(n_4428),
.Y(n_6259)
);

BUFx2_ASAP7_75t_L g6260 ( 
.A(n_4966),
.Y(n_6260)
);

AND2x2_ASAP7_75t_L g6261 ( 
.A(n_5450),
.B(n_4428),
.Y(n_6261)
);

INVx1_ASAP7_75t_L g6262 ( 
.A(n_4860),
.Y(n_6262)
);

BUFx4f_ASAP7_75t_L g6263 ( 
.A(n_5043),
.Y(n_6263)
);

NAND2x1p5_ASAP7_75t_L g6264 ( 
.A(n_5333),
.B(n_4069),
.Y(n_6264)
);

NAND2xp5_ASAP7_75t_L g6265 ( 
.A(n_5155),
.B(n_4592),
.Y(n_6265)
);

NOR2xp33_ASAP7_75t_R g6266 ( 
.A(n_4900),
.B(n_4326),
.Y(n_6266)
);

AOI22xp33_ASAP7_75t_L g6267 ( 
.A1(n_4979),
.A2(n_4553),
.B1(n_4558),
.B2(n_4069),
.Y(n_6267)
);

AND2x4_ASAP7_75t_L g6268 ( 
.A(n_5461),
.B(n_5473),
.Y(n_6268)
);

NAND2xp5_ASAP7_75t_L g6269 ( 
.A(n_5161),
.B(n_4592),
.Y(n_6269)
);

BUFx3_ASAP7_75t_L g6270 ( 
.A(n_5318),
.Y(n_6270)
);

INVx1_ASAP7_75t_L g6271 ( 
.A(n_4860),
.Y(n_6271)
);

INVx1_ASAP7_75t_L g6272 ( 
.A(n_4890),
.Y(n_6272)
);

A2O1A1Ixp33_ASAP7_75t_L g6273 ( 
.A1(n_5099),
.A2(n_3976),
.B(n_3988),
.C(n_3879),
.Y(n_6273)
);

BUFx12f_ASAP7_75t_L g6274 ( 
.A(n_5021),
.Y(n_6274)
);

BUFx12f_ASAP7_75t_L g6275 ( 
.A(n_5131),
.Y(n_6275)
);

BUFx3_ASAP7_75t_L g6276 ( 
.A(n_5318),
.Y(n_6276)
);

AND2x6_ASAP7_75t_L g6277 ( 
.A(n_4715),
.B(n_4558),
.Y(n_6277)
);

A2O1A1Ixp33_ASAP7_75t_L g6278 ( 
.A1(n_5099),
.A2(n_3976),
.B(n_3988),
.C(n_3879),
.Y(n_6278)
);

INVx1_ASAP7_75t_SL g6279 ( 
.A(n_5350),
.Y(n_6279)
);

BUFx12f_ASAP7_75t_L g6280 ( 
.A(n_5131),
.Y(n_6280)
);

NAND2xp33_ASAP7_75t_L g6281 ( 
.A(n_4959),
.B(n_4166),
.Y(n_6281)
);

INVx2_ASAP7_75t_SL g6282 ( 
.A(n_5473),
.Y(n_6282)
);

NOR2xp33_ASAP7_75t_L g6283 ( 
.A(n_5172),
.B(n_5181),
.Y(n_6283)
);

BUFx12f_ASAP7_75t_L g6284 ( 
.A(n_5131),
.Y(n_6284)
);

CKINVDCx8_ASAP7_75t_R g6285 ( 
.A(n_5318),
.Y(n_6285)
);

NOR2xp33_ASAP7_75t_SL g6286 ( 
.A(n_5396),
.B(n_4326),
.Y(n_6286)
);

AOI21xp5_ASAP7_75t_L g6287 ( 
.A1(n_5020),
.A2(n_4655),
.B(n_4604),
.Y(n_6287)
);

CKINVDCx5p33_ASAP7_75t_R g6288 ( 
.A(n_4927),
.Y(n_6288)
);

BUFx2_ASAP7_75t_L g6289 ( 
.A(n_4966),
.Y(n_6289)
);

NAND2xp5_ASAP7_75t_L g6290 ( 
.A(n_5172),
.B(n_4592),
.Y(n_6290)
);

CKINVDCx20_ASAP7_75t_R g6291 ( 
.A(n_4925),
.Y(n_6291)
);

OAI21xp5_ASAP7_75t_L g6292 ( 
.A1(n_4729),
.A2(n_4613),
.B(n_4514),
.Y(n_6292)
);

BUFx12f_ASAP7_75t_L g6293 ( 
.A(n_4927),
.Y(n_6293)
);

INVx1_ASAP7_75t_L g6294 ( 
.A(n_4890),
.Y(n_6294)
);

AND2x6_ASAP7_75t_L g6295 ( 
.A(n_4727),
.B(n_4558),
.Y(n_6295)
);

NOR2xp33_ASAP7_75t_L g6296 ( 
.A(n_5181),
.B(n_5208),
.Y(n_6296)
);

BUFx3_ASAP7_75t_L g6297 ( 
.A(n_5318),
.Y(n_6297)
);

AOI21xp5_ASAP7_75t_L g6298 ( 
.A1(n_5020),
.A2(n_5046),
.B(n_5029),
.Y(n_6298)
);

AOI21xp5_ASAP7_75t_L g6299 ( 
.A1(n_5029),
.A2(n_4655),
.B(n_4604),
.Y(n_6299)
);

AOI21x1_ASAP7_75t_L g6300 ( 
.A1(n_5267),
.A2(n_4237),
.B(n_4221),
.Y(n_6300)
);

BUFx3_ASAP7_75t_L g6301 ( 
.A(n_5318),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_4896),
.Y(n_6302)
);

INVx2_ASAP7_75t_SL g6303 ( 
.A(n_5479),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_4896),
.Y(n_6304)
);

AOI21xp5_ASAP7_75t_L g6305 ( 
.A1(n_5046),
.A2(n_4026),
.B(n_3972),
.Y(n_6305)
);

NAND2xp5_ASAP7_75t_L g6306 ( 
.A(n_5208),
.B(n_4595),
.Y(n_6306)
);

BUFx3_ASAP7_75t_L g6307 ( 
.A(n_5318),
.Y(n_6307)
);

OR2x2_ASAP7_75t_L g6308 ( 
.A(n_4966),
.B(n_4183),
.Y(n_6308)
);

INVx1_ASAP7_75t_L g6309 ( 
.A(n_4898),
.Y(n_6309)
);

OAI22xp5_ASAP7_75t_L g6310 ( 
.A1(n_4778),
.A2(n_4092),
.B1(n_4103),
.B2(n_4089),
.Y(n_6310)
);

OR2x2_ASAP7_75t_L g6311 ( 
.A(n_5026),
.B(n_4192),
.Y(n_6311)
);

OAI22xp5_ASAP7_75t_L g6312 ( 
.A1(n_4693),
.A2(n_4694),
.B1(n_4920),
.B2(n_4893),
.Y(n_6312)
);

INVx2_ASAP7_75t_SL g6313 ( 
.A(n_5479),
.Y(n_6313)
);

HB1xp67_ASAP7_75t_L g6314 ( 
.A(n_4930),
.Y(n_6314)
);

INVx1_ASAP7_75t_SL g6315 ( 
.A(n_5350),
.Y(n_6315)
);

NAND2xp5_ASAP7_75t_L g6316 ( 
.A(n_5215),
.B(n_4595),
.Y(n_6316)
);

NAND2x1p5_ASAP7_75t_L g6317 ( 
.A(n_5259),
.B(n_4012),
.Y(n_6317)
);

NAND2xp5_ASAP7_75t_L g6318 ( 
.A(n_5215),
.B(n_4595),
.Y(n_6318)
);

OR2x6_ASAP7_75t_L g6319 ( 
.A(n_5081),
.B(n_4514),
.Y(n_6319)
);

AOI22xp33_ASAP7_75t_SL g6320 ( 
.A1(n_5196),
.A2(n_3879),
.B1(n_3988),
.B2(n_3976),
.Y(n_6320)
);

INVxp67_ASAP7_75t_L g6321 ( 
.A(n_5026),
.Y(n_6321)
);

INVx1_ASAP7_75t_L g6322 ( 
.A(n_4898),
.Y(n_6322)
);

OAI21xp33_ASAP7_75t_L g6323 ( 
.A1(n_5380),
.A2(n_4197),
.B(n_4193),
.Y(n_6323)
);

A2O1A1Ixp33_ASAP7_75t_L g6324 ( 
.A1(n_4763),
.A2(n_4056),
.B(n_4087),
.C(n_3988),
.Y(n_6324)
);

NAND2x1p5_ASAP7_75t_L g6325 ( 
.A(n_5259),
.B(n_4012),
.Y(n_6325)
);

O2A1O1Ixp33_ASAP7_75t_L g6326 ( 
.A1(n_4737),
.A2(n_4394),
.B(n_4304),
.C(n_4616),
.Y(n_6326)
);

AND2x2_ASAP7_75t_L g6327 ( 
.A(n_5059),
.B(n_5008),
.Y(n_6327)
);

OAI21x1_ASAP7_75t_L g6328 ( 
.A1(n_5176),
.A2(n_4376),
.B(n_4166),
.Y(n_6328)
);

AOI21xp5_ASAP7_75t_L g6329 ( 
.A1(n_5055),
.A2(n_4033),
.B(n_4026),
.Y(n_6329)
);

NOR2xp33_ASAP7_75t_L g6330 ( 
.A(n_5220),
.B(n_4033),
.Y(n_6330)
);

INVx1_ASAP7_75t_L g6331 ( 
.A(n_4909),
.Y(n_6331)
);

BUFx2_ASAP7_75t_L g6332 ( 
.A(n_5026),
.Y(n_6332)
);

AOI222xp33_ASAP7_75t_L g6333 ( 
.A1(n_4821),
.A2(n_4306),
.B1(n_4307),
.B2(n_4303),
.C1(n_4312),
.C2(n_4299),
.Y(n_6333)
);

NOR2xp33_ASAP7_75t_L g6334 ( 
.A(n_5220),
.B(n_3869),
.Y(n_6334)
);

AOI22xp33_ASAP7_75t_L g6335 ( 
.A1(n_4979),
.A2(n_4558),
.B1(n_4056),
.B2(n_4087),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_4909),
.Y(n_6336)
);

INVx1_ASAP7_75t_L g6337 ( 
.A(n_4910),
.Y(n_6337)
);

INVx1_ASAP7_75t_L g6338 ( 
.A(n_4910),
.Y(n_6338)
);

BUFx2_ASAP7_75t_L g6339 ( 
.A(n_5028),
.Y(n_6339)
);

CKINVDCx5p33_ASAP7_75t_R g6340 ( 
.A(n_4981),
.Y(n_6340)
);

AOI22xp33_ASAP7_75t_L g6341 ( 
.A1(n_4992),
.A2(n_4056),
.B1(n_4087),
.B2(n_4581),
.Y(n_6341)
);

BUFx2_ASAP7_75t_L g6342 ( 
.A(n_5028),
.Y(n_6342)
);

NAND2xp5_ASAP7_75t_L g6343 ( 
.A(n_5242),
.B(n_4609),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_4918),
.Y(n_6344)
);

AOI21xp5_ASAP7_75t_L g6345 ( 
.A1(n_5055),
.A2(n_4394),
.B(n_4304),
.Y(n_6345)
);

BUFx2_ASAP7_75t_L g6346 ( 
.A(n_5028),
.Y(n_6346)
);

AOI21xp5_ASAP7_75t_L g6347 ( 
.A1(n_5056),
.A2(n_4394),
.B(n_4304),
.Y(n_6347)
);

OAI21xp5_ASAP7_75t_L g6348 ( 
.A1(n_4729),
.A2(n_4613),
.B(n_3986),
.Y(n_6348)
);

CKINVDCx5p33_ASAP7_75t_R g6349 ( 
.A(n_4981),
.Y(n_6349)
);

NAND2xp5_ASAP7_75t_L g6350 ( 
.A(n_5242),
.B(n_4609),
.Y(n_6350)
);

OAI21xp5_ASAP7_75t_L g6351 ( 
.A1(n_4729),
.A2(n_4613),
.B(n_3986),
.Y(n_6351)
);

CKINVDCx6p67_ASAP7_75t_R g6352 ( 
.A(n_5469),
.Y(n_6352)
);

AND2x2_ASAP7_75t_L g6353 ( 
.A(n_5008),
.B(n_4261),
.Y(n_6353)
);

NAND2xp5_ASAP7_75t_L g6354 ( 
.A(n_5260),
.B(n_5273),
.Y(n_6354)
);

O2A1O1Ixp5_ASAP7_75t_L g6355 ( 
.A1(n_4812),
.A2(n_3890),
.B(n_3900),
.C(n_3869),
.Y(n_6355)
);

BUFx3_ASAP7_75t_L g6356 ( 
.A(n_5410),
.Y(n_6356)
);

OAI22xp5_ASAP7_75t_L g6357 ( 
.A1(n_4693),
.A2(n_4092),
.B1(n_4103),
.B2(n_4089),
.Y(n_6357)
);

INVx1_ASAP7_75t_SL g6358 ( 
.A(n_5419),
.Y(n_6358)
);

INVx1_ASAP7_75t_L g6359 ( 
.A(n_4918),
.Y(n_6359)
);

NAND2xp5_ASAP7_75t_L g6360 ( 
.A(n_5260),
.B(n_4609),
.Y(n_6360)
);

INVx5_ASAP7_75t_L g6361 ( 
.A(n_5410),
.Y(n_6361)
);

AOI21x1_ASAP7_75t_SL g6362 ( 
.A1(n_4777),
.A2(n_4237),
.B(n_4221),
.Y(n_6362)
);

INVx1_ASAP7_75t_L g6363 ( 
.A(n_4931),
.Y(n_6363)
);

A2O1A1Ixp33_ASAP7_75t_L g6364 ( 
.A1(n_4763),
.A2(n_4087),
.B(n_4056),
.C(n_4666),
.Y(n_6364)
);

AND2x2_ASAP7_75t_L g6365 ( 
.A(n_5008),
.B(n_4264),
.Y(n_6365)
);

NAND2xp5_ASAP7_75t_SL g6366 ( 
.A(n_5158),
.B(n_4086),
.Y(n_6366)
);

INVx4_ASAP7_75t_L g6367 ( 
.A(n_4963),
.Y(n_6367)
);

AND2x2_ASAP7_75t_L g6368 ( 
.A(n_5459),
.B(n_5482),
.Y(n_6368)
);

NAND2xp5_ASAP7_75t_L g6369 ( 
.A(n_5273),
.B(n_4617),
.Y(n_6369)
);

HB1xp67_ASAP7_75t_L g6370 ( 
.A(n_4962),
.Y(n_6370)
);

NAND2xp5_ASAP7_75t_L g6371 ( 
.A(n_5275),
.B(n_4617),
.Y(n_6371)
);

AND2x2_ASAP7_75t_L g6372 ( 
.A(n_5459),
.B(n_4264),
.Y(n_6372)
);

INVx2_ASAP7_75t_SL g6373 ( 
.A(n_5488),
.Y(n_6373)
);

AOI21xp33_ASAP7_75t_L g6374 ( 
.A1(n_5314),
.A2(n_4620),
.B(n_4617),
.Y(n_6374)
);

AOI22xp33_ASAP7_75t_L g6375 ( 
.A1(n_5348),
.A2(n_4994),
.B1(n_4813),
.B2(n_4812),
.Y(n_6375)
);

INVx1_ASAP7_75t_L g6376 ( 
.A(n_4931),
.Y(n_6376)
);

O2A1O1Ixp33_ASAP7_75t_L g6377 ( 
.A1(n_4737),
.A2(n_4394),
.B(n_4304),
.C(n_4616),
.Y(n_6377)
);

INVx1_ASAP7_75t_L g6378 ( 
.A(n_4932),
.Y(n_6378)
);

AOI21xp5_ASAP7_75t_L g6379 ( 
.A1(n_5056),
.A2(n_4613),
.B(n_4237),
.Y(n_6379)
);

INVx1_ASAP7_75t_L g6380 ( 
.A(n_4932),
.Y(n_6380)
);

NAND2x1p5_ASAP7_75t_L g6381 ( 
.A(n_5274),
.B(n_4012),
.Y(n_6381)
);

BUFx2_ASAP7_75t_L g6382 ( 
.A(n_5063),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_4935),
.Y(n_6383)
);

INVx2_ASAP7_75t_SL g6384 ( 
.A(n_5493),
.Y(n_6384)
);

OAI22xp5_ASAP7_75t_L g6385 ( 
.A1(n_4694),
.A2(n_4092),
.B1(n_4103),
.B2(n_4089),
.Y(n_6385)
);

NAND2xp5_ASAP7_75t_SL g6386 ( 
.A(n_5541),
.B(n_4086),
.Y(n_6386)
);

NAND2xp5_ASAP7_75t_L g6387 ( 
.A(n_5275),
.B(n_4620),
.Y(n_6387)
);

NOR2xp33_ASAP7_75t_R g6388 ( 
.A(n_4952),
.B(n_4326),
.Y(n_6388)
);

AOI22xp33_ASAP7_75t_L g6389 ( 
.A1(n_5348),
.A2(n_4581),
.B1(n_4339),
.B2(n_4344),
.Y(n_6389)
);

INVx2_ASAP7_75t_SL g6390 ( 
.A(n_5493),
.Y(n_6390)
);

NAND2xp5_ASAP7_75t_L g6391 ( 
.A(n_5284),
.B(n_4620),
.Y(n_6391)
);

BUFx2_ASAP7_75t_L g6392 ( 
.A(n_5063),
.Y(n_6392)
);

OAI22xp5_ASAP7_75t_L g6393 ( 
.A1(n_4920),
.A2(n_4218),
.B1(n_4272),
.B2(n_4220),
.Y(n_6393)
);

AOI21xp5_ASAP7_75t_L g6394 ( 
.A1(n_5532),
.A2(n_4237),
.B(n_4221),
.Y(n_6394)
);

INVx2_ASAP7_75t_SL g6395 ( 
.A(n_5493),
.Y(n_6395)
);

INVx1_ASAP7_75t_L g6396 ( 
.A(n_4935),
.Y(n_6396)
);

BUFx12f_ASAP7_75t_L g6397 ( 
.A(n_4981),
.Y(n_6397)
);

CKINVDCx16_ASAP7_75t_R g6398 ( 
.A(n_5316),
.Y(n_6398)
);

OAI21x1_ASAP7_75t_L g6399 ( 
.A1(n_4713),
.A2(n_4376),
.B(n_4166),
.Y(n_6399)
);

BUFx2_ASAP7_75t_L g6400 ( 
.A(n_5063),
.Y(n_6400)
);

BUFx2_ASAP7_75t_SL g6401 ( 
.A(n_5541),
.Y(n_6401)
);

NAND2xp5_ASAP7_75t_L g6402 ( 
.A(n_5284),
.B(n_3985),
.Y(n_6402)
);

AOI21xp5_ASAP7_75t_L g6403 ( 
.A1(n_5532),
.A2(n_5015),
.B(n_5418),
.Y(n_6403)
);

AND2x2_ASAP7_75t_L g6404 ( 
.A(n_5459),
.B(n_4265),
.Y(n_6404)
);

BUFx12f_ASAP7_75t_L g6405 ( 
.A(n_5469),
.Y(n_6405)
);

CKINVDCx5p33_ASAP7_75t_R g6406 ( 
.A(n_5241),
.Y(n_6406)
);

INVx1_ASAP7_75t_L g6407 ( 
.A(n_4943),
.Y(n_6407)
);

OAI22xp5_ASAP7_75t_L g6408 ( 
.A1(n_4893),
.A2(n_4220),
.B1(n_4272),
.B2(n_4218),
.Y(n_6408)
);

BUFx2_ASAP7_75t_L g6409 ( 
.A(n_5098),
.Y(n_6409)
);

A2O1A1Ixp33_ASAP7_75t_L g6410 ( 
.A1(n_4699),
.A2(n_5413),
.B(n_5373),
.C(n_5298),
.Y(n_6410)
);

BUFx2_ASAP7_75t_L g6411 ( 
.A(n_5098),
.Y(n_6411)
);

HB1xp67_ASAP7_75t_L g6412 ( 
.A(n_4962),
.Y(n_6412)
);

BUFx3_ASAP7_75t_L g6413 ( 
.A(n_5410),
.Y(n_6413)
);

AOI21xp5_ASAP7_75t_L g6414 ( 
.A1(n_5015),
.A2(n_4240),
.B(n_4221),
.Y(n_6414)
);

HAxp5_ASAP7_75t_L g6415 ( 
.A(n_5314),
.B(n_5263),
.CON(n_6415),
.SN(n_6415)
);

HB1xp67_ASAP7_75t_L g6416 ( 
.A(n_4972),
.Y(n_6416)
);

INVx1_ASAP7_75t_L g6417 ( 
.A(n_4943),
.Y(n_6417)
);

BUFx12f_ASAP7_75t_L g6418 ( 
.A(n_5469),
.Y(n_6418)
);

CKINVDCx5p33_ASAP7_75t_R g6419 ( 
.A(n_5255),
.Y(n_6419)
);

AOI21xp5_ASAP7_75t_SL g6420 ( 
.A1(n_4699),
.A2(n_4875),
.B(n_5354),
.Y(n_6420)
);

AND2x2_ASAP7_75t_L g6421 ( 
.A(n_5482),
.B(n_4265),
.Y(n_6421)
);

AOI21xp5_ASAP7_75t_L g6422 ( 
.A1(n_5418),
.A2(n_4240),
.B(n_4221),
.Y(n_6422)
);

AOI21x1_ASAP7_75t_L g6423 ( 
.A1(n_5052),
.A2(n_4240),
.B(n_4348),
.Y(n_6423)
);

CKINVDCx8_ASAP7_75t_R g6424 ( 
.A(n_5410),
.Y(n_6424)
);

NOR2xp33_ASAP7_75t_L g6425 ( 
.A(n_5295),
.B(n_5297),
.Y(n_6425)
);

AOI21xp5_ASAP7_75t_L g6426 ( 
.A1(n_5418),
.A2(n_4240),
.B(n_4376),
.Y(n_6426)
);

NAND3xp33_ASAP7_75t_L g6427 ( 
.A(n_5354),
.B(n_4000),
.C(n_3993),
.Y(n_6427)
);

INVx6_ASAP7_75t_L g6428 ( 
.A(n_4853),
.Y(n_6428)
);

INVx2_ASAP7_75t_SL g6429 ( 
.A(n_5493),
.Y(n_6429)
);

AOI21xp5_ASAP7_75t_L g6430 ( 
.A1(n_5418),
.A2(n_4240),
.B(n_4376),
.Y(n_6430)
);

BUFx2_ASAP7_75t_R g6431 ( 
.A(n_4724),
.Y(n_6431)
);

INVx1_ASAP7_75t_L g6432 ( 
.A(n_4944),
.Y(n_6432)
);

BUFx3_ASAP7_75t_L g6433 ( 
.A(n_5410),
.Y(n_6433)
);

AOI221xp5_ASAP7_75t_L g6434 ( 
.A1(n_5319),
.A2(n_4295),
.B1(n_4299),
.B2(n_4284),
.C(n_4283),
.Y(n_6434)
);

INVx1_ASAP7_75t_SL g6435 ( 
.A(n_5419),
.Y(n_6435)
);

INVx1_ASAP7_75t_SL g6436 ( 
.A(n_5440),
.Y(n_6436)
);

INVx3_ASAP7_75t_L g6437 ( 
.A(n_5142),
.Y(n_6437)
);

NAND2xp5_ASAP7_75t_L g6438 ( 
.A(n_5295),
.B(n_3993),
.Y(n_6438)
);

OAI222xp33_ASAP7_75t_L g6439 ( 
.A1(n_5328),
.A2(n_5274),
.B1(n_4727),
.B2(n_5524),
.C1(n_5298),
.C2(n_5337),
.Y(n_6439)
);

INVx1_ASAP7_75t_L g6440 ( 
.A(n_4944),
.Y(n_6440)
);

AOI22xp33_ASAP7_75t_L g6441 ( 
.A1(n_4994),
.A2(n_4581),
.B1(n_4339),
.B2(n_4344),
.Y(n_6441)
);

INVx1_ASAP7_75t_L g6442 ( 
.A(n_6144),
.Y(n_6442)
);

OA21x2_ASAP7_75t_L g6443 ( 
.A1(n_6403),
.A2(n_5270),
.B(n_5417),
.Y(n_6443)
);

OAI21x1_ASAP7_75t_L g6444 ( 
.A1(n_6097),
.A2(n_5285),
.B(n_5270),
.Y(n_6444)
);

AOI21xp5_ASAP7_75t_L g6445 ( 
.A1(n_5770),
.A2(n_5418),
.B(n_4800),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_6144),
.Y(n_6446)
);

NAND2xp5_ASAP7_75t_L g6447 ( 
.A(n_5560),
.B(n_5098),
.Y(n_6447)
);

AND2x2_ASAP7_75t_L g6448 ( 
.A(n_5713),
.B(n_5482),
.Y(n_6448)
);

AO21x1_ASAP7_75t_L g6449 ( 
.A1(n_5682),
.A2(n_5358),
.B(n_4965),
.Y(n_6449)
);

OAI21x1_ASAP7_75t_L g6450 ( 
.A1(n_6097),
.A2(n_5285),
.B(n_4750),
.Y(n_6450)
);

NOR2xp33_ASAP7_75t_L g6451 ( 
.A(n_5705),
.B(n_5682),
.Y(n_6451)
);

NAND2xp5_ASAP7_75t_L g6452 ( 
.A(n_5560),
.B(n_5115),
.Y(n_6452)
);

OR2x2_ASAP7_75t_L g6453 ( 
.A(n_5654),
.B(n_5115),
.Y(n_6453)
);

AO31x2_ASAP7_75t_L g6454 ( 
.A1(n_6117),
.A2(n_5344),
.A3(n_5000),
.B(n_5023),
.Y(n_6454)
);

INVx2_ASAP7_75t_L g6455 ( 
.A(n_5553),
.Y(n_6455)
);

BUFx2_ASAP7_75t_L g6456 ( 
.A(n_6128),
.Y(n_6456)
);

BUFx2_ASAP7_75t_L g6457 ( 
.A(n_6128),
.Y(n_6457)
);

INVx6_ASAP7_75t_L g6458 ( 
.A(n_6246),
.Y(n_6458)
);

INVx1_ASAP7_75t_L g6459 ( 
.A(n_6154),
.Y(n_6459)
);

OAI21x1_ASAP7_75t_L g6460 ( 
.A1(n_6097),
.A2(n_5285),
.B(n_4750),
.Y(n_6460)
);

AOI22xp33_ASAP7_75t_L g6461 ( 
.A1(n_5664),
.A2(n_5196),
.B1(n_4869),
.B2(n_4826),
.Y(n_6461)
);

AO31x2_ASAP7_75t_L g6462 ( 
.A1(n_6117),
.A2(n_5344),
.A3(n_5023),
.B(n_5358),
.Y(n_6462)
);

AOI21xp5_ASAP7_75t_L g6463 ( 
.A1(n_5770),
.A2(n_5418),
.B(n_4983),
.Y(n_6463)
);

INVx1_ASAP7_75t_L g6464 ( 
.A(n_6154),
.Y(n_6464)
);

OA21x2_ASAP7_75t_L g6465 ( 
.A1(n_6403),
.A2(n_5065),
.B(n_5052),
.Y(n_6465)
);

INVx1_ASAP7_75t_L g6466 ( 
.A(n_6157),
.Y(n_6466)
);

OAI21xp33_ASAP7_75t_SL g6467 ( 
.A1(n_5575),
.A2(n_5140),
.B(n_5184),
.Y(n_6467)
);

INVx6_ASAP7_75t_L g6468 ( 
.A(n_6246),
.Y(n_6468)
);

NAND2xp5_ASAP7_75t_L g6469 ( 
.A(n_5672),
.B(n_5115),
.Y(n_6469)
);

AO21x2_ASAP7_75t_L g6470 ( 
.A1(n_5894),
.A2(n_5037),
.B(n_5030),
.Y(n_6470)
);

INVx2_ASAP7_75t_L g6471 ( 
.A(n_5553),
.Y(n_6471)
);

OAI21x1_ASAP7_75t_L g6472 ( 
.A1(n_6423),
.A2(n_4750),
.B(n_5426),
.Y(n_6472)
);

INVx2_ASAP7_75t_SL g6473 ( 
.A(n_6246),
.Y(n_6473)
);

OAI21x1_ASAP7_75t_L g6474 ( 
.A1(n_6423),
.A2(n_5426),
.B(n_5289),
.Y(n_6474)
);

OR2x2_ASAP7_75t_L g6475 ( 
.A(n_5654),
.B(n_5124),
.Y(n_6475)
);

OAI21x1_ASAP7_75t_L g6476 ( 
.A1(n_6423),
.A2(n_6300),
.B(n_6170),
.Y(n_6476)
);

NAND2x1p5_ASAP7_75t_L g6477 ( 
.A(n_5598),
.B(n_4963),
.Y(n_6477)
);

NAND2x1p5_ASAP7_75t_L g6478 ( 
.A(n_5598),
.B(n_4963),
.Y(n_6478)
);

INVx2_ASAP7_75t_L g6479 ( 
.A(n_5553),
.Y(n_6479)
);

OAI221xp5_ASAP7_75t_L g6480 ( 
.A1(n_5951),
.A2(n_5337),
.B1(n_5380),
.B2(n_5442),
.C(n_5413),
.Y(n_6480)
);

BUFx2_ASAP7_75t_L g6481 ( 
.A(n_6128),
.Y(n_6481)
);

INVx1_ASAP7_75t_L g6482 ( 
.A(n_6157),
.Y(n_6482)
);

OAI21x1_ASAP7_75t_L g6483 ( 
.A1(n_6170),
.A2(n_5289),
.B(n_4742),
.Y(n_6483)
);

NOR2xp33_ASAP7_75t_L g6484 ( 
.A(n_5705),
.B(n_5359),
.Y(n_6484)
);

INVx1_ASAP7_75t_L g6485 ( 
.A(n_6159),
.Y(n_6485)
);

OAI21x1_ASAP7_75t_L g6486 ( 
.A1(n_6170),
.A2(n_5289),
.B(n_4742),
.Y(n_6486)
);

AND2x2_ASAP7_75t_L g6487 ( 
.A(n_5713),
.B(n_5499),
.Y(n_6487)
);

INVx2_ASAP7_75t_L g6488 ( 
.A(n_5553),
.Y(n_6488)
);

HB1xp67_ASAP7_75t_L g6489 ( 
.A(n_5812),
.Y(n_6489)
);

NAND2x1p5_ASAP7_75t_L g6490 ( 
.A(n_5598),
.B(n_4963),
.Y(n_6490)
);

INVx6_ASAP7_75t_L g6491 ( 
.A(n_6246),
.Y(n_6491)
);

AOI22xp33_ASAP7_75t_L g6492 ( 
.A1(n_5664),
.A2(n_4826),
.B1(n_4813),
.B2(n_5359),
.Y(n_6492)
);

AO21x2_ASAP7_75t_L g6493 ( 
.A1(n_5894),
.A2(n_5037),
.B(n_5030),
.Y(n_6493)
);

HB1xp67_ASAP7_75t_L g6494 ( 
.A(n_5812),
.Y(n_6494)
);

INVx1_ASAP7_75t_L g6495 ( 
.A(n_6159),
.Y(n_6495)
);

INVx3_ASAP7_75t_L g6496 ( 
.A(n_5636),
.Y(n_6496)
);

AND2x4_ASAP7_75t_L g6497 ( 
.A(n_5822),
.B(n_5493),
.Y(n_6497)
);

INVx1_ASAP7_75t_L g6498 ( 
.A(n_6173),
.Y(n_6498)
);

AO31x2_ASAP7_75t_L g6499 ( 
.A1(n_6117),
.A2(n_4961),
.A3(n_5517),
.B(n_5514),
.Y(n_6499)
);

OA21x2_ASAP7_75t_L g6500 ( 
.A1(n_5579),
.A2(n_5072),
.B(n_5065),
.Y(n_6500)
);

OAI21x1_ASAP7_75t_L g6501 ( 
.A1(n_6300),
.A2(n_4713),
.B(n_5072),
.Y(n_6501)
);

CKINVDCx5p33_ASAP7_75t_R g6502 ( 
.A(n_5619),
.Y(n_6502)
);

NOR2xp67_ASAP7_75t_L g6503 ( 
.A(n_6246),
.B(n_6257),
.Y(n_6503)
);

OAI21x1_ASAP7_75t_L g6504 ( 
.A1(n_6300),
.A2(n_5089),
.B(n_5079),
.Y(n_6504)
);

OAI22xp5_ASAP7_75t_L g6505 ( 
.A1(n_6006),
.A2(n_5442),
.B1(n_5124),
.B2(n_4833),
.Y(n_6505)
);

INVx4_ASAP7_75t_SL g6506 ( 
.A(n_5573),
.Y(n_6506)
);

NAND2xp5_ASAP7_75t_L g6507 ( 
.A(n_5672),
.B(n_5124),
.Y(n_6507)
);

BUFx2_ASAP7_75t_L g6508 ( 
.A(n_5670),
.Y(n_6508)
);

AND2x2_ASAP7_75t_L g6509 ( 
.A(n_5713),
.B(n_5499),
.Y(n_6509)
);

OA21x2_ASAP7_75t_L g6510 ( 
.A1(n_5579),
.A2(n_5089),
.B(n_5079),
.Y(n_6510)
);

OAI21x1_ASAP7_75t_L g6511 ( 
.A1(n_6298),
.A2(n_5129),
.B(n_5116),
.Y(n_6511)
);

INVx1_ASAP7_75t_L g6512 ( 
.A(n_6173),
.Y(n_6512)
);

BUFx6f_ASAP7_75t_L g6513 ( 
.A(n_5598),
.Y(n_6513)
);

OAI22xp5_ASAP7_75t_L g6514 ( 
.A1(n_6006),
.A2(n_4833),
.B1(n_4915),
.B2(n_4908),
.Y(n_6514)
);

O2A1O1Ixp33_ASAP7_75t_SL g6515 ( 
.A1(n_5951),
.A2(n_5263),
.B(n_4952),
.C(n_5422),
.Y(n_6515)
);

AOI21x1_ASAP7_75t_L g6516 ( 
.A1(n_5572),
.A2(n_5140),
.B(n_5311),
.Y(n_6516)
);

INVx1_ASAP7_75t_L g6517 ( 
.A(n_6183),
.Y(n_6517)
);

INVx1_ASAP7_75t_L g6518 ( 
.A(n_6183),
.Y(n_6518)
);

BUFx3_ASAP7_75t_L g6519 ( 
.A(n_5628),
.Y(n_6519)
);

BUFx3_ASAP7_75t_L g6520 ( 
.A(n_5628),
.Y(n_6520)
);

AO32x2_ASAP7_75t_L g6521 ( 
.A1(n_6039),
.A2(n_5303),
.A3(n_5306),
.B1(n_5277),
.B2(n_5261),
.Y(n_6521)
);

OAI21x1_ASAP7_75t_L g6522 ( 
.A1(n_6298),
.A2(n_5129),
.B(n_5116),
.Y(n_6522)
);

OAI21x1_ASAP7_75t_L g6523 ( 
.A1(n_6345),
.A2(n_5164),
.B(n_5143),
.Y(n_6523)
);

INVx2_ASAP7_75t_L g6524 ( 
.A(n_5555),
.Y(n_6524)
);

OAI21x1_ASAP7_75t_L g6525 ( 
.A1(n_6345),
.A2(n_5164),
.B(n_5143),
.Y(n_6525)
);

OAI21x1_ASAP7_75t_L g6526 ( 
.A1(n_6347),
.A2(n_5462),
.B(n_5311),
.Y(n_6526)
);

OAI21x1_ASAP7_75t_L g6527 ( 
.A1(n_6347),
.A2(n_5462),
.B(n_4967),
.Y(n_6527)
);

INVx3_ASAP7_75t_L g6528 ( 
.A(n_5636),
.Y(n_6528)
);

NAND2xp5_ASAP7_75t_SL g6529 ( 
.A(n_5629),
.B(n_4963),
.Y(n_6529)
);

INVx2_ASAP7_75t_L g6530 ( 
.A(n_5555),
.Y(n_6530)
);

AOI22xp33_ASAP7_75t_SL g6531 ( 
.A1(n_6116),
.A2(n_6210),
.B1(n_6174),
.B2(n_6005),
.Y(n_6531)
);

OAI21x1_ASAP7_75t_L g6532 ( 
.A1(n_6082),
.A2(n_5462),
.B(n_4967),
.Y(n_6532)
);

NAND2xp5_ASAP7_75t_L g6533 ( 
.A(n_5672),
.B(n_5401),
.Y(n_6533)
);

BUFx3_ASAP7_75t_L g6534 ( 
.A(n_5628),
.Y(n_6534)
);

OAI21x1_ASAP7_75t_L g6535 ( 
.A1(n_6082),
.A2(n_4941),
.B(n_4864),
.Y(n_6535)
);

AOI22xp33_ASAP7_75t_L g6536 ( 
.A1(n_5809),
.A2(n_6116),
.B1(n_6210),
.B2(n_6005),
.Y(n_6536)
);

OAI21x1_ASAP7_75t_L g6537 ( 
.A1(n_6090),
.A2(n_4941),
.B(n_4864),
.Y(n_6537)
);

CKINVDCx11_ASAP7_75t_R g6538 ( 
.A(n_5867),
.Y(n_6538)
);

INVx4_ASAP7_75t_L g6539 ( 
.A(n_5548),
.Y(n_6539)
);

AND2x4_ASAP7_75t_L g6540 ( 
.A(n_5822),
.B(n_5526),
.Y(n_6540)
);

NOR2xp33_ASAP7_75t_L g6541 ( 
.A(n_5632),
.B(n_5297),
.Y(n_6541)
);

HB1xp67_ASAP7_75t_L g6542 ( 
.A(n_5816),
.Y(n_6542)
);

OAI21xp5_ASAP7_75t_L g6543 ( 
.A1(n_5975),
.A2(n_5184),
.B(n_4802),
.Y(n_6543)
);

BUFx3_ASAP7_75t_L g6544 ( 
.A(n_5628),
.Y(n_6544)
);

AND2x2_ASAP7_75t_L g6545 ( 
.A(n_5730),
.B(n_5499),
.Y(n_6545)
);

BUFx2_ASAP7_75t_L g6546 ( 
.A(n_5670),
.Y(n_6546)
);

INVx2_ASAP7_75t_L g6547 ( 
.A(n_5555),
.Y(n_6547)
);

INVx1_ASAP7_75t_L g6548 ( 
.A(n_6184),
.Y(n_6548)
);

AOI22xp33_ASAP7_75t_L g6549 ( 
.A1(n_5809),
.A2(n_5940),
.B1(n_5938),
.B2(n_5632),
.Y(n_6549)
);

AO21x2_ASAP7_75t_L g6550 ( 
.A1(n_5920),
.A2(n_5030),
.B(n_4983),
.Y(n_6550)
);

OAI21xp5_ASAP7_75t_L g6551 ( 
.A1(n_5975),
.A2(n_4802),
.B(n_5389),
.Y(n_6551)
);

NAND2xp5_ASAP7_75t_L g6552 ( 
.A(n_5912),
.B(n_5401),
.Y(n_6552)
);

HB1xp67_ASAP7_75t_L g6553 ( 
.A(n_5816),
.Y(n_6553)
);

INVx1_ASAP7_75t_L g6554 ( 
.A(n_6184),
.Y(n_6554)
);

INVx1_ASAP7_75t_L g6555 ( 
.A(n_6187),
.Y(n_6555)
);

AO31x2_ASAP7_75t_L g6556 ( 
.A1(n_5730),
.A2(n_4961),
.A3(n_5517),
.B(n_5514),
.Y(n_6556)
);

INVx2_ASAP7_75t_SL g6557 ( 
.A(n_6246),
.Y(n_6557)
);

NAND2xp5_ASAP7_75t_L g6558 ( 
.A(n_5912),
.B(n_5411),
.Y(n_6558)
);

AO21x2_ASAP7_75t_L g6559 ( 
.A1(n_5920),
.A2(n_5030),
.B(n_5007),
.Y(n_6559)
);

INVx1_ASAP7_75t_L g6560 ( 
.A(n_6187),
.Y(n_6560)
);

INVx2_ASAP7_75t_L g6561 ( 
.A(n_5555),
.Y(n_6561)
);

OAI21x1_ASAP7_75t_L g6562 ( 
.A1(n_6090),
.A2(n_4824),
.B(n_4823),
.Y(n_6562)
);

OAI22xp33_ASAP7_75t_L g6563 ( 
.A1(n_6014),
.A2(n_5524),
.B1(n_5328),
.B2(n_5522),
.Y(n_6563)
);

INVxp67_ASAP7_75t_SL g6564 ( 
.A(n_5959),
.Y(n_6564)
);

NOR2xp67_ASAP7_75t_SL g6565 ( 
.A(n_5548),
.B(n_5477),
.Y(n_6565)
);

AOI22xp5_ASAP7_75t_L g6566 ( 
.A1(n_6014),
.A2(n_5522),
.B1(n_4929),
.B2(n_4831),
.Y(n_6566)
);

AOI21xp33_ASAP7_75t_L g6567 ( 
.A1(n_5938),
.A2(n_5389),
.B(n_4946),
.Y(n_6567)
);

INVx5_ASAP7_75t_SL g6568 ( 
.A(n_6352),
.Y(n_6568)
);

BUFx2_ASAP7_75t_L g6569 ( 
.A(n_5670),
.Y(n_6569)
);

AOI22xp33_ASAP7_75t_L g6570 ( 
.A1(n_5940),
.A2(n_5224),
.B1(n_4831),
.B2(n_4929),
.Y(n_6570)
);

OAI21xp5_ASAP7_75t_L g6571 ( 
.A1(n_6420),
.A2(n_4875),
.B(n_4895),
.Y(n_6571)
);

OAI21x1_ASAP7_75t_L g6572 ( 
.A1(n_6100),
.A2(n_6111),
.B(n_6107),
.Y(n_6572)
);

OAI21x1_ASAP7_75t_SL g6573 ( 
.A1(n_5543),
.A2(n_5310),
.B(n_5188),
.Y(n_6573)
);

BUFx3_ASAP7_75t_L g6574 ( 
.A(n_5548),
.Y(n_6574)
);

INVx1_ASAP7_75t_L g6575 ( 
.A(n_6189),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_6189),
.Y(n_6576)
);

OAI21x1_ASAP7_75t_L g6577 ( 
.A1(n_6100),
.A2(n_4824),
.B(n_4823),
.Y(n_6577)
);

NAND2x1_ASAP7_75t_L g6578 ( 
.A(n_6104),
.B(n_5114),
.Y(n_6578)
);

OAI21x1_ASAP7_75t_L g6579 ( 
.A1(n_6107),
.A2(n_6119),
.B(n_6111),
.Y(n_6579)
);

OAI222xp33_ASAP7_75t_L g6580 ( 
.A1(n_6099),
.A2(n_5483),
.B1(n_5484),
.B2(n_5081),
.C1(n_5266),
.C2(n_5542),
.Y(n_6580)
);

NAND2x1_ASAP7_75t_L g6581 ( 
.A(n_6104),
.B(n_5114),
.Y(n_6581)
);

HB1xp67_ASAP7_75t_L g6582 ( 
.A(n_5848),
.Y(n_6582)
);

A2O1A1Ixp33_ASAP7_75t_L g6583 ( 
.A1(n_6174),
.A2(n_6410),
.B(n_6099),
.C(n_5693),
.Y(n_6583)
);

INVx3_ASAP7_75t_L g6584 ( 
.A(n_5636),
.Y(n_6584)
);

OR2x2_ASAP7_75t_L g6585 ( 
.A(n_5654),
.B(n_5421),
.Y(n_6585)
);

NAND3x1_ASAP7_75t_L g6586 ( 
.A(n_5806),
.B(n_5483),
.C(n_4905),
.Y(n_6586)
);

OAI22xp5_ASAP7_75t_L g6587 ( 
.A1(n_5570),
.A2(n_4915),
.B1(n_4908),
.B2(n_5353),
.Y(n_6587)
);

OAI21x1_ASAP7_75t_L g6588 ( 
.A1(n_6119),
.A2(n_4876),
.B(n_4873),
.Y(n_6588)
);

INVx2_ASAP7_75t_L g6589 ( 
.A(n_5562),
.Y(n_6589)
);

INVx1_ASAP7_75t_L g6590 ( 
.A(n_6190),
.Y(n_6590)
);

AND2x2_ASAP7_75t_L g6591 ( 
.A(n_5730),
.B(n_5503),
.Y(n_6591)
);

HB1xp67_ASAP7_75t_L g6592 ( 
.A(n_5848),
.Y(n_6592)
);

INVx1_ASAP7_75t_SL g6593 ( 
.A(n_5748),
.Y(n_6593)
);

OAI21x1_ASAP7_75t_L g6594 ( 
.A1(n_6120),
.A2(n_4876),
.B(n_4873),
.Y(n_6594)
);

OAI21xp5_ASAP7_75t_L g6595 ( 
.A1(n_6410),
.A2(n_4895),
.B(n_4734),
.Y(n_6595)
);

OAI21xp5_ASAP7_75t_L g6596 ( 
.A1(n_5862),
.A2(n_4734),
.B(n_4916),
.Y(n_6596)
);

INVx1_ASAP7_75t_L g6597 ( 
.A(n_6190),
.Y(n_6597)
);

INVx3_ASAP7_75t_L g6598 ( 
.A(n_5636),
.Y(n_6598)
);

OAI211xp5_ASAP7_75t_L g6599 ( 
.A1(n_5575),
.A2(n_4815),
.B(n_4905),
.C(n_4897),
.Y(n_6599)
);

BUFx2_ASAP7_75t_L g6600 ( 
.A(n_5670),
.Y(n_6600)
);

AOI21xp5_ASAP7_75t_L g6601 ( 
.A1(n_6247),
.A2(n_5418),
.B(n_4863),
.Y(n_6601)
);

OAI21x1_ASAP7_75t_L g6602 ( 
.A1(n_6120),
.A2(n_4706),
.B(n_5456),
.Y(n_6602)
);

OAI22xp33_ASAP7_75t_SL g6603 ( 
.A1(n_6155),
.A2(n_4928),
.B1(n_5006),
.B2(n_4870),
.Y(n_6603)
);

OAI21x1_ASAP7_75t_L g6604 ( 
.A1(n_6232),
.A2(n_4706),
.B(n_5456),
.Y(n_6604)
);

OAI21x1_ASAP7_75t_L g6605 ( 
.A1(n_6232),
.A2(n_5480),
.B(n_5467),
.Y(n_6605)
);

AOI21xp5_ASAP7_75t_L g6606 ( 
.A1(n_6247),
.A2(n_4863),
.B(n_5373),
.Y(n_6606)
);

AOI21xp5_ASAP7_75t_L g6607 ( 
.A1(n_5563),
.A2(n_5423),
.B(n_5409),
.Y(n_6607)
);

AOI22xp33_ASAP7_75t_L g6608 ( 
.A1(n_5693),
.A2(n_5224),
.B1(n_4977),
.B2(n_4815),
.Y(n_6608)
);

NAND2xp5_ASAP7_75t_L g6609 ( 
.A(n_5918),
.B(n_5411),
.Y(n_6609)
);

INVx2_ASAP7_75t_L g6610 ( 
.A(n_5562),
.Y(n_6610)
);

AOI22xp33_ASAP7_75t_L g6611 ( 
.A1(n_5806),
.A2(n_5224),
.B1(n_4977),
.B2(n_4926),
.Y(n_6611)
);

INVx1_ASAP7_75t_L g6612 ( 
.A(n_6196),
.Y(n_6612)
);

NAND3xp33_ASAP7_75t_L g6613 ( 
.A(n_6023),
.B(n_4897),
.C(n_5388),
.Y(n_6613)
);

NAND2x1p5_ASAP7_75t_L g6614 ( 
.A(n_5598),
.B(n_5114),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_6196),
.Y(n_6615)
);

OA21x2_ASAP7_75t_L g6616 ( 
.A1(n_6422),
.A2(n_5423),
.B(n_5007),
.Y(n_6616)
);

OR2x6_ASAP7_75t_L g6617 ( 
.A(n_6244),
.B(n_5081),
.Y(n_6617)
);

AOI22xp33_ASAP7_75t_L g6618 ( 
.A1(n_6231),
.A2(n_5626),
.B1(n_5708),
.B2(n_6375),
.Y(n_6618)
);

AOI22xp33_ASAP7_75t_SL g6619 ( 
.A1(n_5778),
.A2(n_5224),
.B1(n_5378),
.B2(n_5476),
.Y(n_6619)
);

AND2x2_ASAP7_75t_L g6620 ( 
.A(n_5778),
.B(n_5503),
.Y(n_6620)
);

INVx1_ASAP7_75t_L g6621 ( 
.A(n_6201),
.Y(n_6621)
);

BUFx3_ASAP7_75t_L g6622 ( 
.A(n_5548),
.Y(n_6622)
);

OAI22xp33_ASAP7_75t_L g6623 ( 
.A1(n_6155),
.A2(n_5501),
.B1(n_5353),
.B2(n_5188),
.Y(n_6623)
);

INVx1_ASAP7_75t_L g6624 ( 
.A(n_6201),
.Y(n_6624)
);

OR2x6_ASAP7_75t_L g6625 ( 
.A(n_6244),
.B(n_5081),
.Y(n_6625)
);

INVx2_ASAP7_75t_L g6626 ( 
.A(n_5562),
.Y(n_6626)
);

INVx2_ASAP7_75t_L g6627 ( 
.A(n_5562),
.Y(n_6627)
);

AND2x4_ASAP7_75t_L g6628 ( 
.A(n_5822),
.B(n_5526),
.Y(n_6628)
);

OAI21x1_ASAP7_75t_L g6629 ( 
.A1(n_6287),
.A2(n_5480),
.B(n_5467),
.Y(n_6629)
);

OAI21x1_ASAP7_75t_L g6630 ( 
.A1(n_6287),
.A2(n_5485),
.B(n_5481),
.Y(n_6630)
);

OAI21x1_ASAP7_75t_L g6631 ( 
.A1(n_6299),
.A2(n_5485),
.B(n_5481),
.Y(n_6631)
);

INVx4_ASAP7_75t_L g6632 ( 
.A(n_5589),
.Y(n_6632)
);

INVx1_ASAP7_75t_L g6633 ( 
.A(n_6203),
.Y(n_6633)
);

OAI21x1_ASAP7_75t_L g6634 ( 
.A1(n_6299),
.A2(n_4837),
.B(n_4838),
.Y(n_6634)
);

AOI22xp33_ASAP7_75t_L g6635 ( 
.A1(n_6231),
.A2(n_5224),
.B1(n_4926),
.B2(n_4882),
.Y(n_6635)
);

INVx1_ASAP7_75t_L g6636 ( 
.A(n_6203),
.Y(n_6636)
);

NAND2xp5_ASAP7_75t_L g6637 ( 
.A(n_5918),
.B(n_5416),
.Y(n_6637)
);

OAI21x1_ASAP7_75t_L g6638 ( 
.A1(n_5572),
.A2(n_4837),
.B(n_4838),
.Y(n_6638)
);

AND2x2_ASAP7_75t_L g6639 ( 
.A(n_5778),
.B(n_5503),
.Y(n_6639)
);

INVx4_ASAP7_75t_L g6640 ( 
.A(n_5589),
.Y(n_6640)
);

BUFx3_ASAP7_75t_L g6641 ( 
.A(n_5942),
.Y(n_6641)
);

INVx3_ASAP7_75t_L g6642 ( 
.A(n_5636),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6205),
.Y(n_6643)
);

OA21x2_ASAP7_75t_L g6644 ( 
.A1(n_6422),
.A2(n_5388),
.B(n_5034),
.Y(n_6644)
);

NOR2xp33_ASAP7_75t_L g6645 ( 
.A(n_6023),
.B(n_5300),
.Y(n_6645)
);

INVx3_ASAP7_75t_L g6646 ( 
.A(n_5670),
.Y(n_6646)
);

OAI22xp33_ASAP7_75t_L g6647 ( 
.A1(n_5723),
.A2(n_5501),
.B1(n_5353),
.B2(n_5188),
.Y(n_6647)
);

AOI22xp33_ASAP7_75t_L g6648 ( 
.A1(n_5626),
.A2(n_4882),
.B1(n_4937),
.B2(n_5490),
.Y(n_6648)
);

NAND2xp5_ASAP7_75t_L g6649 ( 
.A(n_5585),
.B(n_5416),
.Y(n_6649)
);

AOI21xp5_ASAP7_75t_L g6650 ( 
.A1(n_5563),
.A2(n_5409),
.B(n_5402),
.Y(n_6650)
);

AO21x1_ASAP7_75t_L g6651 ( 
.A1(n_6032),
.A2(n_5452),
.B(n_5448),
.Y(n_6651)
);

OAI211xp5_ASAP7_75t_SL g6652 ( 
.A1(n_5739),
.A2(n_5422),
.B(n_4878),
.C(n_5447),
.Y(n_6652)
);

AND2x6_ASAP7_75t_L g6653 ( 
.A(n_5554),
.B(n_4870),
.Y(n_6653)
);

INVx2_ASAP7_75t_L g6654 ( 
.A(n_5567),
.Y(n_6654)
);

NOR2xp33_ASAP7_75t_L g6655 ( 
.A(n_6032),
.B(n_5300),
.Y(n_6655)
);

AOI21xp5_ASAP7_75t_L g6656 ( 
.A1(n_6213),
.A2(n_5402),
.B(n_5398),
.Y(n_6656)
);

AOI22xp33_ASAP7_75t_SL g6657 ( 
.A1(n_5788),
.A2(n_5476),
.B1(n_4959),
.B2(n_5035),
.Y(n_6657)
);

INVx1_ASAP7_75t_L g6658 ( 
.A(n_6205),
.Y(n_6658)
);

OAI21x1_ASAP7_75t_L g6659 ( 
.A1(n_5572),
.A2(n_4950),
.B(n_5465),
.Y(n_6659)
);

OAI22xp5_ASAP7_75t_SL g6660 ( 
.A1(n_5760),
.A2(n_5414),
.B1(n_5173),
.B2(n_5336),
.Y(n_6660)
);

BUFx3_ASAP7_75t_L g6661 ( 
.A(n_5942),
.Y(n_6661)
);

OAI21x1_ASAP7_75t_L g6662 ( 
.A1(n_5552),
.A2(n_4950),
.B(n_5465),
.Y(n_6662)
);

CKINVDCx5p33_ASAP7_75t_R g6663 ( 
.A(n_5619),
.Y(n_6663)
);

AOI21xp33_ASAP7_75t_L g6664 ( 
.A1(n_6427),
.A2(n_4946),
.B(n_5448),
.Y(n_6664)
);

BUFx10_ASAP7_75t_L g6665 ( 
.A(n_6018),
.Y(n_6665)
);

NAND2xp5_ASAP7_75t_L g6666 ( 
.A(n_5585),
.B(n_5305),
.Y(n_6666)
);

BUFx12f_ASAP7_75t_L g6667 ( 
.A(n_5914),
.Y(n_6667)
);

OAI21x1_ASAP7_75t_L g6668 ( 
.A1(n_5552),
.A2(n_5777),
.B(n_5620),
.Y(n_6668)
);

AO21x2_ASAP7_75t_L g6669 ( 
.A1(n_5920),
.A2(n_6056),
.B(n_6292),
.Y(n_6669)
);

OAI21x1_ASAP7_75t_L g6670 ( 
.A1(n_5552),
.A2(n_5474),
.B(n_5465),
.Y(n_6670)
);

OAI21x1_ASAP7_75t_L g6671 ( 
.A1(n_5620),
.A2(n_5474),
.B(n_5465),
.Y(n_6671)
);

BUFx2_ASAP7_75t_L g6672 ( 
.A(n_5549),
.Y(n_6672)
);

AOI21xp5_ASAP7_75t_L g6673 ( 
.A1(n_6213),
.A2(n_5708),
.B(n_6197),
.Y(n_6673)
);

HB1xp67_ASAP7_75t_L g6674 ( 
.A(n_5890),
.Y(n_6674)
);

OAI21x1_ASAP7_75t_L g6675 ( 
.A1(n_5620),
.A2(n_5498),
.B(n_5474),
.Y(n_6675)
);

AOI21xp5_ASAP7_75t_L g6676 ( 
.A1(n_6197),
.A2(n_5398),
.B(n_4791),
.Y(n_6676)
);

INVx1_ASAP7_75t_L g6677 ( 
.A(n_6208),
.Y(n_6677)
);

OAI21xp5_ASAP7_75t_L g6678 ( 
.A1(n_6427),
.A2(n_4916),
.B(n_4780),
.Y(n_6678)
);

INVx3_ASAP7_75t_L g6679 ( 
.A(n_5641),
.Y(n_6679)
);

CKINVDCx6p67_ASAP7_75t_R g6680 ( 
.A(n_5698),
.Y(n_6680)
);

INVx1_ASAP7_75t_L g6681 ( 
.A(n_6208),
.Y(n_6681)
);

INVx2_ASAP7_75t_L g6682 ( 
.A(n_5567),
.Y(n_6682)
);

BUFx3_ASAP7_75t_L g6683 ( 
.A(n_5942),
.Y(n_6683)
);

OAI21x1_ASAP7_75t_SL g6684 ( 
.A1(n_5543),
.A2(n_5310),
.B(n_5188),
.Y(n_6684)
);

OAI21x1_ASAP7_75t_L g6685 ( 
.A1(n_5777),
.A2(n_5498),
.B(n_4878),
.Y(n_6685)
);

AOI21xp5_ASAP7_75t_L g6686 ( 
.A1(n_6326),
.A2(n_4791),
.B(n_4948),
.Y(n_6686)
);

NAND2xp33_ASAP7_75t_L g6687 ( 
.A(n_5754),
.B(n_4959),
.Y(n_6687)
);

OAI21x1_ASAP7_75t_L g6688 ( 
.A1(n_6426),
.A2(n_5498),
.B(n_4844),
.Y(n_6688)
);

INVx1_ASAP7_75t_L g6689 ( 
.A(n_6248),
.Y(n_6689)
);

INVx1_ASAP7_75t_SL g6690 ( 
.A(n_5748),
.Y(n_6690)
);

AND2x4_ASAP7_75t_L g6691 ( 
.A(n_5822),
.B(n_5526),
.Y(n_6691)
);

INVx2_ASAP7_75t_SL g6692 ( 
.A(n_6246),
.Y(n_6692)
);

OR2x2_ASAP7_75t_L g6693 ( 
.A(n_5892),
.B(n_5421),
.Y(n_6693)
);

OA21x2_ASAP7_75t_L g6694 ( 
.A1(n_6426),
.A2(n_5034),
.B(n_4711),
.Y(n_6694)
);

NOR2xp33_ASAP7_75t_L g6695 ( 
.A(n_5977),
.B(n_5305),
.Y(n_6695)
);

A2O1A1Ixp33_ASAP7_75t_L g6696 ( 
.A1(n_6326),
.A2(n_4948),
.B(n_4780),
.C(n_4928),
.Y(n_6696)
);

NAND2xp5_ASAP7_75t_L g6697 ( 
.A(n_5616),
.B(n_5313),
.Y(n_6697)
);

AOI22xp33_ASAP7_75t_L g6698 ( 
.A1(n_6375),
.A2(n_4937),
.B1(n_5520),
.B2(n_5490),
.Y(n_6698)
);

AOI222xp33_ASAP7_75t_L g6699 ( 
.A1(n_6042),
.A2(n_5424),
.B1(n_5064),
.B2(n_5067),
.C1(n_5009),
.C2(n_5012),
.Y(n_6699)
);

OAI21x1_ASAP7_75t_L g6700 ( 
.A1(n_6430),
.A2(n_4844),
.B(n_5003),
.Y(n_6700)
);

INVx2_ASAP7_75t_L g6701 ( 
.A(n_5567),
.Y(n_6701)
);

OAI21x1_ASAP7_75t_L g6702 ( 
.A1(n_6430),
.A2(n_6329),
.B(n_6305),
.Y(n_6702)
);

A2O1A1Ixp33_ASAP7_75t_L g6703 ( 
.A1(n_6377),
.A2(n_5006),
.B(n_4870),
.C(n_4773),
.Y(n_6703)
);

CKINVDCx5p33_ASAP7_75t_R g6704 ( 
.A(n_5659),
.Y(n_6704)
);

OAI22xp5_ASAP7_75t_SL g6705 ( 
.A1(n_5760),
.A2(n_5414),
.B1(n_5173),
.B2(n_5336),
.Y(n_6705)
);

INVx1_ASAP7_75t_L g6706 ( 
.A(n_6248),
.Y(n_6706)
);

INVx1_ASAP7_75t_L g6707 ( 
.A(n_6249),
.Y(n_6707)
);

OAI22xp5_ASAP7_75t_L g6708 ( 
.A1(n_5570),
.A2(n_5501),
.B1(n_5353),
.B2(n_5188),
.Y(n_6708)
);

OR2x2_ASAP7_75t_L g6709 ( 
.A(n_5892),
.B(n_5421),
.Y(n_6709)
);

OAI21xp5_ASAP7_75t_L g6710 ( 
.A1(n_5732),
.A2(n_4934),
.B(n_4773),
.Y(n_6710)
);

NAND2x1p5_ASAP7_75t_L g6711 ( 
.A(n_5598),
.B(n_5114),
.Y(n_6711)
);

INVx1_ASAP7_75t_L g6712 ( 
.A(n_6249),
.Y(n_6712)
);

INVx2_ASAP7_75t_L g6713 ( 
.A(n_5567),
.Y(n_6713)
);

OAI21x1_ASAP7_75t_L g6714 ( 
.A1(n_6305),
.A2(n_5003),
.B(n_4769),
.Y(n_6714)
);

OAI221xp5_ASAP7_75t_L g6715 ( 
.A1(n_6221),
.A2(n_4951),
.B1(n_5366),
.B2(n_5012),
.C(n_5009),
.Y(n_6715)
);

OAI22xp33_ASAP7_75t_SL g6716 ( 
.A1(n_6221),
.A2(n_5067),
.B1(n_5064),
.B2(n_5051),
.Y(n_6716)
);

O2A1O1Ixp33_ASAP7_75t_L g6717 ( 
.A1(n_6415),
.A2(n_5403),
.B(n_5430),
.C(n_4934),
.Y(n_6717)
);

OAI21xp5_ASAP7_75t_L g6718 ( 
.A1(n_5732),
.A2(n_5430),
.B(n_4958),
.Y(n_6718)
);

OA21x2_ASAP7_75t_L g6719 ( 
.A1(n_5788),
.A2(n_4711),
.B(n_4696),
.Y(n_6719)
);

BUFx6f_ASAP7_75t_L g6720 ( 
.A(n_5598),
.Y(n_6720)
);

INVx2_ASAP7_75t_L g6721 ( 
.A(n_5590),
.Y(n_6721)
);

BUFx6f_ASAP7_75t_L g6722 ( 
.A(n_5598),
.Y(n_6722)
);

OAI21x1_ASAP7_75t_L g6723 ( 
.A1(n_6329),
.A2(n_5003),
.B(n_4769),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_6250),
.Y(n_6724)
);

INVx2_ASAP7_75t_SL g6725 ( 
.A(n_6246),
.Y(n_6725)
);

A2O1A1Ixp33_ASAP7_75t_L g6726 ( 
.A1(n_6377),
.A2(n_5542),
.B(n_5520),
.C(n_5476),
.Y(n_6726)
);

AOI22xp33_ASAP7_75t_L g6727 ( 
.A1(n_6216),
.A2(n_4912),
.B1(n_4939),
.B2(n_4959),
.Y(n_6727)
);

OA21x2_ASAP7_75t_L g6728 ( 
.A1(n_5788),
.A2(n_4696),
.B(n_5445),
.Y(n_6728)
);

INVx1_ASAP7_75t_SL g6729 ( 
.A(n_5756),
.Y(n_6729)
);

OAI21x1_ASAP7_75t_L g6730 ( 
.A1(n_6414),
.A2(n_5003),
.B(n_5049),
.Y(n_6730)
);

AOI221xp5_ASAP7_75t_L g6731 ( 
.A1(n_6042),
.A2(n_5500),
.B1(n_5529),
.B2(n_5497),
.C(n_5452),
.Y(n_6731)
);

INVx2_ASAP7_75t_L g6732 ( 
.A(n_5590),
.Y(n_6732)
);

INVx2_ASAP7_75t_L g6733 ( 
.A(n_5590),
.Y(n_6733)
);

INVx2_ASAP7_75t_L g6734 ( 
.A(n_5590),
.Y(n_6734)
);

INVx2_ASAP7_75t_SL g6735 ( 
.A(n_6246),
.Y(n_6735)
);

AOI22xp33_ASAP7_75t_L g6736 ( 
.A1(n_6216),
.A2(n_4912),
.B1(n_4939),
.B2(n_4959),
.Y(n_6736)
);

AND2x2_ASAP7_75t_L g6737 ( 
.A(n_5789),
.B(n_5523),
.Y(n_6737)
);

BUFx6f_ASAP7_75t_L g6738 ( 
.A(n_5598),
.Y(n_6738)
);

INVx1_ASAP7_75t_L g6739 ( 
.A(n_6250),
.Y(n_6739)
);

OR2x2_ASAP7_75t_L g6740 ( 
.A(n_5892),
.B(n_5304),
.Y(n_6740)
);

INVx2_ASAP7_75t_SL g6741 ( 
.A(n_6257),
.Y(n_6741)
);

OAI21xp5_ASAP7_75t_L g6742 ( 
.A1(n_5783),
.A2(n_4958),
.B(n_5403),
.Y(n_6742)
);

AO21x2_ASAP7_75t_L g6743 ( 
.A1(n_5920),
.A2(n_5030),
.B(n_5445),
.Y(n_6743)
);

AOI22xp5_ASAP7_75t_L g6744 ( 
.A1(n_5723),
.A2(n_5533),
.B1(n_4809),
.B2(n_4722),
.Y(n_6744)
);

AOI22xp33_ASAP7_75t_L g6745 ( 
.A1(n_5953),
.A2(n_4959),
.B1(n_5035),
.B2(n_4722),
.Y(n_6745)
);

AO222x2_ASAP7_75t_L g6746 ( 
.A1(n_6211),
.A2(n_5536),
.B1(n_5500),
.B2(n_5529),
.C1(n_5497),
.C2(n_5341),
.Y(n_6746)
);

NAND2x1p5_ASAP7_75t_L g6747 ( 
.A(n_5776),
.B(n_5114),
.Y(n_6747)
);

INVx2_ASAP7_75t_L g6748 ( 
.A(n_5594),
.Y(n_6748)
);

INVx2_ASAP7_75t_L g6749 ( 
.A(n_5594),
.Y(n_6749)
);

AND2x2_ASAP7_75t_L g6750 ( 
.A(n_5789),
.B(n_5523),
.Y(n_6750)
);

INVx2_ASAP7_75t_SL g6751 ( 
.A(n_6257),
.Y(n_6751)
);

O2A1O1Ixp33_ASAP7_75t_SL g6752 ( 
.A1(n_6222),
.A2(n_4792),
.B(n_4808),
.C(n_4744),
.Y(n_6752)
);

INVx1_ASAP7_75t_L g6753 ( 
.A(n_6262),
.Y(n_6753)
);

INVx2_ASAP7_75t_SL g6754 ( 
.A(n_6257),
.Y(n_6754)
);

OAI21x1_ASAP7_75t_L g6755 ( 
.A1(n_6414),
.A2(n_5049),
.B(n_4933),
.Y(n_6755)
);

AOI22xp33_ASAP7_75t_L g6756 ( 
.A1(n_5953),
.A2(n_4959),
.B1(n_4697),
.B2(n_4752),
.Y(n_6756)
);

AO31x2_ASAP7_75t_L g6757 ( 
.A1(n_5789),
.A2(n_4951),
.A3(n_5053),
.B(n_5051),
.Y(n_6757)
);

AOI22xp33_ASAP7_75t_L g6758 ( 
.A1(n_5947),
.A2(n_4959),
.B1(n_4697),
.B2(n_4752),
.Y(n_6758)
);

INVx3_ASAP7_75t_L g6759 ( 
.A(n_5641),
.Y(n_6759)
);

BUFx2_ASAP7_75t_SL g6760 ( 
.A(n_5629),
.Y(n_6760)
);

OAI21x1_ASAP7_75t_L g6761 ( 
.A1(n_6292),
.A2(n_5049),
.B(n_4933),
.Y(n_6761)
);

NAND2xp5_ASAP7_75t_L g6762 ( 
.A(n_5616),
.B(n_5313),
.Y(n_6762)
);

INVx1_ASAP7_75t_L g6763 ( 
.A(n_6262),
.Y(n_6763)
);

OAI21x1_ASAP7_75t_L g6764 ( 
.A1(n_5969),
.A2(n_5049),
.B(n_4904),
.Y(n_6764)
);

OAI21x1_ASAP7_75t_L g6765 ( 
.A1(n_5969),
.A2(n_4904),
.B(n_4949),
.Y(n_6765)
);

INVx1_ASAP7_75t_L g6766 ( 
.A(n_6271),
.Y(n_6766)
);

INVxp67_ASAP7_75t_L g6767 ( 
.A(n_6175),
.Y(n_6767)
);

NOR2xp67_ASAP7_75t_L g6768 ( 
.A(n_6257),
.B(n_4721),
.Y(n_6768)
);

A2O1A1Ixp33_ASAP7_75t_L g6769 ( 
.A1(n_6254),
.A2(n_5476),
.B(n_5533),
.C(n_4709),
.Y(n_6769)
);

OA21x2_ASAP7_75t_L g6770 ( 
.A1(n_5802),
.A2(n_5053),
.B(n_5169),
.Y(n_6770)
);

NAND2x1p5_ASAP7_75t_L g6771 ( 
.A(n_5776),
.B(n_5457),
.Y(n_6771)
);

NAND3xp33_ASAP7_75t_L g6772 ( 
.A(n_6374),
.B(n_5536),
.C(n_5062),
.Y(n_6772)
);

OR2x6_ASAP7_75t_L g6773 ( 
.A(n_6244),
.B(n_5081),
.Y(n_6773)
);

BUFx8_ASAP7_75t_L g6774 ( 
.A(n_6405),
.Y(n_6774)
);

INVx2_ASAP7_75t_L g6775 ( 
.A(n_5594),
.Y(n_6775)
);

O2A1O1Ixp33_ASAP7_75t_SL g6776 ( 
.A1(n_6222),
.A2(n_4744),
.B(n_4808),
.C(n_4792),
.Y(n_6776)
);

OAI21x1_ASAP7_75t_L g6777 ( 
.A1(n_5969),
.A2(n_4949),
.B(n_4762),
.Y(n_6777)
);

INVx2_ASAP7_75t_L g6778 ( 
.A(n_5594),
.Y(n_6778)
);

INVx1_ASAP7_75t_L g6779 ( 
.A(n_6271),
.Y(n_6779)
);

BUFx12f_ASAP7_75t_L g6780 ( 
.A(n_5914),
.Y(n_6780)
);

INVx2_ASAP7_75t_L g6781 ( 
.A(n_5601),
.Y(n_6781)
);

INVx1_ASAP7_75t_L g6782 ( 
.A(n_6272),
.Y(n_6782)
);

AND2x4_ASAP7_75t_L g6783 ( 
.A(n_5822),
.B(n_5526),
.Y(n_6783)
);

OAI21x1_ASAP7_75t_L g6784 ( 
.A1(n_6080),
.A2(n_4762),
.B(n_4677),
.Y(n_6784)
);

OAI21x1_ASAP7_75t_L g6785 ( 
.A1(n_6080),
.A2(n_4807),
.B(n_4677),
.Y(n_6785)
);

OAI21x1_ASAP7_75t_L g6786 ( 
.A1(n_6080),
.A2(n_4807),
.B(n_4677),
.Y(n_6786)
);

AOI222xp33_ASAP7_75t_L g6787 ( 
.A1(n_5947),
.A2(n_5424),
.B1(n_5331),
.B2(n_5341),
.C1(n_5347),
.C2(n_5346),
.Y(n_6787)
);

OAI21x1_ASAP7_75t_L g6788 ( 
.A1(n_6328),
.A2(n_4807),
.B(n_4677),
.Y(n_6788)
);

AOI22xp33_ASAP7_75t_L g6789 ( 
.A1(n_5974),
.A2(n_4959),
.B1(n_4701),
.B2(n_5362),
.Y(n_6789)
);

INVx1_ASAP7_75t_L g6790 ( 
.A(n_6272),
.Y(n_6790)
);

A2O1A1Ixp33_ASAP7_75t_L g6791 ( 
.A1(n_6254),
.A2(n_4709),
.B(n_4953),
.C(n_5400),
.Y(n_6791)
);

OAI21x1_ASAP7_75t_L g6792 ( 
.A1(n_6328),
.A2(n_6399),
.B(n_6053),
.Y(n_6792)
);

OAI21x1_ASAP7_75t_L g6793 ( 
.A1(n_6328),
.A2(n_4807),
.B(n_4677),
.Y(n_6793)
);

OA21x2_ASAP7_75t_L g6794 ( 
.A1(n_5802),
.A2(n_5186),
.B(n_5169),
.Y(n_6794)
);

OAI21x1_ASAP7_75t_L g6795 ( 
.A1(n_6399),
.A2(n_4807),
.B(n_5400),
.Y(n_6795)
);

AOI21xp5_ASAP7_75t_L g6796 ( 
.A1(n_5613),
.A2(n_6364),
.B(n_6053),
.Y(n_6796)
);

OR2x6_ASAP7_75t_L g6797 ( 
.A(n_6244),
.B(n_5266),
.Y(n_6797)
);

NAND2xp5_ASAP7_75t_L g6798 ( 
.A(n_5640),
.B(n_5329),
.Y(n_6798)
);

BUFx12f_ASAP7_75t_L g6799 ( 
.A(n_5845),
.Y(n_6799)
);

OAI21x1_ASAP7_75t_L g6800 ( 
.A1(n_6399),
.A2(n_5404),
.B(n_5491),
.Y(n_6800)
);

NOR2x1_ASAP7_75t_SL g6801 ( 
.A(n_6165),
.B(n_5463),
.Y(n_6801)
);

AOI22xp33_ASAP7_75t_L g6802 ( 
.A1(n_5974),
.A2(n_4959),
.B1(n_4701),
.B2(n_5362),
.Y(n_6802)
);

OAI21x1_ASAP7_75t_SL g6803 ( 
.A1(n_5543),
.A2(n_5464),
.B(n_5463),
.Y(n_6803)
);

INVx1_ASAP7_75t_L g6804 ( 
.A(n_6294),
.Y(n_6804)
);

OAI22xp5_ASAP7_75t_L g6805 ( 
.A1(n_5570),
.A2(n_5501),
.B1(n_4809),
.B2(n_5366),
.Y(n_6805)
);

AO31x2_ASAP7_75t_L g6806 ( 
.A1(n_5802),
.A2(n_5432),
.A3(n_4982),
.B(n_4978),
.Y(n_6806)
);

OAI21x1_ASAP7_75t_L g6807 ( 
.A1(n_6348),
.A2(n_5404),
.B(n_5491),
.Y(n_6807)
);

AOI21x1_ASAP7_75t_L g6808 ( 
.A1(n_5843),
.A2(n_6180),
.B(n_6175),
.Y(n_6808)
);

OAI21x1_ASAP7_75t_L g6809 ( 
.A1(n_6348),
.A2(n_5495),
.B(n_5492),
.Y(n_6809)
);

INVx1_ASAP7_75t_L g6810 ( 
.A(n_6294),
.Y(n_6810)
);

OAI21x1_ASAP7_75t_L g6811 ( 
.A1(n_6351),
.A2(n_5495),
.B(n_5492),
.Y(n_6811)
);

INVx3_ASAP7_75t_L g6812 ( 
.A(n_5641),
.Y(n_6812)
);

OA21x2_ASAP7_75t_L g6813 ( 
.A1(n_5815),
.A2(n_5265),
.B(n_5186),
.Y(n_6813)
);

BUFx6f_ASAP7_75t_L g6814 ( 
.A(n_5776),
.Y(n_6814)
);

AOI21xp5_ASAP7_75t_L g6815 ( 
.A1(n_5613),
.A2(n_5384),
.B(n_5538),
.Y(n_6815)
);

OAI21x1_ASAP7_75t_L g6816 ( 
.A1(n_6351),
.A2(n_5510),
.B(n_5507),
.Y(n_6816)
);

AND2x4_ASAP7_75t_L g6817 ( 
.A(n_5822),
.B(n_5526),
.Y(n_6817)
);

OAI21x1_ASAP7_75t_L g6818 ( 
.A1(n_6355),
.A2(n_5510),
.B(n_5507),
.Y(n_6818)
);

OAI21x1_ASAP7_75t_L g6819 ( 
.A1(n_6355),
.A2(n_4989),
.B(n_4825),
.Y(n_6819)
);

OAI21x1_ASAP7_75t_SL g6820 ( 
.A1(n_6129),
.A2(n_5464),
.B(n_5437),
.Y(n_6820)
);

INVx2_ASAP7_75t_L g6821 ( 
.A(n_5601),
.Y(n_6821)
);

AO21x2_ASAP7_75t_L g6822 ( 
.A1(n_5920),
.A2(n_4982),
.B(n_4978),
.Y(n_6822)
);

OAI21x1_ASAP7_75t_L g6823 ( 
.A1(n_6067),
.A2(n_4989),
.B(n_4825),
.Y(n_6823)
);

INVx8_ASAP7_75t_L g6824 ( 
.A(n_6405),
.Y(n_6824)
);

OA21x2_ASAP7_75t_L g6825 ( 
.A1(n_5815),
.A2(n_5837),
.B(n_5569),
.Y(n_6825)
);

HB1xp67_ASAP7_75t_L g6826 ( 
.A(n_5890),
.Y(n_6826)
);

OAI21x1_ASAP7_75t_L g6827 ( 
.A1(n_6067),
.A2(n_4989),
.B(n_4825),
.Y(n_6827)
);

HB1xp67_ASAP7_75t_L g6828 ( 
.A(n_5905),
.Y(n_6828)
);

HB1xp67_ASAP7_75t_L g6829 ( 
.A(n_5905),
.Y(n_6829)
);

A2O1A1Ixp33_ASAP7_75t_L g6830 ( 
.A1(n_5815),
.A2(n_4953),
.B(n_4903),
.C(n_5379),
.Y(n_6830)
);

AND2x4_ASAP7_75t_L g6831 ( 
.A(n_5822),
.B(n_4681),
.Y(n_6831)
);

INVx1_ASAP7_75t_L g6832 ( 
.A(n_6302),
.Y(n_6832)
);

NAND2xp5_ASAP7_75t_L g6833 ( 
.A(n_5640),
.B(n_5329),
.Y(n_6833)
);

OAI21x1_ASAP7_75t_L g6834 ( 
.A1(n_6071),
.A2(n_4989),
.B(n_4825),
.Y(n_6834)
);

INVx1_ASAP7_75t_L g6835 ( 
.A(n_6302),
.Y(n_6835)
);

CKINVDCx5p33_ASAP7_75t_R g6836 ( 
.A(n_5659),
.Y(n_6836)
);

O2A1O1Ixp33_ASAP7_75t_L g6837 ( 
.A1(n_6415),
.A2(n_5331),
.B(n_5347),
.C(n_5346),
.Y(n_6837)
);

OAI21x1_ASAP7_75t_L g6838 ( 
.A1(n_6071),
.A2(n_6379),
.B(n_6362),
.Y(n_6838)
);

AO21x2_ASAP7_75t_L g6839 ( 
.A1(n_6056),
.A2(n_5451),
.B(n_5024),
.Y(n_6839)
);

OAI22xp5_ASAP7_75t_L g6840 ( 
.A1(n_5645),
.A2(n_5351),
.B1(n_4827),
.B2(n_5437),
.Y(n_6840)
);

AND2x4_ASAP7_75t_L g6841 ( 
.A(n_5996),
.B(n_5997),
.Y(n_6841)
);

OAI21x1_ASAP7_75t_L g6842 ( 
.A1(n_6379),
.A2(n_5376),
.B(n_5251),
.Y(n_6842)
);

NOR2xp33_ASAP7_75t_SL g6843 ( 
.A(n_6398),
.B(n_5439),
.Y(n_6843)
);

NAND2x1p5_ASAP7_75t_L g6844 ( 
.A(n_5776),
.B(n_5457),
.Y(n_6844)
);

INVx1_ASAP7_75t_L g6845 ( 
.A(n_6304),
.Y(n_6845)
);

OA21x2_ASAP7_75t_L g6846 ( 
.A1(n_5837),
.A2(n_5569),
.B(n_5549),
.Y(n_6846)
);

BUFx10_ASAP7_75t_L g6847 ( 
.A(n_6018),
.Y(n_6847)
);

INVx1_ASAP7_75t_L g6848 ( 
.A(n_6304),
.Y(n_6848)
);

OAI21x1_ASAP7_75t_L g6849 ( 
.A1(n_6362),
.A2(n_5376),
.B(n_5251),
.Y(n_6849)
);

AND2x4_ASAP7_75t_L g6850 ( 
.A(n_5996),
.B(n_4681),
.Y(n_6850)
);

CKINVDCx20_ASAP7_75t_R g6851 ( 
.A(n_5583),
.Y(n_6851)
);

AO31x2_ASAP7_75t_L g6852 ( 
.A1(n_5837),
.A2(n_5432),
.A3(n_5198),
.B(n_5201),
.Y(n_6852)
);

OAI21x1_ASAP7_75t_L g6853 ( 
.A1(n_5684),
.A2(n_5376),
.B(n_5251),
.Y(n_6853)
);

BUFx3_ASAP7_75t_L g6854 ( 
.A(n_5942),
.Y(n_6854)
);

OA21x2_ASAP7_75t_L g6855 ( 
.A1(n_5549),
.A2(n_5265),
.B(n_5538),
.Y(n_6855)
);

INVx2_ASAP7_75t_L g6856 ( 
.A(n_5601),
.Y(n_6856)
);

OAI21xp5_ASAP7_75t_L g6857 ( 
.A1(n_5783),
.A2(n_4907),
.B(n_4705),
.Y(n_6857)
);

AOI22xp33_ASAP7_75t_L g6858 ( 
.A1(n_5961),
.A2(n_4959),
.B1(n_5477),
.B2(n_4776),
.Y(n_6858)
);

OAI22xp5_ASAP7_75t_L g6859 ( 
.A1(n_5645),
.A2(n_5351),
.B1(n_4827),
.B2(n_5379),
.Y(n_6859)
);

NAND2x1p5_ASAP7_75t_L g6860 ( 
.A(n_5776),
.B(n_5457),
.Y(n_6860)
);

INVxp67_ASAP7_75t_SL g6861 ( 
.A(n_5959),
.Y(n_6861)
);

AO21x2_ASAP7_75t_L g6862 ( 
.A1(n_6056),
.A2(n_6374),
.B(n_6439),
.Y(n_6862)
);

AOI22xp33_ASAP7_75t_L g6863 ( 
.A1(n_5961),
.A2(n_5477),
.B1(n_4776),
.B2(n_5384),
.Y(n_6863)
);

INVx2_ASAP7_75t_L g6864 ( 
.A(n_5601),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_6309),
.Y(n_6865)
);

AOI22xp33_ASAP7_75t_L g6866 ( 
.A1(n_5976),
.A2(n_4855),
.B1(n_4851),
.B2(n_4789),
.Y(n_6866)
);

AND2x4_ASAP7_75t_L g6867 ( 
.A(n_5996),
.B(n_4698),
.Y(n_6867)
);

INVx1_ASAP7_75t_L g6868 ( 
.A(n_6309),
.Y(n_6868)
);

OAI21x1_ASAP7_75t_L g6869 ( 
.A1(n_5684),
.A2(n_5376),
.B(n_5251),
.Y(n_6869)
);

OR2x2_ASAP7_75t_L g6870 ( 
.A(n_5941),
.B(n_5304),
.Y(n_6870)
);

INVx2_ASAP7_75t_SL g6871 ( 
.A(n_6257),
.Y(n_6871)
);

OAI21x1_ASAP7_75t_L g6872 ( 
.A1(n_5835),
.A2(n_4856),
.B(n_4705),
.Y(n_6872)
);

OAI21x1_ASAP7_75t_L g6873 ( 
.A1(n_5835),
.A2(n_4856),
.B(n_4676),
.Y(n_6873)
);

NOR2xp33_ASAP7_75t_L g6874 ( 
.A(n_5977),
.B(n_5391),
.Y(n_6874)
);

NAND2xp5_ASAP7_75t_L g6875 ( 
.A(n_5643),
.B(n_5435),
.Y(n_6875)
);

OAI21x1_ASAP7_75t_SL g6876 ( 
.A1(n_6129),
.A2(n_5518),
.B(n_5502),
.Y(n_6876)
);

OAI22xp33_ASAP7_75t_L g6877 ( 
.A1(n_5964),
.A2(n_6161),
.B1(n_5804),
.B2(n_5695),
.Y(n_6877)
);

NOR2xp33_ASAP7_75t_L g6878 ( 
.A(n_5979),
.B(n_5391),
.Y(n_6878)
);

CKINVDCx20_ASAP7_75t_R g6879 ( 
.A(n_5583),
.Y(n_6879)
);

INVx1_ASAP7_75t_L g6880 ( 
.A(n_6322),
.Y(n_6880)
);

OA21x2_ASAP7_75t_L g6881 ( 
.A1(n_5569),
.A2(n_5024),
.B(n_5451),
.Y(n_6881)
);

AOI21xp5_ASAP7_75t_L g6882 ( 
.A1(n_6364),
.A2(n_4903),
.B(n_4907),
.Y(n_6882)
);

CKINVDCx5p33_ASAP7_75t_R g6883 ( 
.A(n_5746),
.Y(n_6883)
);

AOI22xp5_ASAP7_75t_L g6884 ( 
.A1(n_6161),
.A2(n_5964),
.B1(n_5990),
.B2(n_5976),
.Y(n_6884)
);

INVx6_ASAP7_75t_L g6885 ( 
.A(n_6257),
.Y(n_6885)
);

INVx1_ASAP7_75t_L g6886 ( 
.A(n_6322),
.Y(n_6886)
);

BUFx12f_ASAP7_75t_L g6887 ( 
.A(n_5845),
.Y(n_6887)
);

NAND2x1p5_ASAP7_75t_L g6888 ( 
.A(n_5776),
.B(n_5457),
.Y(n_6888)
);

INVx2_ASAP7_75t_L g6889 ( 
.A(n_5605),
.Y(n_6889)
);

NAND2xp5_ASAP7_75t_L g6890 ( 
.A(n_5643),
.B(n_5984),
.Y(n_6890)
);

BUFx12f_ASAP7_75t_L g6891 ( 
.A(n_5611),
.Y(n_6891)
);

AND2x2_ASAP7_75t_L g6892 ( 
.A(n_6368),
.B(n_5523),
.Y(n_6892)
);

OAI21x1_ASAP7_75t_L g6893 ( 
.A1(n_5835),
.A2(n_4676),
.B(n_5218),
.Y(n_6893)
);

AO21x2_ASAP7_75t_L g6894 ( 
.A1(n_6056),
.A2(n_4997),
.B(n_4995),
.Y(n_6894)
);

OA21x2_ASAP7_75t_L g6895 ( 
.A1(n_5612),
.A2(n_5024),
.B(n_5435),
.Y(n_6895)
);

AOI22xp33_ASAP7_75t_L g6896 ( 
.A1(n_6295),
.A2(n_4855),
.B1(n_4851),
.B2(n_4789),
.Y(n_6896)
);

AO21x2_ASAP7_75t_L g6897 ( 
.A1(n_6056),
.A2(n_5024),
.B(n_4997),
.Y(n_6897)
);

OAI21x1_ASAP7_75t_L g6898 ( 
.A1(n_5835),
.A2(n_5228),
.B(n_5218),
.Y(n_6898)
);

AOI21x1_ASAP7_75t_L g6899 ( 
.A1(n_5843),
.A2(n_5439),
.B(n_5144),
.Y(n_6899)
);

INVx1_ASAP7_75t_L g6900 ( 
.A(n_6331),
.Y(n_6900)
);

OAI21x1_ASAP7_75t_L g6901 ( 
.A1(n_6101),
.A2(n_5228),
.B(n_5218),
.Y(n_6901)
);

HB1xp67_ASAP7_75t_L g6902 ( 
.A(n_5939),
.Y(n_6902)
);

OAI21x1_ASAP7_75t_L g6903 ( 
.A1(n_6101),
.A2(n_5228),
.B(n_5218),
.Y(n_6903)
);

INVx3_ASAP7_75t_L g6904 ( 
.A(n_5641),
.Y(n_6904)
);

INVx1_ASAP7_75t_L g6905 ( 
.A(n_6331),
.Y(n_6905)
);

INVx3_ASAP7_75t_L g6906 ( 
.A(n_5642),
.Y(n_6906)
);

AND2x2_ASAP7_75t_L g6907 ( 
.A(n_6368),
.B(n_5530),
.Y(n_6907)
);

INVx2_ASAP7_75t_L g6908 ( 
.A(n_5605),
.Y(n_6908)
);

AOI22xp33_ASAP7_75t_L g6909 ( 
.A1(n_6295),
.A2(n_5651),
.B1(n_6389),
.B2(n_5791),
.Y(n_6909)
);

INVx2_ASAP7_75t_L g6910 ( 
.A(n_5605),
.Y(n_6910)
);

NAND2xp5_ASAP7_75t_L g6911 ( 
.A(n_5984),
.B(n_5372),
.Y(n_6911)
);

NAND2xp5_ASAP7_75t_L g6912 ( 
.A(n_5986),
.B(n_5372),
.Y(n_6912)
);

INVx6_ASAP7_75t_L g6913 ( 
.A(n_6257),
.Y(n_6913)
);

AND2x2_ASAP7_75t_L g6914 ( 
.A(n_6368),
.B(n_5530),
.Y(n_6914)
);

OAI22xp33_ASAP7_75t_SL g6915 ( 
.A1(n_6195),
.A2(n_5010),
.B1(n_5415),
.B2(n_5412),
.Y(n_6915)
);

OAI21x1_ASAP7_75t_SL g6916 ( 
.A1(n_5592),
.A2(n_5518),
.B(n_5502),
.Y(n_6916)
);

AOI22xp33_ASAP7_75t_SL g6917 ( 
.A1(n_5599),
.A2(n_5316),
.B1(n_5410),
.B2(n_5024),
.Y(n_6917)
);

NOR2xp33_ASAP7_75t_L g6918 ( 
.A(n_5979),
.B(n_5394),
.Y(n_6918)
);

BUFx6f_ASAP7_75t_L g6919 ( 
.A(n_5776),
.Y(n_6919)
);

OAI21x1_ASAP7_75t_L g6920 ( 
.A1(n_6101),
.A2(n_5228),
.B(n_5218),
.Y(n_6920)
);

CKINVDCx5p33_ASAP7_75t_R g6921 ( 
.A(n_5746),
.Y(n_6921)
);

OAI21x1_ASAP7_75t_L g6922 ( 
.A1(n_6101),
.A2(n_5230),
.B(n_5228),
.Y(n_6922)
);

OAI21x1_ASAP7_75t_L g6923 ( 
.A1(n_5578),
.A2(n_5239),
.B(n_5230),
.Y(n_6923)
);

OAI21x1_ASAP7_75t_L g6924 ( 
.A1(n_5578),
.A2(n_5239),
.B(n_5230),
.Y(n_6924)
);

AND2x2_ASAP7_75t_L g6925 ( 
.A(n_5612),
.B(n_5530),
.Y(n_6925)
);

CKINVDCx5p33_ASAP7_75t_R g6926 ( 
.A(n_5831),
.Y(n_6926)
);

A2O1A1Ixp33_ASAP7_75t_L g6927 ( 
.A1(n_6028),
.A2(n_5386),
.B(n_5010),
.C(n_5039),
.Y(n_6927)
);

AOI21x1_ASAP7_75t_L g6928 ( 
.A1(n_6180),
.A2(n_5144),
.B(n_5128),
.Y(n_6928)
);

AND2x4_ASAP7_75t_L g6929 ( 
.A(n_5996),
.B(n_5997),
.Y(n_6929)
);

INVx4_ASAP7_75t_SL g6930 ( 
.A(n_5573),
.Y(n_6930)
);

INVx4_ASAP7_75t_L g6931 ( 
.A(n_5698),
.Y(n_6931)
);

OAI21x1_ASAP7_75t_L g6932 ( 
.A1(n_5581),
.A2(n_5239),
.B(n_5230),
.Y(n_6932)
);

OA21x2_ASAP7_75t_L g6933 ( 
.A1(n_5612),
.A2(n_5637),
.B(n_5623),
.Y(n_6933)
);

INVx1_ASAP7_75t_L g6934 ( 
.A(n_6336),
.Y(n_6934)
);

NAND2xp5_ASAP7_75t_L g6935 ( 
.A(n_5986),
.B(n_4972),
.Y(n_6935)
);

OA21x2_ASAP7_75t_L g6936 ( 
.A1(n_5623),
.A2(n_5144),
.B(n_5128),
.Y(n_6936)
);

AOI22xp33_ASAP7_75t_L g6937 ( 
.A1(n_6295),
.A2(n_4855),
.B1(n_4851),
.B2(n_4789),
.Y(n_6937)
);

OR2x2_ASAP7_75t_L g6938 ( 
.A(n_5941),
.B(n_5062),
.Y(n_6938)
);

OAI21x1_ASAP7_75t_L g6939 ( 
.A1(n_5581),
.A2(n_5239),
.B(n_5230),
.Y(n_6939)
);

NAND2xp5_ASAP7_75t_L g6940 ( 
.A(n_6015),
.B(n_5082),
.Y(n_6940)
);

NAND2x1p5_ASAP7_75t_L g6941 ( 
.A(n_5776),
.B(n_5457),
.Y(n_6941)
);

CKINVDCx20_ASAP7_75t_R g6942 ( 
.A(n_5867),
.Y(n_6942)
);

OR2x6_ASAP7_75t_L g6943 ( 
.A(n_6244),
.B(n_5266),
.Y(n_6943)
);

AO31x2_ASAP7_75t_L g6944 ( 
.A1(n_5738),
.A2(n_5198),
.A3(n_5201),
.B(n_5195),
.Y(n_6944)
);

AOI221xp5_ASAP7_75t_SL g6945 ( 
.A1(n_5739),
.A2(n_5386),
.B1(n_5405),
.B2(n_5394),
.C(n_5412),
.Y(n_6945)
);

NAND2xp5_ASAP7_75t_L g6946 ( 
.A(n_6015),
.B(n_5082),
.Y(n_6946)
);

AND2x2_ASAP7_75t_L g6947 ( 
.A(n_5623),
.B(n_5637),
.Y(n_6947)
);

AOI22xp33_ASAP7_75t_L g6948 ( 
.A1(n_6295),
.A2(n_4855),
.B1(n_4851),
.B2(n_4789),
.Y(n_6948)
);

A2O1A1Ixp33_ASAP7_75t_L g6949 ( 
.A1(n_6028),
.A2(n_5010),
.B(n_5039),
.C(n_5038),
.Y(n_6949)
);

AND2x4_ASAP7_75t_L g6950 ( 
.A(n_5997),
.B(n_4698),
.Y(n_6950)
);

INVx4_ASAP7_75t_SL g6951 ( 
.A(n_5573),
.Y(n_6951)
);

INVx2_ASAP7_75t_L g6952 ( 
.A(n_5605),
.Y(n_6952)
);

AND2x2_ASAP7_75t_L g6953 ( 
.A(n_5637),
.B(n_5427),
.Y(n_6953)
);

CKINVDCx16_ASAP7_75t_R g6954 ( 
.A(n_6398),
.Y(n_6954)
);

BUFx2_ASAP7_75t_SL g6955 ( 
.A(n_5629),
.Y(n_6955)
);

AO21x1_ASAP7_75t_L g6956 ( 
.A1(n_5941),
.A2(n_5537),
.B(n_5471),
.Y(n_6956)
);

AND2x2_ASAP7_75t_L g6957 ( 
.A(n_5646),
.B(n_5427),
.Y(n_6957)
);

INVx1_ASAP7_75t_L g6958 ( 
.A(n_6336),
.Y(n_6958)
);

OA21x2_ASAP7_75t_L g6959 ( 
.A1(n_5646),
.A2(n_5145),
.B(n_5128),
.Y(n_6959)
);

AOI22xp5_ASAP7_75t_L g6960 ( 
.A1(n_5990),
.A2(n_5381),
.B1(n_5406),
.B2(n_5385),
.Y(n_6960)
);

INVx2_ASAP7_75t_L g6961 ( 
.A(n_5607),
.Y(n_6961)
);

CKINVDCx6p67_ASAP7_75t_R g6962 ( 
.A(n_5823),
.Y(n_6962)
);

OAI22xp5_ASAP7_75t_L g6963 ( 
.A1(n_5600),
.A2(n_5405),
.B1(n_5433),
.B2(n_5415),
.Y(n_6963)
);

AND2x2_ASAP7_75t_L g6964 ( 
.A(n_5646),
.B(n_5427),
.Y(n_6964)
);

INVx3_ASAP7_75t_L g6965 ( 
.A(n_5642),
.Y(n_6965)
);

AND2x4_ASAP7_75t_L g6966 ( 
.A(n_5997),
.B(n_4698),
.Y(n_6966)
);

BUFx12f_ASAP7_75t_L g6967 ( 
.A(n_5611),
.Y(n_6967)
);

BUFx2_ASAP7_75t_L g6968 ( 
.A(n_5663),
.Y(n_6968)
);

INVx2_ASAP7_75t_L g6969 ( 
.A(n_5607),
.Y(n_6969)
);

INVx1_ASAP7_75t_L g6970 ( 
.A(n_6337),
.Y(n_6970)
);

NOR3xp33_ASAP7_75t_SL g6971 ( 
.A(n_5615),
.B(n_4917),
.C(n_4894),
.Y(n_6971)
);

A2O1A1Ixp33_ASAP7_75t_L g6972 ( 
.A1(n_6145),
.A2(n_5039),
.B(n_5038),
.C(n_5381),
.Y(n_6972)
);

INVx1_ASAP7_75t_L g6973 ( 
.A(n_6337),
.Y(n_6973)
);

NOR2xp33_ASAP7_75t_L g6974 ( 
.A(n_5830),
.B(n_5433),
.Y(n_6974)
);

INVx2_ASAP7_75t_L g6975 ( 
.A(n_5607),
.Y(n_6975)
);

AND2x2_ASAP7_75t_L g6976 ( 
.A(n_5663),
.B(n_5429),
.Y(n_6976)
);

BUFx2_ASAP7_75t_L g6977 ( 
.A(n_5663),
.Y(n_6977)
);

OAI22xp33_ASAP7_75t_L g6978 ( 
.A1(n_5804),
.A2(n_5406),
.B1(n_5385),
.B2(n_5531),
.Y(n_6978)
);

AOI21xp5_ASAP7_75t_L g6979 ( 
.A1(n_5648),
.A2(n_5147),
.B(n_5145),
.Y(n_6979)
);

INVx3_ASAP7_75t_L g6980 ( 
.A(n_5642),
.Y(n_6980)
);

NAND2xp5_ASAP7_75t_L g6981 ( 
.A(n_5544),
.B(n_5146),
.Y(n_6981)
);

INVx2_ASAP7_75t_L g6982 ( 
.A(n_5607),
.Y(n_6982)
);

OAI21x1_ASAP7_75t_L g6983 ( 
.A1(n_5839),
.A2(n_5276),
.B(n_5245),
.Y(n_6983)
);

BUFx10_ASAP7_75t_L g6984 ( 
.A(n_6018),
.Y(n_6984)
);

INVx1_ASAP7_75t_L g6985 ( 
.A(n_6338),
.Y(n_6985)
);

OAI21x1_ASAP7_75t_L g6986 ( 
.A1(n_5839),
.A2(n_5649),
.B(n_5711),
.Y(n_6986)
);

INVx1_ASAP7_75t_L g6987 ( 
.A(n_6338),
.Y(n_6987)
);

OA21x2_ASAP7_75t_L g6988 ( 
.A1(n_5692),
.A2(n_5147),
.B(n_5145),
.Y(n_6988)
);

INVx1_ASAP7_75t_L g6989 ( 
.A(n_6344),
.Y(n_6989)
);

INVx2_ASAP7_75t_L g6990 ( 
.A(n_5618),
.Y(n_6990)
);

CKINVDCx20_ASAP7_75t_R g6991 ( 
.A(n_6020),
.Y(n_6991)
);

AO31x2_ASAP7_75t_L g6992 ( 
.A1(n_5738),
.A2(n_5202),
.A3(n_5205),
.B(n_5195),
.Y(n_6992)
);

AND2x6_ASAP7_75t_L g6993 ( 
.A(n_5554),
.B(n_4541),
.Y(n_6993)
);

INVx2_ASAP7_75t_L g6994 ( 
.A(n_5618),
.Y(n_6994)
);

OAI21x1_ASAP7_75t_SL g6995 ( 
.A1(n_5592),
.A2(n_5518),
.B(n_5471),
.Y(n_6995)
);

OAI21x1_ASAP7_75t_L g6996 ( 
.A1(n_5649),
.A2(n_5307),
.B(n_5276),
.Y(n_6996)
);

OAI21x1_ASAP7_75t_L g6997 ( 
.A1(n_5711),
.A2(n_5312),
.B(n_5307),
.Y(n_6997)
);

INVx1_ASAP7_75t_L g6998 ( 
.A(n_6344),
.Y(n_6998)
);

INVx1_ASAP7_75t_L g6999 ( 
.A(n_6359),
.Y(n_6999)
);

BUFx3_ASAP7_75t_L g7000 ( 
.A(n_5991),
.Y(n_7000)
);

OAI21xp5_ASAP7_75t_L g7001 ( 
.A1(n_5651),
.A2(n_5146),
.B(n_5335),
.Y(n_7001)
);

OAI22xp5_ASAP7_75t_L g7002 ( 
.A1(n_5600),
.A2(n_5444),
.B1(n_5443),
.B2(n_5429),
.Y(n_7002)
);

OAI21x1_ASAP7_75t_L g7003 ( 
.A1(n_6437),
.A2(n_5686),
.B(n_5683),
.Y(n_7003)
);

BUFx8_ASAP7_75t_L g7004 ( 
.A(n_6405),
.Y(n_7004)
);

NAND3xp33_ASAP7_75t_L g7005 ( 
.A(n_5725),
.B(n_4877),
.C(n_4848),
.Y(n_7005)
);

O2A1O1Ixp33_ASAP7_75t_L g7006 ( 
.A1(n_6415),
.A2(n_5335),
.B(n_4877),
.C(n_4886),
.Y(n_7006)
);

OAI221xp5_ASAP7_75t_L g7007 ( 
.A1(n_6389),
.A2(n_5453),
.B1(n_5440),
.B2(n_5444),
.C(n_5443),
.Y(n_7007)
);

INVx5_ASAP7_75t_L g7008 ( 
.A(n_6295),
.Y(n_7008)
);

INVx1_ASAP7_75t_L g7009 ( 
.A(n_6359),
.Y(n_7009)
);

OAI22xp5_ASAP7_75t_L g7010 ( 
.A1(n_5725),
.A2(n_5429),
.B1(n_5470),
.B2(n_5468),
.Y(n_7010)
);

INVx1_ASAP7_75t_L g7011 ( 
.A(n_6363),
.Y(n_7011)
);

INVx2_ASAP7_75t_SL g7012 ( 
.A(n_6257),
.Y(n_7012)
);

NOR2xp33_ASAP7_75t_L g7013 ( 
.A(n_5830),
.B(n_5527),
.Y(n_7013)
);

OAI22xp33_ASAP7_75t_SL g7014 ( 
.A1(n_6195),
.A2(n_5484),
.B1(n_5266),
.B2(n_5458),
.Y(n_7014)
);

NAND2xp5_ASAP7_75t_L g7015 ( 
.A(n_5544),
.B(n_5557),
.Y(n_7015)
);

NOR2xp67_ASAP7_75t_L g7016 ( 
.A(n_6361),
.B(n_6394),
.Y(n_7016)
);

CKINVDCx16_ASAP7_75t_R g7017 ( 
.A(n_6020),
.Y(n_7017)
);

AO21x2_ASAP7_75t_L g7018 ( 
.A1(n_6439),
.A2(n_4997),
.B(n_4995),
.Y(n_7018)
);

NOR2xp33_ASAP7_75t_L g7019 ( 
.A(n_5836),
.B(n_5527),
.Y(n_7019)
);

OA21x2_ASAP7_75t_L g7020 ( 
.A1(n_5692),
.A2(n_5148),
.B(n_5147),
.Y(n_7020)
);

OAI22xp5_ASAP7_75t_L g7021 ( 
.A1(n_5735),
.A2(n_5468),
.B1(n_5487),
.B2(n_5470),
.Y(n_7021)
);

OA21x2_ASAP7_75t_L g7022 ( 
.A1(n_5692),
.A2(n_5742),
.B(n_6394),
.Y(n_7022)
);

NOR2xp67_ASAP7_75t_L g7023 ( 
.A(n_6361),
.B(n_4721),
.Y(n_7023)
);

OAI22xp33_ASAP7_75t_L g7024 ( 
.A1(n_5695),
.A2(n_5531),
.B1(n_5525),
.B2(n_4789),
.Y(n_7024)
);

NOR2xp33_ASAP7_75t_SL g7025 ( 
.A(n_5671),
.B(n_5360),
.Y(n_7025)
);

INVxp67_ASAP7_75t_L g7026 ( 
.A(n_5557),
.Y(n_7026)
);

INVx1_ASAP7_75t_L g7027 ( 
.A(n_6363),
.Y(n_7027)
);

CKINVDCx5p33_ASAP7_75t_R g7028 ( 
.A(n_5831),
.Y(n_7028)
);

AOI22xp5_ASAP7_75t_L g7029 ( 
.A1(n_5671),
.A2(n_4702),
.B1(n_4725),
.B2(n_4720),
.Y(n_7029)
);

A2O1A1Ixp33_ASAP7_75t_L g7030 ( 
.A1(n_6145),
.A2(n_5039),
.B(n_5038),
.C(n_4717),
.Y(n_7030)
);

OAI21xp5_ASAP7_75t_L g7031 ( 
.A1(n_6017),
.A2(n_4886),
.B(n_4848),
.Y(n_7031)
);

AND2x4_ASAP7_75t_L g7032 ( 
.A(n_6037),
.B(n_4698),
.Y(n_7032)
);

OA21x2_ASAP7_75t_L g7033 ( 
.A1(n_5742),
.A2(n_5177),
.B(n_5148),
.Y(n_7033)
);

INVx2_ASAP7_75t_SL g7034 ( 
.A(n_6361),
.Y(n_7034)
);

INVx1_ASAP7_75t_L g7035 ( 
.A(n_6376),
.Y(n_7035)
);

OAI21xp5_ASAP7_75t_L g7036 ( 
.A1(n_6017),
.A2(n_4892),
.B(n_4888),
.Y(n_7036)
);

OA21x2_ASAP7_75t_L g7037 ( 
.A1(n_6176),
.A2(n_5768),
.B(n_6178),
.Y(n_7037)
);

BUFx6f_ASAP7_75t_L g7038 ( 
.A(n_5776),
.Y(n_7038)
);

A2O1A1Ixp33_ASAP7_75t_L g7039 ( 
.A1(n_6176),
.A2(n_5039),
.B(n_5038),
.C(n_4717),
.Y(n_7039)
);

INVx2_ASAP7_75t_L g7040 ( 
.A(n_5618),
.Y(n_7040)
);

OR2x2_ASAP7_75t_L g7041 ( 
.A(n_5689),
.B(n_5453),
.Y(n_7041)
);

BUFx3_ASAP7_75t_L g7042 ( 
.A(n_5991),
.Y(n_7042)
);

INVx1_ASAP7_75t_L g7043 ( 
.A(n_6376),
.Y(n_7043)
);

AOI221xp5_ASAP7_75t_L g7044 ( 
.A1(n_5948),
.A2(n_5458),
.B1(n_5454),
.B2(n_5537),
.C(n_4725),
.Y(n_7044)
);

NAND2x1p5_ASAP7_75t_L g7045 ( 
.A(n_5878),
.B(n_4721),
.Y(n_7045)
);

NAND2x1_ASAP7_75t_L g7046 ( 
.A(n_6104),
.B(n_5148),
.Y(n_7046)
);

AND2x4_ASAP7_75t_L g7047 ( 
.A(n_6037),
.B(n_4698),
.Y(n_7047)
);

INVx2_ASAP7_75t_L g7048 ( 
.A(n_5618),
.Y(n_7048)
);

OA21x2_ASAP7_75t_L g7049 ( 
.A1(n_5768),
.A2(n_5209),
.B(n_5177),
.Y(n_7049)
);

AND2x4_ASAP7_75t_L g7050 ( 
.A(n_6037),
.B(n_4704),
.Y(n_7050)
);

INVxp67_ASAP7_75t_L g7051 ( 
.A(n_6044),
.Y(n_7051)
);

BUFx6f_ASAP7_75t_L g7052 ( 
.A(n_5878),
.Y(n_7052)
);

OAI21xp5_ASAP7_75t_L g7053 ( 
.A1(n_6081),
.A2(n_4892),
.B(n_4888),
.Y(n_7053)
);

OR2x2_ASAP7_75t_L g7054 ( 
.A(n_5689),
.B(n_5454),
.Y(n_7054)
);

OR2x6_ASAP7_75t_L g7055 ( 
.A(n_6244),
.B(n_5266),
.Y(n_7055)
);

AOI22xp33_ASAP7_75t_L g7056 ( 
.A1(n_6295),
.A2(n_4855),
.B1(n_4851),
.B2(n_4789),
.Y(n_7056)
);

INVx4_ASAP7_75t_L g7057 ( 
.A(n_5991),
.Y(n_7057)
);

INVx1_ASAP7_75t_L g7058 ( 
.A(n_6378),
.Y(n_7058)
);

AO21x2_ASAP7_75t_L g7059 ( 
.A1(n_5556),
.A2(n_4999),
.B(n_4995),
.Y(n_7059)
);

AOI221xp5_ASAP7_75t_L g7060 ( 
.A1(n_5948),
.A2(n_4725),
.B1(n_4756),
.B2(n_4720),
.C(n_4702),
.Y(n_7060)
);

INVx5_ASAP7_75t_L g7061 ( 
.A(n_6295),
.Y(n_7061)
);

NOR2x1_ASAP7_75t_SL g7062 ( 
.A(n_6165),
.B(n_5489),
.Y(n_7062)
);

AOI21xp33_ASAP7_75t_SL g7063 ( 
.A1(n_5615),
.A2(n_5171),
.B(n_5005),
.Y(n_7063)
);

NAND2x1p5_ASAP7_75t_L g7064 ( 
.A(n_5878),
.B(n_4721),
.Y(n_7064)
);

AO21x2_ASAP7_75t_L g7065 ( 
.A1(n_5556),
.A2(n_5002),
.B(n_4999),
.Y(n_7065)
);

AND2x2_ASAP7_75t_L g7066 ( 
.A(n_6327),
.B(n_5468),
.Y(n_7066)
);

AOI221xp5_ASAP7_75t_L g7067 ( 
.A1(n_6044),
.A2(n_4756),
.B1(n_4767),
.B2(n_4720),
.C(n_4702),
.Y(n_7067)
);

INVx2_ASAP7_75t_SL g7068 ( 
.A(n_6361),
.Y(n_7068)
);

NAND2xp5_ASAP7_75t_L g7069 ( 
.A(n_5690),
.B(n_4798),
.Y(n_7069)
);

INVx1_ASAP7_75t_L g7070 ( 
.A(n_6378),
.Y(n_7070)
);

INVx1_ASAP7_75t_L g7071 ( 
.A(n_6380),
.Y(n_7071)
);

OR2x2_ASAP7_75t_L g7072 ( 
.A(n_5690),
.B(n_5177),
.Y(n_7072)
);

OAI21x1_ASAP7_75t_SL g7073 ( 
.A1(n_5592),
.A2(n_5363),
.B(n_5360),
.Y(n_7073)
);

INVx2_ASAP7_75t_L g7074 ( 
.A(n_5652),
.Y(n_7074)
);

O2A1O1Ixp33_ASAP7_75t_SL g7075 ( 
.A1(n_5566),
.A2(n_5466),
.B(n_5369),
.C(n_5535),
.Y(n_7075)
);

AOI221xp5_ASAP7_75t_L g7076 ( 
.A1(n_6031),
.A2(n_4786),
.B1(n_4767),
.B2(n_4756),
.C(n_5202),
.Y(n_7076)
);

NOR2xp33_ASAP7_75t_L g7077 ( 
.A(n_5836),
.B(n_6031),
.Y(n_7077)
);

INVx1_ASAP7_75t_L g7078 ( 
.A(n_6380),
.Y(n_7078)
);

OAI22xp5_ASAP7_75t_L g7079 ( 
.A1(n_5735),
.A2(n_5470),
.B1(n_5504),
.B2(n_5487),
.Y(n_7079)
);

AO21x2_ASAP7_75t_L g7080 ( 
.A1(n_5556),
.A2(n_5002),
.B(n_4999),
.Y(n_7080)
);

INVx2_ASAP7_75t_L g7081 ( 
.A(n_5652),
.Y(n_7081)
);

OAI21xp5_ASAP7_75t_L g7082 ( 
.A1(n_5710),
.A2(n_4795),
.B(n_4777),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_6383),
.Y(n_7083)
);

INVx3_ASAP7_75t_L g7084 ( 
.A(n_5642),
.Y(n_7084)
);

HB1xp67_ASAP7_75t_L g7085 ( 
.A(n_5939),
.Y(n_7085)
);

NAND2xp5_ASAP7_75t_L g7086 ( 
.A(n_6105),
.B(n_4798),
.Y(n_7086)
);

INVx1_ASAP7_75t_L g7087 ( 
.A(n_6383),
.Y(n_7087)
);

AOI22xp33_ASAP7_75t_L g7088 ( 
.A1(n_6295),
.A2(n_4855),
.B1(n_4851),
.B2(n_4775),
.Y(n_7088)
);

INVx1_ASAP7_75t_L g7089 ( 
.A(n_6396),
.Y(n_7089)
);

INVx2_ASAP7_75t_L g7090 ( 
.A(n_5652),
.Y(n_7090)
);

BUFx2_ASAP7_75t_L g7091 ( 
.A(n_6195),
.Y(n_7091)
);

INVx1_ASAP7_75t_L g7092 ( 
.A(n_6396),
.Y(n_7092)
);

AO21x2_ASAP7_75t_L g7093 ( 
.A1(n_5556),
.A2(n_5011),
.B(n_5002),
.Y(n_7093)
);

AND2x4_ASAP7_75t_L g7094 ( 
.A(n_6037),
.B(n_4704),
.Y(n_7094)
);

AOI22x1_ASAP7_75t_L g7095 ( 
.A1(n_6077),
.A2(n_5527),
.B1(n_5217),
.B2(n_5223),
.Y(n_7095)
);

OAI21x1_ASAP7_75t_L g7096 ( 
.A1(n_5701),
.A2(n_5728),
.B(n_5727),
.Y(n_7096)
);

NAND3xp33_ASAP7_75t_L g7097 ( 
.A(n_5896),
.B(n_4830),
.C(n_4795),
.Y(n_7097)
);

NOR2xp33_ASAP7_75t_L g7098 ( 
.A(n_6038),
.B(n_5466),
.Y(n_7098)
);

OR2x2_ASAP7_75t_L g7099 ( 
.A(n_6064),
.B(n_5662),
.Y(n_7099)
);

INVx1_ASAP7_75t_L g7100 ( 
.A(n_6407),
.Y(n_7100)
);

INVx2_ASAP7_75t_L g7101 ( 
.A(n_5652),
.Y(n_7101)
);

OA21x2_ASAP7_75t_L g7102 ( 
.A1(n_6178),
.A2(n_5217),
.B(n_5209),
.Y(n_7102)
);

OAI22xp33_ASAP7_75t_L g7103 ( 
.A1(n_6286),
.A2(n_5525),
.B1(n_4789),
.B2(n_4775),
.Y(n_7103)
);

NOR2xp67_ASAP7_75t_L g7104 ( 
.A(n_6361),
.B(n_4721),
.Y(n_7104)
);

INVx2_ASAP7_75t_SL g7105 ( 
.A(n_6361),
.Y(n_7105)
);

BUFx2_ASAP7_75t_L g7106 ( 
.A(n_5568),
.Y(n_7106)
);

NAND2xp5_ASAP7_75t_L g7107 ( 
.A(n_6105),
.B(n_4798),
.Y(n_7107)
);

AND2x4_ASAP7_75t_L g7108 ( 
.A(n_6126),
.B(n_4704),
.Y(n_7108)
);

AOI22xp33_ASAP7_75t_L g7109 ( 
.A1(n_6295),
.A2(n_4855),
.B1(n_4851),
.B2(n_4775),
.Y(n_7109)
);

CKINVDCx8_ASAP7_75t_R g7110 ( 
.A(n_6165),
.Y(n_7110)
);

AND2x2_ASAP7_75t_L g7111 ( 
.A(n_6327),
.B(n_5487),
.Y(n_7111)
);

AOI22xp33_ASAP7_75t_L g7112 ( 
.A1(n_6295),
.A2(n_4775),
.B1(n_5484),
.B2(n_5266),
.Y(n_7112)
);

BUFx3_ASAP7_75t_L g7113 ( 
.A(n_5991),
.Y(n_7113)
);

AO21x2_ASAP7_75t_L g7114 ( 
.A1(n_5556),
.A2(n_5027),
.B(n_5011),
.Y(n_7114)
);

OA21x2_ASAP7_75t_L g7115 ( 
.A1(n_6186),
.A2(n_5217),
.B(n_5209),
.Y(n_7115)
);

INVx1_ASAP7_75t_L g7116 ( 
.A(n_6407),
.Y(n_7116)
);

AO21x2_ASAP7_75t_L g7117 ( 
.A1(n_6055),
.A2(n_5027),
.B(n_5011),
.Y(n_7117)
);

INVx2_ASAP7_75t_L g7118 ( 
.A(n_5653),
.Y(n_7118)
);

AOI21xp5_ASAP7_75t_L g7119 ( 
.A1(n_5648),
.A2(n_5237),
.B(n_5223),
.Y(n_7119)
);

CKINVDCx5p33_ASAP7_75t_R g7120 ( 
.A(n_5756),
.Y(n_7120)
);

INVx2_ASAP7_75t_L g7121 ( 
.A(n_5653),
.Y(n_7121)
);

NAND2x1p5_ASAP7_75t_L g7122 ( 
.A(n_5878),
.B(n_5880),
.Y(n_7122)
);

NAND2xp5_ASAP7_75t_L g7123 ( 
.A(n_6146),
.B(n_4801),
.Y(n_7123)
);

AOI22xp33_ASAP7_75t_SL g7124 ( 
.A1(n_5599),
.A2(n_5410),
.B1(n_5038),
.B2(n_4745),
.Y(n_7124)
);

OAI222xp33_ASAP7_75t_L g7125 ( 
.A1(n_5588),
.A2(n_5597),
.B1(n_5791),
.B2(n_5785),
.C1(n_5864),
.C2(n_5671),
.Y(n_7125)
);

BUFx2_ASAP7_75t_L g7126 ( 
.A(n_5568),
.Y(n_7126)
);

BUFx10_ASAP7_75t_L g7127 ( 
.A(n_6018),
.Y(n_7127)
);

INVx2_ASAP7_75t_SL g7128 ( 
.A(n_6361),
.Y(n_7128)
);

AOI21xp5_ASAP7_75t_L g7129 ( 
.A1(n_5624),
.A2(n_5879),
.B(n_5710),
.Y(n_7129)
);

AOI221xp5_ASAP7_75t_L g7130 ( 
.A1(n_6038),
.A2(n_5857),
.B1(n_5847),
.B2(n_5903),
.C(n_5896),
.Y(n_7130)
);

AO31x2_ASAP7_75t_L g7131 ( 
.A1(n_5738),
.A2(n_5206),
.A3(n_5213),
.B(n_5205),
.Y(n_7131)
);

AOI222xp33_ASAP7_75t_L g7132 ( 
.A1(n_6039),
.A2(n_4786),
.B1(n_4767),
.B2(n_4303),
.C1(n_4284),
.C2(n_4306),
.Y(n_7132)
);

INVx1_ASAP7_75t_L g7133 ( 
.A(n_6417),
.Y(n_7133)
);

INVx1_ASAP7_75t_L g7134 ( 
.A(n_6417),
.Y(n_7134)
);

OAI21xp5_ASAP7_75t_L g7135 ( 
.A1(n_6312),
.A2(n_5857),
.B(n_5847),
.Y(n_7135)
);

NOR2xp67_ASAP7_75t_L g7136 ( 
.A(n_6361),
.B(n_4721),
.Y(n_7136)
);

AOI221xp5_ASAP7_75t_L g7137 ( 
.A1(n_5903),
.A2(n_5842),
.B1(n_5853),
.B2(n_6323),
.C(n_5874),
.Y(n_7137)
);

NAND2x1p5_ASAP7_75t_L g7138 ( 
.A(n_5878),
.B(n_4721),
.Y(n_7138)
);

AOI21xp5_ASAP7_75t_L g7139 ( 
.A1(n_5624),
.A2(n_5237),
.B(n_5223),
.Y(n_7139)
);

INVx2_ASAP7_75t_L g7140 ( 
.A(n_5653),
.Y(n_7140)
);

INVx1_ASAP7_75t_L g7141 ( 
.A(n_6432),
.Y(n_7141)
);

BUFx4f_ASAP7_75t_SL g7142 ( 
.A(n_5823),
.Y(n_7142)
);

AO21x2_ASAP7_75t_L g7143 ( 
.A1(n_6055),
.A2(n_5031),
.B(n_5027),
.Y(n_7143)
);

INVx2_ASAP7_75t_L g7144 ( 
.A(n_5653),
.Y(n_7144)
);

AND2x4_ASAP7_75t_L g7145 ( 
.A(n_6126),
.B(n_4704),
.Y(n_7145)
);

AO21x2_ASAP7_75t_L g7146 ( 
.A1(n_6186),
.A2(n_5040),
.B(n_5031),
.Y(n_7146)
);

INVx1_ASAP7_75t_L g7147 ( 
.A(n_6432),
.Y(n_7147)
);

NAND2xp5_ASAP7_75t_L g7148 ( 
.A(n_6146),
.B(n_4801),
.Y(n_7148)
);

NAND2x1p5_ASAP7_75t_L g7149 ( 
.A(n_5878),
.B(n_4721),
.Y(n_7149)
);

AND2x2_ASAP7_75t_L g7150 ( 
.A(n_6327),
.B(n_5504),
.Y(n_7150)
);

INVx2_ASAP7_75t_L g7151 ( 
.A(n_5696),
.Y(n_7151)
);

OA21x2_ASAP7_75t_L g7152 ( 
.A1(n_5842),
.A2(n_5252),
.B(n_5237),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_6440),
.Y(n_7153)
);

AOI21x1_ASAP7_75t_L g7154 ( 
.A1(n_5913),
.A2(n_5268),
.B(n_5252),
.Y(n_7154)
);

INVx1_ASAP7_75t_L g7155 ( 
.A(n_6440),
.Y(n_7155)
);

OAI22xp5_ASAP7_75t_L g7156 ( 
.A1(n_6312),
.A2(n_5504),
.B1(n_5512),
.B2(n_5509),
.Y(n_7156)
);

AO21x2_ASAP7_75t_L g7157 ( 
.A1(n_5577),
.A2(n_5703),
.B(n_5700),
.Y(n_7157)
);

O2A1O1Ixp33_ASAP7_75t_SL g7158 ( 
.A1(n_5566),
.A2(n_5369),
.B(n_5535),
.C(n_4723),
.Y(n_7158)
);

AOI22xp33_ASAP7_75t_SL g7159 ( 
.A1(n_5599),
.A2(n_5410),
.B1(n_4797),
.B2(n_4817),
.Y(n_7159)
);

INVx1_ASAP7_75t_L g7160 ( 
.A(n_5661),
.Y(n_7160)
);

OAI22xp5_ASAP7_75t_L g7161 ( 
.A1(n_5631),
.A2(n_5509),
.B1(n_5512),
.B2(n_5540),
.Y(n_7161)
);

NAND3xp33_ASAP7_75t_L g7162 ( 
.A(n_6046),
.B(n_4840),
.C(n_4830),
.Y(n_7162)
);

CKINVDCx5p33_ASAP7_75t_R g7163 ( 
.A(n_5846),
.Y(n_7163)
);

INVx4_ASAP7_75t_SL g7164 ( 
.A(n_5573),
.Y(n_7164)
);

INVx2_ASAP7_75t_SL g7165 ( 
.A(n_6361),
.Y(n_7165)
);

INVx2_ASAP7_75t_SL g7166 ( 
.A(n_6126),
.Y(n_7166)
);

NAND2xp5_ASAP7_75t_L g7167 ( 
.A(n_6064),
.B(n_5874),
.Y(n_7167)
);

NAND2xp5_ASAP7_75t_L g7168 ( 
.A(n_5853),
.B(n_4801),
.Y(n_7168)
);

INVx8_ASAP7_75t_L g7169 ( 
.A(n_6405),
.Y(n_7169)
);

OAI21xp5_ASAP7_75t_L g7170 ( 
.A1(n_5608),
.A2(n_4841),
.B(n_4840),
.Y(n_7170)
);

INVx2_ASAP7_75t_L g7171 ( 
.A(n_5696),
.Y(n_7171)
);

AOI22xp33_ASAP7_75t_L g7172 ( 
.A1(n_6295),
.A2(n_4775),
.B1(n_5484),
.B2(n_4786),
.Y(n_7172)
);

INVx1_ASAP7_75t_L g7173 ( 
.A(n_5661),
.Y(n_7173)
);

INVx1_ASAP7_75t_L g7174 ( 
.A(n_5669),
.Y(n_7174)
);

O2A1O1Ixp33_ASAP7_75t_SL g7175 ( 
.A1(n_6291),
.A2(n_4723),
.B(n_5431),
.C(n_5349),
.Y(n_7175)
);

INVx1_ASAP7_75t_SL g7176 ( 
.A(n_5602),
.Y(n_7176)
);

AND2x4_ASAP7_75t_L g7177 ( 
.A(n_6126),
.B(n_4704),
.Y(n_7177)
);

OA21x2_ASAP7_75t_L g7178 ( 
.A1(n_6323),
.A2(n_5268),
.B(n_5252),
.Y(n_7178)
);

CKINVDCx16_ASAP7_75t_R g7179 ( 
.A(n_6291),
.Y(n_7179)
);

AOI21x1_ASAP7_75t_L g7180 ( 
.A1(n_5913),
.A2(n_5282),
.B(n_5268),
.Y(n_7180)
);

AOI22xp33_ASAP7_75t_L g7181 ( 
.A1(n_5785),
.A2(n_4775),
.B1(n_5484),
.B2(n_4581),
.Y(n_7181)
);

HB1xp67_ASAP7_75t_L g7182 ( 
.A(n_5978),
.Y(n_7182)
);

OAI21xp5_ASAP7_75t_L g7183 ( 
.A1(n_5608),
.A2(n_4845),
.B(n_4841),
.Y(n_7183)
);

NOR2xp33_ASAP7_75t_L g7184 ( 
.A(n_6283),
.B(n_5282),
.Y(n_7184)
);

INVx2_ASAP7_75t_L g7185 ( 
.A(n_5696),
.Y(n_7185)
);

O2A1O1Ixp33_ASAP7_75t_SL g7186 ( 
.A1(n_6074),
.A2(n_4885),
.B(n_4956),
.C(n_4736),
.Y(n_7186)
);

INVx2_ASAP7_75t_L g7187 ( 
.A(n_5696),
.Y(n_7187)
);

NOR2xp33_ASAP7_75t_L g7188 ( 
.A(n_6283),
.B(n_5282),
.Y(n_7188)
);

INVx2_ASAP7_75t_SL g7189 ( 
.A(n_6137),
.Y(n_7189)
);

O2A1O1Ixp33_ASAP7_75t_L g7190 ( 
.A1(n_6415),
.A2(n_4845),
.B(n_5322),
.C(n_5308),
.Y(n_7190)
);

INVx1_ASAP7_75t_SL g7191 ( 
.A(n_5602),
.Y(n_7191)
);

AOI22xp33_ASAP7_75t_L g7192 ( 
.A1(n_5588),
.A2(n_4775),
.B1(n_5484),
.B2(n_5410),
.Y(n_7192)
);

AO31x2_ASAP7_75t_L g7193 ( 
.A1(n_5870),
.A2(n_5213),
.A3(n_5216),
.B(n_5206),
.Y(n_7193)
);

INVx3_ASAP7_75t_L g7194 ( 
.A(n_5650),
.Y(n_7194)
);

INVx4_ASAP7_75t_SL g7195 ( 
.A(n_5573),
.Y(n_7195)
);

BUFx2_ASAP7_75t_SL g7196 ( 
.A(n_5801),
.Y(n_7196)
);

AOI22xp33_ASAP7_75t_L g7197 ( 
.A1(n_5597),
.A2(n_5484),
.B1(n_5410),
.B2(n_4541),
.Y(n_7197)
);

INVx5_ASAP7_75t_L g7198 ( 
.A(n_5573),
.Y(n_7198)
);

INVx1_ASAP7_75t_L g7199 ( 
.A(n_5669),
.Y(n_7199)
);

INVx2_ASAP7_75t_L g7200 ( 
.A(n_5700),
.Y(n_7200)
);

OAI21x1_ASAP7_75t_L g7201 ( 
.A1(n_5811),
.A2(n_5506),
.B(n_4220),
.Y(n_7201)
);

BUFx2_ASAP7_75t_L g7202 ( 
.A(n_5879),
.Y(n_7202)
);

INVx1_ASAP7_75t_L g7203 ( 
.A(n_5676),
.Y(n_7203)
);

O2A1O1Ixp33_ASAP7_75t_SL g7204 ( 
.A1(n_6074),
.A2(n_4859),
.B(n_4901),
.C(n_4736),
.Y(n_7204)
);

AOI22xp33_ASAP7_75t_L g7205 ( 
.A1(n_5864),
.A2(n_4541),
.B1(n_5489),
.B2(n_4717),
.Y(n_7205)
);

OAI21x1_ASAP7_75t_L g7206 ( 
.A1(n_5819),
.A2(n_5506),
.B(n_4220),
.Y(n_7206)
);

AO22x2_ASAP7_75t_L g7207 ( 
.A1(n_5610),
.A2(n_5656),
.B1(n_5662),
.B2(n_5681),
.Y(n_7207)
);

OA21x2_ASAP7_75t_L g7208 ( 
.A1(n_6324),
.A2(n_5322),
.B(n_5308),
.Y(n_7208)
);

AO31x2_ASAP7_75t_L g7209 ( 
.A1(n_5870),
.A2(n_6051),
.A3(n_5610),
.B(n_6273),
.Y(n_7209)
);

INVx1_ASAP7_75t_L g7210 ( 
.A(n_5676),
.Y(n_7210)
);

INVx1_ASAP7_75t_SL g7211 ( 
.A(n_5846),
.Y(n_7211)
);

INVx1_ASAP7_75t_L g7212 ( 
.A(n_5687),
.Y(n_7212)
);

OAI22xp5_ASAP7_75t_L g7213 ( 
.A1(n_5631),
.A2(n_5509),
.B1(n_5512),
.B2(n_5540),
.Y(n_7213)
);

OAI222xp33_ASAP7_75t_L g7214 ( 
.A1(n_5741),
.A2(n_5489),
.B1(n_4945),
.B2(n_4849),
.C1(n_4906),
.C2(n_4922),
.Y(n_7214)
);

BUFx2_ASAP7_75t_R g7215 ( 
.A(n_6188),
.Y(n_7215)
);

NAND2xp5_ASAP7_75t_L g7216 ( 
.A(n_6046),
.B(n_4849),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_5687),
.Y(n_7217)
);

AOI22xp33_ASAP7_75t_SL g7218 ( 
.A1(n_5599),
.A2(n_6121),
.B1(n_6211),
.B2(n_6277),
.Y(n_7218)
);

INVx3_ASAP7_75t_L g7219 ( 
.A(n_5650),
.Y(n_7219)
);

OAI21x1_ASAP7_75t_L g7220 ( 
.A1(n_5819),
.A2(n_5506),
.B(n_4220),
.Y(n_7220)
);

AOI21xp5_ASAP7_75t_L g7221 ( 
.A1(n_6324),
.A2(n_5322),
.B(n_5308),
.Y(n_7221)
);

OAI22xp5_ASAP7_75t_L g7222 ( 
.A1(n_5658),
.A2(n_5540),
.B1(n_4688),
.B2(n_5355),
.Y(n_7222)
);

OR2x6_ASAP7_75t_L g7223 ( 
.A(n_6244),
.B(n_5489),
.Y(n_7223)
);

CKINVDCx20_ASAP7_75t_R g7224 ( 
.A(n_5758),
.Y(n_7224)
);

OA21x2_ASAP7_75t_L g7225 ( 
.A1(n_5665),
.A2(n_5355),
.B(n_5326),
.Y(n_7225)
);

INVx1_ASAP7_75t_L g7226 ( 
.A(n_5709),
.Y(n_7226)
);

INVx1_ASAP7_75t_L g7227 ( 
.A(n_5709),
.Y(n_7227)
);

OAI21x1_ASAP7_75t_SL g7228 ( 
.A1(n_6073),
.A2(n_5363),
.B(n_5360),
.Y(n_7228)
);

INVx1_ASAP7_75t_L g7229 ( 
.A(n_5712),
.Y(n_7229)
);

AND2x2_ASAP7_75t_L g7230 ( 
.A(n_5821),
.B(n_5326),
.Y(n_7230)
);

INVx1_ASAP7_75t_L g7231 ( 
.A(n_5712),
.Y(n_7231)
);

INVx1_ASAP7_75t_L g7232 ( 
.A(n_5724),
.Y(n_7232)
);

INVx2_ASAP7_75t_L g7233 ( 
.A(n_5700),
.Y(n_7233)
);

NOR2x1_ASAP7_75t_R g7234 ( 
.A(n_6033),
.B(n_4724),
.Y(n_7234)
);

BUFx3_ASAP7_75t_L g7235 ( 
.A(n_6033),
.Y(n_7235)
);

HB1xp67_ASAP7_75t_L g7236 ( 
.A(n_5978),
.Y(n_7236)
);

NOR2xp67_ASAP7_75t_SL g7237 ( 
.A(n_6418),
.B(n_4724),
.Y(n_7237)
);

AND2x2_ASAP7_75t_L g7238 ( 
.A(n_5821),
.B(n_5326),
.Y(n_7238)
);

INVx1_ASAP7_75t_L g7239 ( 
.A(n_5724),
.Y(n_7239)
);

AOI22xp33_ASAP7_75t_L g7240 ( 
.A1(n_5658),
.A2(n_5489),
.B1(n_4717),
.B2(n_4678),
.Y(n_7240)
);

INVx1_ASAP7_75t_L g7241 ( 
.A(n_5734),
.Y(n_7241)
);

HB1xp67_ASAP7_75t_L g7242 ( 
.A(n_6009),
.Y(n_7242)
);

O2A1O1Ixp33_ASAP7_75t_L g7243 ( 
.A1(n_6047),
.A2(n_5656),
.B(n_5993),
.C(n_5577),
.Y(n_7243)
);

OA21x2_ASAP7_75t_L g7244 ( 
.A1(n_5665),
.A2(n_5357),
.B(n_5355),
.Y(n_7244)
);

INVx3_ASAP7_75t_L g7245 ( 
.A(n_5650),
.Y(n_7245)
);

AND2x4_ASAP7_75t_L g7246 ( 
.A(n_6137),
.B(n_4761),
.Y(n_7246)
);

INVx2_ASAP7_75t_L g7247 ( 
.A(n_5700),
.Y(n_7247)
);

OAI21x1_ASAP7_75t_SL g7248 ( 
.A1(n_6073),
.A2(n_5363),
.B(n_5360),
.Y(n_7248)
);

AO21x2_ASAP7_75t_L g7249 ( 
.A1(n_5703),
.A2(n_5040),
.B(n_5031),
.Y(n_7249)
);

BUFx3_ASAP7_75t_L g7250 ( 
.A(n_6033),
.Y(n_7250)
);

OAI21x1_ASAP7_75t_L g7251 ( 
.A1(n_5826),
.A2(n_5871),
.B(n_5840),
.Y(n_7251)
);

AND2x2_ASAP7_75t_L g7252 ( 
.A(n_5821),
.B(n_5357),
.Y(n_7252)
);

AOI21xp5_ASAP7_75t_L g7253 ( 
.A1(n_6281),
.A2(n_5370),
.B(n_5357),
.Y(n_7253)
);

INVx1_ASAP7_75t_L g7254 ( 
.A(n_5734),
.Y(n_7254)
);

INVx1_ASAP7_75t_L g7255 ( 
.A(n_5761),
.Y(n_7255)
);

INVx2_ASAP7_75t_L g7256 ( 
.A(n_5731),
.Y(n_7256)
);

NAND2x1_ASAP7_75t_L g7257 ( 
.A(n_6104),
.B(n_5370),
.Y(n_7257)
);

AO31x2_ASAP7_75t_L g7258 ( 
.A1(n_5870),
.A2(n_5229),
.A3(n_5234),
.B(n_5216),
.Y(n_7258)
);

INVx2_ASAP7_75t_L g7259 ( 
.A(n_5731),
.Y(n_7259)
);

AO21x2_ASAP7_75t_L g7260 ( 
.A1(n_5731),
.A2(n_5047),
.B(n_5040),
.Y(n_7260)
);

OAI21x1_ASAP7_75t_L g7261 ( 
.A1(n_5826),
.A2(n_4766),
.B(n_4761),
.Y(n_7261)
);

INVx2_ASAP7_75t_L g7262 ( 
.A(n_5731),
.Y(n_7262)
);

INVx1_ASAP7_75t_L g7263 ( 
.A(n_5761),
.Y(n_7263)
);

OAI21x1_ASAP7_75t_L g7264 ( 
.A1(n_5826),
.A2(n_4834),
.B(n_4766),
.Y(n_7264)
);

OAI22xp5_ASAP7_75t_L g7265 ( 
.A1(n_5801),
.A2(n_4688),
.B1(n_5420),
.B2(n_5370),
.Y(n_7265)
);

INVx1_ASAP7_75t_L g7266 ( 
.A(n_5773),
.Y(n_7266)
);

INVx2_ASAP7_75t_L g7267 ( 
.A(n_5737),
.Y(n_7267)
);

INVx1_ASAP7_75t_L g7268 ( 
.A(n_5773),
.Y(n_7268)
);

NAND2xp5_ASAP7_75t_L g7269 ( 
.A(n_6047),
.B(n_4849),
.Y(n_7269)
);

OAI21xp5_ASAP7_75t_L g7270 ( 
.A1(n_6219),
.A2(n_5420),
.B(n_4957),
.Y(n_7270)
);

AOI22xp33_ASAP7_75t_L g7271 ( 
.A1(n_5741),
.A2(n_6277),
.B1(n_5960),
.B2(n_6441),
.Y(n_7271)
);

AOI22xp33_ASAP7_75t_SL g7272 ( 
.A1(n_6121),
.A2(n_4797),
.B1(n_4817),
.B2(n_4745),
.Y(n_7272)
);

NOR2xp67_ASAP7_75t_L g7273 ( 
.A(n_5878),
.B(n_4850),
.Y(n_7273)
);

AO21x2_ASAP7_75t_L g7274 ( 
.A1(n_5737),
.A2(n_5050),
.B(n_5047),
.Y(n_7274)
);

OAI21x1_ASAP7_75t_SL g7275 ( 
.A1(n_6051),
.A2(n_6156),
.B(n_6130),
.Y(n_7275)
);

INVx2_ASAP7_75t_L g7276 ( 
.A(n_5737),
.Y(n_7276)
);

INVx2_ASAP7_75t_R g7277 ( 
.A(n_5957),
.Y(n_7277)
);

OAI21xp5_ASAP7_75t_L g7278 ( 
.A1(n_6219),
.A2(n_5420),
.B(n_4957),
.Y(n_7278)
);

OA21x2_ASAP7_75t_L g7279 ( 
.A1(n_5678),
.A2(n_4998),
.B(n_5047),
.Y(n_7279)
);

AO21x2_ASAP7_75t_L g7280 ( 
.A1(n_5737),
.A2(n_5054),
.B(n_5050),
.Y(n_7280)
);

INVx1_ASAP7_75t_L g7281 ( 
.A(n_5775),
.Y(n_7281)
);

OAI21x1_ASAP7_75t_SL g7282 ( 
.A1(n_6051),
.A2(n_5363),
.B(n_5360),
.Y(n_7282)
);

AO31x2_ASAP7_75t_L g7283 ( 
.A1(n_6273),
.A2(n_5234),
.A3(n_5238),
.B(n_5229),
.Y(n_7283)
);

BUFx3_ASAP7_75t_L g7284 ( 
.A(n_6033),
.Y(n_7284)
);

INVx3_ASAP7_75t_L g7285 ( 
.A(n_5650),
.Y(n_7285)
);

OAI22xp5_ASAP7_75t_L g7286 ( 
.A1(n_5801),
.A2(n_4688),
.B1(n_5043),
.B2(n_5363),
.Y(n_7286)
);

AO21x2_ASAP7_75t_L g7287 ( 
.A1(n_5743),
.A2(n_5054),
.B(n_5050),
.Y(n_7287)
);

AOI22xp33_ASAP7_75t_SL g7288 ( 
.A1(n_6121),
.A2(n_4797),
.B1(n_4817),
.B2(n_4745),
.Y(n_7288)
);

AOI22xp33_ASAP7_75t_L g7289 ( 
.A1(n_5960),
.A2(n_4717),
.B1(n_4678),
.B2(n_4358),
.Y(n_7289)
);

INVx1_ASAP7_75t_L g7290 ( 
.A(n_5775),
.Y(n_7290)
);

INVx4_ASAP7_75t_L g7291 ( 
.A(n_6293),
.Y(n_7291)
);

INVx2_ASAP7_75t_L g7292 ( 
.A(n_5743),
.Y(n_7292)
);

AOI21x1_ASAP7_75t_L g7293 ( 
.A1(n_5913),
.A2(n_5061),
.B(n_5054),
.Y(n_7293)
);

AND2x4_ASAP7_75t_L g7294 ( 
.A(n_6137),
.B(n_4913),
.Y(n_7294)
);

AND2x2_ASAP7_75t_L g7295 ( 
.A(n_6012),
.B(n_6211),
.Y(n_7295)
);

OA21x2_ASAP7_75t_L g7296 ( 
.A1(n_5678),
.A2(n_4998),
.B(n_5061),
.Y(n_7296)
);

OAI22xp5_ASAP7_75t_L g7297 ( 
.A1(n_5814),
.A2(n_5043),
.B1(n_5438),
.B2(n_4757),
.Y(n_7297)
);

AOI22xp33_ASAP7_75t_L g7298 ( 
.A1(n_5960),
.A2(n_4678),
.B1(n_4358),
.B2(n_4379),
.Y(n_7298)
);

AOI21x1_ASAP7_75t_L g7299 ( 
.A1(n_5919),
.A2(n_5066),
.B(n_5061),
.Y(n_7299)
);

INVx2_ASAP7_75t_L g7300 ( 
.A(n_5743),
.Y(n_7300)
);

AND2x4_ASAP7_75t_L g7301 ( 
.A(n_6137),
.B(n_4913),
.Y(n_7301)
);

CKINVDCx5p33_ASAP7_75t_R g7302 ( 
.A(n_5899),
.Y(n_7302)
);

NOR3xp33_ASAP7_75t_L g7303 ( 
.A(n_5627),
.B(n_5244),
.C(n_5238),
.Y(n_7303)
);

INVx2_ASAP7_75t_L g7304 ( 
.A(n_5743),
.Y(n_7304)
);

AO21x2_ASAP7_75t_L g7305 ( 
.A1(n_5744),
.A2(n_5070),
.B(n_5066),
.Y(n_7305)
);

BUFx3_ASAP7_75t_L g7306 ( 
.A(n_6188),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_5786),
.Y(n_7307)
);

A2O1A1Ixp33_ASAP7_75t_L g7308 ( 
.A1(n_6121),
.A2(n_5751),
.B(n_5668),
.C(n_6079),
.Y(n_7308)
);

A2O1A1Ixp33_ASAP7_75t_L g7309 ( 
.A1(n_5751),
.A2(n_4678),
.B(n_4998),
.C(n_4740),
.Y(n_7309)
);

OR2x2_ASAP7_75t_L g7310 ( 
.A(n_5662),
.B(n_4874),
.Y(n_7310)
);

INVx2_ASAP7_75t_L g7311 ( 
.A(n_5744),
.Y(n_7311)
);

AOI221xp5_ASAP7_75t_L g7312 ( 
.A1(n_5993),
.A2(n_5539),
.B1(n_5256),
.B2(n_5257),
.C(n_5250),
.Y(n_7312)
);

INVx8_ASAP7_75t_L g7313 ( 
.A(n_6418),
.Y(n_7313)
);

NAND2x1p5_ASAP7_75t_L g7314 ( 
.A(n_5878),
.B(n_4850),
.Y(n_7314)
);

OAI21xp5_ASAP7_75t_L g7315 ( 
.A1(n_6219),
.A2(n_6202),
.B(n_6233),
.Y(n_7315)
);

AOI221xp5_ASAP7_75t_L g7316 ( 
.A1(n_6434),
.A2(n_5539),
.B1(n_5256),
.B2(n_5257),
.C(n_5250),
.Y(n_7316)
);

AOI221xp5_ASAP7_75t_L g7317 ( 
.A1(n_6434),
.A2(n_5679),
.B1(n_6425),
.B2(n_6296),
.C(n_5685),
.Y(n_7317)
);

HB1xp67_ASAP7_75t_L g7318 ( 
.A(n_6009),
.Y(n_7318)
);

AND2x4_ASAP7_75t_L g7319 ( 
.A(n_6138),
.B(n_4938),
.Y(n_7319)
);

AOI21xp5_ASAP7_75t_L g7320 ( 
.A1(n_6281),
.A2(n_4723),
.B(n_4714),
.Y(n_7320)
);

BUFx2_ASAP7_75t_L g7321 ( 
.A(n_6211),
.Y(n_7321)
);

NAND2xp5_ASAP7_75t_L g7322 ( 
.A(n_5904),
.B(n_4874),
.Y(n_7322)
);

OA21x2_ASAP7_75t_L g7323 ( 
.A1(n_5681),
.A2(n_4998),
.B(n_5066),
.Y(n_7323)
);

AOI21x1_ASAP7_75t_L g7324 ( 
.A1(n_5919),
.A2(n_5970),
.B(n_5925),
.Y(n_7324)
);

OR2x2_ASAP7_75t_L g7325 ( 
.A(n_5745),
.B(n_4874),
.Y(n_7325)
);

AOI221xp5_ASAP7_75t_L g7326 ( 
.A1(n_5679),
.A2(n_5534),
.B1(n_5519),
.B2(n_5515),
.C(n_5288),
.Y(n_7326)
);

INVx2_ASAP7_75t_L g7327 ( 
.A(n_5744),
.Y(n_7327)
);

INVx1_ASAP7_75t_L g7328 ( 
.A(n_5786),
.Y(n_7328)
);

NAND2x1_ASAP7_75t_L g7329 ( 
.A(n_6104),
.B(n_4968),
.Y(n_7329)
);

NAND2xp5_ASAP7_75t_L g7330 ( 
.A(n_5904),
.B(n_4906),
.Y(n_7330)
);

OAI22xp5_ASAP7_75t_L g7331 ( 
.A1(n_5814),
.A2(n_5438),
.B1(n_4757),
.B2(n_4835),
.Y(n_7331)
);

AOI22xp33_ASAP7_75t_L g7332 ( 
.A1(n_5960),
.A2(n_4678),
.B1(n_4358),
.B2(n_4379),
.Y(n_7332)
);

AOI22xp33_ASAP7_75t_L g7333 ( 
.A1(n_5960),
.A2(n_4379),
.B1(n_4430),
.B2(n_4348),
.Y(n_7333)
);

AND2x2_ASAP7_75t_L g7334 ( 
.A(n_6012),
.B(n_5017),
.Y(n_7334)
);

INVx1_ASAP7_75t_L g7335 ( 
.A(n_5813),
.Y(n_7335)
);

AOI21xp5_ASAP7_75t_L g7336 ( 
.A1(n_6024),
.A2(n_5660),
.B(n_6202),
.Y(n_7336)
);

AO31x2_ASAP7_75t_L g7337 ( 
.A1(n_6278),
.A2(n_5258),
.A3(n_5288),
.B(n_5244),
.Y(n_7337)
);

OA21x2_ASAP7_75t_L g7338 ( 
.A1(n_5685),
.A2(n_6057),
.B(n_6048),
.Y(n_7338)
);

INVx1_ASAP7_75t_L g7339 ( 
.A(n_5813),
.Y(n_7339)
);

INVx1_ASAP7_75t_L g7340 ( 
.A(n_5825),
.Y(n_7340)
);

AND2x4_ASAP7_75t_L g7341 ( 
.A(n_6138),
.B(n_6142),
.Y(n_7341)
);

AO31x2_ASAP7_75t_L g7342 ( 
.A1(n_6278),
.A2(n_5321),
.A3(n_5323),
.B(n_5258),
.Y(n_7342)
);

AND2x4_ASAP7_75t_L g7343 ( 
.A(n_6138),
.B(n_6142),
.Y(n_7343)
);

O2A1O1Ixp33_ASAP7_75t_L g7344 ( 
.A1(n_6233),
.A2(n_5323),
.B(n_5327),
.C(n_5321),
.Y(n_7344)
);

AOI22xp33_ASAP7_75t_L g7345 ( 
.A1(n_5960),
.A2(n_4430),
.B1(n_4439),
.B2(n_4348),
.Y(n_7345)
);

NOR2xp33_ASAP7_75t_R g7346 ( 
.A(n_5716),
.B(n_4853),
.Y(n_7346)
);

INVx3_ASAP7_75t_L g7347 ( 
.A(n_5666),
.Y(n_7347)
);

AOI22xp33_ASAP7_75t_L g7348 ( 
.A1(n_5960),
.A2(n_6277),
.B1(n_6441),
.B2(n_5668),
.Y(n_7348)
);

AO21x2_ASAP7_75t_L g7349 ( 
.A1(n_5744),
.A2(n_5076),
.B(n_5070),
.Y(n_7349)
);

OAI21xp5_ASAP7_75t_L g7350 ( 
.A1(n_6219),
.A2(n_4960),
.B(n_4947),
.Y(n_7350)
);

OAI21xp5_ASAP7_75t_L g7351 ( 
.A1(n_6008),
.A2(n_4960),
.B(n_4947),
.Y(n_7351)
);

NAND2xp5_ASAP7_75t_L g7352 ( 
.A(n_5908),
.B(n_4906),
.Y(n_7352)
);

INVx1_ASAP7_75t_L g7353 ( 
.A(n_5825),
.Y(n_7353)
);

OAI21xp5_ASAP7_75t_L g7354 ( 
.A1(n_6008),
.A2(n_5790),
.B(n_5759),
.Y(n_7354)
);

AO21x2_ASAP7_75t_L g7355 ( 
.A1(n_5749),
.A2(n_5076),
.B(n_5070),
.Y(n_7355)
);

INVx2_ASAP7_75t_L g7356 ( 
.A(n_5749),
.Y(n_7356)
);

OA21x2_ASAP7_75t_L g7357 ( 
.A1(n_6048),
.A2(n_4998),
.B(n_5076),
.Y(n_7357)
);

INVx2_ASAP7_75t_L g7358 ( 
.A(n_5749),
.Y(n_7358)
);

OAI21x1_ASAP7_75t_L g7359 ( 
.A1(n_5893),
.A2(n_5937),
.B(n_5935),
.Y(n_7359)
);

HB1xp67_ASAP7_75t_L g7360 ( 
.A(n_5574),
.Y(n_7360)
);

NAND2xp5_ASAP7_75t_L g7361 ( 
.A(n_5908),
.B(n_4922),
.Y(n_7361)
);

AO21x2_ASAP7_75t_L g7362 ( 
.A1(n_5749),
.A2(n_5767),
.B(n_5763),
.Y(n_7362)
);

NAND2xp5_ASAP7_75t_L g7363 ( 
.A(n_5922),
.B(n_4922),
.Y(n_7363)
);

AND2x4_ASAP7_75t_L g7364 ( 
.A(n_6138),
.B(n_5088),
.Y(n_7364)
);

AND2x4_ASAP7_75t_L g7365 ( 
.A(n_6142),
.B(n_5088),
.Y(n_7365)
);

INVx2_ASAP7_75t_L g7366 ( 
.A(n_5763),
.Y(n_7366)
);

OA21x2_ASAP7_75t_L g7367 ( 
.A1(n_6057),
.A2(n_5080),
.B(n_5078),
.Y(n_7367)
);

AO21x2_ASAP7_75t_L g7368 ( 
.A1(n_5763),
.A2(n_5080),
.B(n_5078),
.Y(n_7368)
);

INVx1_ASAP7_75t_L g7369 ( 
.A(n_5829),
.Y(n_7369)
);

AOI22xp33_ASAP7_75t_L g7370 ( 
.A1(n_5960),
.A2(n_4439),
.B1(n_4488),
.B2(n_4430),
.Y(n_7370)
);

NAND2xp5_ASAP7_75t_SL g7371 ( 
.A(n_5861),
.B(n_5203),
.Y(n_7371)
);

OAI21xp5_ASAP7_75t_L g7372 ( 
.A1(n_5759),
.A2(n_4969),
.B(n_4964),
.Y(n_7372)
);

INVxp67_ASAP7_75t_L g7373 ( 
.A(n_6206),
.Y(n_7373)
);

AOI22xp33_ASAP7_75t_L g7374 ( 
.A1(n_5960),
.A2(n_4488),
.B1(n_4497),
.B2(n_4439),
.Y(n_7374)
);

NAND2xp5_ASAP7_75t_L g7375 ( 
.A(n_5922),
.B(n_4976),
.Y(n_7375)
);

CKINVDCx16_ASAP7_75t_R g7376 ( 
.A(n_5716),
.Y(n_7376)
);

NAND2x1p5_ASAP7_75t_L g7377 ( 
.A(n_5878),
.B(n_4850),
.Y(n_7377)
);

AO21x2_ASAP7_75t_L g7378 ( 
.A1(n_5767),
.A2(n_5105),
.B(n_5092),
.Y(n_7378)
);

AO31x2_ASAP7_75t_L g7379 ( 
.A1(n_6007),
.A2(n_5343),
.A3(n_5345),
.B(n_5327),
.Y(n_7379)
);

INVx1_ASAP7_75t_L g7380 ( 
.A(n_5829),
.Y(n_7380)
);

NOR3xp33_ASAP7_75t_SL g7381 ( 
.A(n_5897),
.B(n_5968),
.C(n_5952),
.Y(n_7381)
);

BUFx12f_ASAP7_75t_L g7382 ( 
.A(n_5823),
.Y(n_7382)
);

INVx1_ASAP7_75t_L g7383 ( 
.A(n_5838),
.Y(n_7383)
);

BUFx2_ASAP7_75t_L g7384 ( 
.A(n_6211),
.Y(n_7384)
);

NAND2xp5_ASAP7_75t_L g7385 ( 
.A(n_5745),
.B(n_4976),
.Y(n_7385)
);

NOR2xp67_ASAP7_75t_L g7386 ( 
.A(n_5880),
.B(n_4850),
.Y(n_7386)
);

NAND2xp5_ASAP7_75t_L g7387 ( 
.A(n_5766),
.B(n_4976),
.Y(n_7387)
);

HB1xp67_ASAP7_75t_L g7388 ( 
.A(n_5574),
.Y(n_7388)
);

CKINVDCx14_ASAP7_75t_R g7389 ( 
.A(n_5754),
.Y(n_7389)
);

AOI22xp33_ASAP7_75t_L g7390 ( 
.A1(n_5960),
.A2(n_6277),
.B1(n_5911),
.B2(n_5946),
.Y(n_7390)
);

INVx1_ASAP7_75t_L g7391 ( 
.A(n_5838),
.Y(n_7391)
);

AND2x2_ASAP7_75t_L g7392 ( 
.A(n_6012),
.B(n_5097),
.Y(n_7392)
);

AOI221xp5_ASAP7_75t_L g7393 ( 
.A1(n_6296),
.A2(n_5361),
.B1(n_5365),
.B2(n_5345),
.C(n_5343),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_5854),
.Y(n_7394)
);

AOI21xp5_ASAP7_75t_L g7395 ( 
.A1(n_6024),
.A2(n_4736),
.B(n_4714),
.Y(n_7395)
);

INVx1_ASAP7_75t_L g7396 ( 
.A(n_5854),
.Y(n_7396)
);

NOR2xp67_ASAP7_75t_L g7397 ( 
.A(n_5880),
.B(n_4850),
.Y(n_7397)
);

NOR2xp33_ASAP7_75t_SL g7398 ( 
.A(n_6431),
.B(n_5438),
.Y(n_7398)
);

INVx2_ASAP7_75t_L g7399 ( 
.A(n_5767),
.Y(n_7399)
);

OA21x2_ASAP7_75t_L g7400 ( 
.A1(n_6060),
.A2(n_5105),
.B(n_5092),
.Y(n_7400)
);

OAI22xp5_ASAP7_75t_L g7401 ( 
.A1(n_5814),
.A2(n_5438),
.B1(n_4757),
.B2(n_4835),
.Y(n_7401)
);

OAI21xp5_ASAP7_75t_L g7402 ( 
.A1(n_5790),
.A2(n_4969),
.B(n_4964),
.Y(n_7402)
);

AND2x2_ASAP7_75t_L g7403 ( 
.A(n_6211),
.B(n_5097),
.Y(n_7403)
);

OAI21xp5_ASAP7_75t_L g7404 ( 
.A1(n_5934),
.A2(n_6045),
.B(n_5954),
.Y(n_7404)
);

INVx1_ASAP7_75t_L g7405 ( 
.A(n_5866),
.Y(n_7405)
);

OA21x2_ASAP7_75t_L g7406 ( 
.A1(n_6060),
.A2(n_5105),
.B(n_5092),
.Y(n_7406)
);

AOI21xp5_ASAP7_75t_L g7407 ( 
.A1(n_5660),
.A2(n_4859),
.B(n_4714),
.Y(n_7407)
);

AO21x2_ASAP7_75t_L g7408 ( 
.A1(n_5767),
.A2(n_5119),
.B(n_5113),
.Y(n_7408)
);

NAND2xp5_ASAP7_75t_L g7409 ( 
.A(n_5766),
.B(n_4971),
.Y(n_7409)
);

AOI22xp5_ASAP7_75t_L g7410 ( 
.A1(n_5818),
.A2(n_4497),
.B1(n_4506),
.B2(n_4488),
.Y(n_7410)
);

AOI22xp33_ASAP7_75t_SL g7411 ( 
.A1(n_7321),
.A2(n_6211),
.B1(n_6277),
.B2(n_5960),
.Y(n_7411)
);

BUFx3_ASAP7_75t_L g7412 ( 
.A(n_6667),
.Y(n_7412)
);

CKINVDCx20_ASAP7_75t_R g7413 ( 
.A(n_6991),
.Y(n_7413)
);

OR2x2_ASAP7_75t_L g7414 ( 
.A(n_7321),
.B(n_5779),
.Y(n_7414)
);

BUFx3_ASAP7_75t_L g7415 ( 
.A(n_6667),
.Y(n_7415)
);

OAI21xp33_ASAP7_75t_L g7416 ( 
.A1(n_6536),
.A2(n_6211),
.B(n_6153),
.Y(n_7416)
);

INVx1_ASAP7_75t_L g7417 ( 
.A(n_6442),
.Y(n_7417)
);

BUFx3_ASAP7_75t_L g7418 ( 
.A(n_6667),
.Y(n_7418)
);

INVx1_ASAP7_75t_L g7419 ( 
.A(n_6442),
.Y(n_7419)
);

OAI22xp33_ASAP7_75t_L g7420 ( 
.A1(n_7321),
.A2(n_6079),
.B1(n_6083),
.B2(n_5930),
.Y(n_7420)
);

INVxp67_ASAP7_75t_SL g7421 ( 
.A(n_6956),
.Y(n_7421)
);

OR2x6_ASAP7_75t_L g7422 ( 
.A(n_6445),
.B(n_6124),
.Y(n_7422)
);

INVx3_ASAP7_75t_L g7423 ( 
.A(n_6855),
.Y(n_7423)
);

AO21x1_ASAP7_75t_SL g7424 ( 
.A1(n_6571),
.A2(n_6092),
.B(n_6078),
.Y(n_7424)
);

INVx1_ASAP7_75t_L g7425 ( 
.A(n_6446),
.Y(n_7425)
);

OAI22xp33_ASAP7_75t_L g7426 ( 
.A1(n_7384),
.A2(n_6083),
.B1(n_5930),
.B2(n_6241),
.Y(n_7426)
);

OAI21x1_ASAP7_75t_L g7427 ( 
.A1(n_6808),
.A2(n_5949),
.B(n_5937),
.Y(n_7427)
);

INVx2_ASAP7_75t_L g7428 ( 
.A(n_7293),
.Y(n_7428)
);

INVx2_ASAP7_75t_L g7429 ( 
.A(n_7293),
.Y(n_7429)
);

AOI22xp33_ASAP7_75t_L g7430 ( 
.A1(n_7384),
.A2(n_6277),
.B1(n_5911),
.B2(n_5946),
.Y(n_7430)
);

AOI21x1_ASAP7_75t_L g7431 ( 
.A1(n_6565),
.A2(n_5925),
.B(n_5919),
.Y(n_7431)
);

INVx2_ASAP7_75t_L g7432 ( 
.A(n_7299),
.Y(n_7432)
);

BUFx2_ASAP7_75t_L g7433 ( 
.A(n_6467),
.Y(n_7433)
);

HB1xp67_ASAP7_75t_L g7434 ( 
.A(n_7051),
.Y(n_7434)
);

AOI22xp33_ASAP7_75t_L g7435 ( 
.A1(n_7384),
.A2(n_6531),
.B1(n_6618),
.B2(n_6449),
.Y(n_7435)
);

AOI21x1_ASAP7_75t_L g7436 ( 
.A1(n_6565),
.A2(n_5970),
.B(n_5925),
.Y(n_7436)
);

INVx1_ASAP7_75t_SL g7437 ( 
.A(n_6538),
.Y(n_7437)
);

BUFx3_ASAP7_75t_L g7438 ( 
.A(n_6780),
.Y(n_7438)
);

AOI22xp33_ASAP7_75t_L g7439 ( 
.A1(n_6531),
.A2(n_6277),
.B1(n_5911),
.B2(n_5946),
.Y(n_7439)
);

INVx1_ASAP7_75t_L g7440 ( 
.A(n_6446),
.Y(n_7440)
);

INVx1_ASAP7_75t_L g7441 ( 
.A(n_6459),
.Y(n_7441)
);

INVx1_ASAP7_75t_L g7442 ( 
.A(n_6459),
.Y(n_7442)
);

INVx1_ASAP7_75t_L g7443 ( 
.A(n_6464),
.Y(n_7443)
);

OAI21x1_ASAP7_75t_L g7444 ( 
.A1(n_6808),
.A2(n_6986),
.B(n_6476),
.Y(n_7444)
);

NAND2xp5_ASAP7_75t_L g7445 ( 
.A(n_7077),
.B(n_6425),
.Y(n_7445)
);

HB1xp67_ASAP7_75t_L g7446 ( 
.A(n_7051),
.Y(n_7446)
);

INVx2_ASAP7_75t_L g7447 ( 
.A(n_7299),
.Y(n_7447)
);

INVx2_ASAP7_75t_L g7448 ( 
.A(n_7323),
.Y(n_7448)
);

BUFx6f_ASAP7_75t_L g7449 ( 
.A(n_6780),
.Y(n_7449)
);

NAND2x1p5_ASAP7_75t_L g7450 ( 
.A(n_7198),
.B(n_5880),
.Y(n_7450)
);

INVx1_ASAP7_75t_L g7451 ( 
.A(n_6464),
.Y(n_7451)
);

AND2x2_ASAP7_75t_L g7452 ( 
.A(n_7091),
.B(n_6238),
.Y(n_7452)
);

INVx1_ASAP7_75t_L g7453 ( 
.A(n_6466),
.Y(n_7453)
);

INVx2_ASAP7_75t_L g7454 ( 
.A(n_7323),
.Y(n_7454)
);

AND2x2_ASAP7_75t_L g7455 ( 
.A(n_7091),
.B(n_6238),
.Y(n_7455)
);

INVx1_ASAP7_75t_L g7456 ( 
.A(n_6466),
.Y(n_7456)
);

INVx3_ASAP7_75t_L g7457 ( 
.A(n_6855),
.Y(n_7457)
);

INVx2_ASAP7_75t_SL g7458 ( 
.A(n_7376),
.Y(n_7458)
);

AOI22xp33_ASAP7_75t_L g7459 ( 
.A1(n_6618),
.A2(n_6277),
.B1(n_5911),
.B2(n_5946),
.Y(n_7459)
);

INVx2_ASAP7_75t_L g7460 ( 
.A(n_7323),
.Y(n_7460)
);

INVx2_ASAP7_75t_L g7461 ( 
.A(n_7323),
.Y(n_7461)
);

INVx4_ASAP7_75t_L g7462 ( 
.A(n_6780),
.Y(n_7462)
);

BUFx2_ASAP7_75t_L g7463 ( 
.A(n_6467),
.Y(n_7463)
);

AOI22xp33_ASAP7_75t_SL g7464 ( 
.A1(n_6746),
.A2(n_6277),
.B1(n_5946),
.B2(n_5911),
.Y(n_7464)
);

INVx1_ASAP7_75t_L g7465 ( 
.A(n_6482),
.Y(n_7465)
);

AOI21x1_ASAP7_75t_L g7466 ( 
.A1(n_7091),
.A2(n_6010),
.B(n_5970),
.Y(n_7466)
);

OAI22xp33_ASAP7_75t_L g7467 ( 
.A1(n_6480),
.A2(n_6241),
.B1(n_6251),
.B2(n_6286),
.Y(n_7467)
);

AND2x2_ASAP7_75t_L g7468 ( 
.A(n_7403),
.B(n_7295),
.Y(n_7468)
);

AOI21x1_ASAP7_75t_L g7469 ( 
.A1(n_6651),
.A2(n_6112),
.B(n_6010),
.Y(n_7469)
);

INVx2_ASAP7_75t_L g7470 ( 
.A(n_6669),
.Y(n_7470)
);

NAND2x1p5_ASAP7_75t_L g7471 ( 
.A(n_7198),
.B(n_5880),
.Y(n_7471)
);

BUFx2_ASAP7_75t_L g7472 ( 
.A(n_6521),
.Y(n_7472)
);

AOI22xp33_ASAP7_75t_L g7473 ( 
.A1(n_6449),
.A2(n_6277),
.B1(n_5911),
.B2(n_5946),
.Y(n_7473)
);

BUFx12f_ASAP7_75t_L g7474 ( 
.A(n_6538),
.Y(n_7474)
);

AND2x4_ASAP7_75t_L g7475 ( 
.A(n_6506),
.B(n_6142),
.Y(n_7475)
);

INVx2_ASAP7_75t_L g7476 ( 
.A(n_7323),
.Y(n_7476)
);

INVx2_ASAP7_75t_L g7477 ( 
.A(n_7279),
.Y(n_7477)
);

INVx1_ASAP7_75t_L g7478 ( 
.A(n_6482),
.Y(n_7478)
);

AOI21x1_ASAP7_75t_L g7479 ( 
.A1(n_6651),
.A2(n_6112),
.B(n_6010),
.Y(n_7479)
);

INVx2_ASAP7_75t_L g7480 ( 
.A(n_6669),
.Y(n_7480)
);

INVx2_ASAP7_75t_L g7481 ( 
.A(n_6669),
.Y(n_7481)
);

AOI22xp33_ASAP7_75t_L g7482 ( 
.A1(n_6449),
.A2(n_6277),
.B1(n_5911),
.B2(n_5946),
.Y(n_7482)
);

INVx2_ASAP7_75t_L g7483 ( 
.A(n_6669),
.Y(n_7483)
);

INVx1_ASAP7_75t_L g7484 ( 
.A(n_6485),
.Y(n_7484)
);

OAI21x1_ASAP7_75t_SL g7485 ( 
.A1(n_6801),
.A2(n_6130),
.B(n_6122),
.Y(n_7485)
);

AOI22xp33_ASAP7_75t_L g7486 ( 
.A1(n_6651),
.A2(n_5911),
.B1(n_5946),
.B2(n_6124),
.Y(n_7486)
);

OA21x2_ASAP7_75t_L g7487 ( 
.A1(n_6702),
.A2(n_5954),
.B(n_5934),
.Y(n_7487)
);

AOI22xp5_ASAP7_75t_L g7488 ( 
.A1(n_6451),
.A2(n_5818),
.B1(n_5714),
.B2(n_5688),
.Y(n_7488)
);

INVx3_ASAP7_75t_L g7489 ( 
.A(n_6855),
.Y(n_7489)
);

AOI21xp5_ASAP7_75t_L g7490 ( 
.A1(n_6571),
.A2(n_5603),
.B(n_5547),
.Y(n_7490)
);

AND2x2_ASAP7_75t_L g7491 ( 
.A(n_7403),
.B(n_6238),
.Y(n_7491)
);

INVx2_ASAP7_75t_L g7492 ( 
.A(n_6669),
.Y(n_7492)
);

OAI22xp33_ASAP7_75t_L g7493 ( 
.A1(n_6480),
.A2(n_6251),
.B1(n_6230),
.B2(n_6013),
.Y(n_7493)
);

AOI22xp33_ASAP7_75t_L g7494 ( 
.A1(n_7218),
.A2(n_5946),
.B1(n_5911),
.B2(n_6124),
.Y(n_7494)
);

AO21x2_ASAP7_75t_L g7495 ( 
.A1(n_6862),
.A2(n_5784),
.B(n_5779),
.Y(n_7495)
);

INVx2_ASAP7_75t_L g7496 ( 
.A(n_6894),
.Y(n_7496)
);

AOI22xp33_ASAP7_75t_L g7497 ( 
.A1(n_7218),
.A2(n_5946),
.B1(n_5911),
.B2(n_6124),
.Y(n_7497)
);

OAI21x1_ASAP7_75t_L g7498 ( 
.A1(n_6986),
.A2(n_5956),
.B(n_5949),
.Y(n_7498)
);

HB1xp67_ASAP7_75t_L g7499 ( 
.A(n_6489),
.Y(n_7499)
);

INVx1_ASAP7_75t_L g7500 ( 
.A(n_6485),
.Y(n_7500)
);

INVx2_ASAP7_75t_L g7501 ( 
.A(n_6894),
.Y(n_7501)
);

AOI22xp33_ASAP7_75t_L g7502 ( 
.A1(n_6451),
.A2(n_5946),
.B1(n_5911),
.B2(n_5677),
.Y(n_7502)
);

AOI22xp5_ASAP7_75t_L g7503 ( 
.A1(n_6536),
.A2(n_5714),
.B1(n_5688),
.B2(n_5627),
.Y(n_7503)
);

INVx1_ASAP7_75t_SL g7504 ( 
.A(n_6991),
.Y(n_7504)
);

NOR2x1_ASAP7_75t_R g7505 ( 
.A(n_7306),
.B(n_6293),
.Y(n_7505)
);

AOI22xp33_ASAP7_75t_SL g7506 ( 
.A1(n_6746),
.A2(n_5573),
.B1(n_5677),
.B2(n_5861),
.Y(n_7506)
);

INVx2_ASAP7_75t_L g7507 ( 
.A(n_6894),
.Y(n_7507)
);

OR2x2_ASAP7_75t_L g7508 ( 
.A(n_6585),
.B(n_5784),
.Y(n_7508)
);

BUFx2_ASAP7_75t_L g7509 ( 
.A(n_6521),
.Y(n_7509)
);

INVx3_ASAP7_75t_L g7510 ( 
.A(n_6855),
.Y(n_7510)
);

OAI22xp5_ASAP7_75t_L g7511 ( 
.A1(n_6549),
.A2(n_5916),
.B1(n_5895),
.B2(n_6320),
.Y(n_7511)
);

INVx2_ASAP7_75t_L g7512 ( 
.A(n_6894),
.Y(n_7512)
);

INVx1_ASAP7_75t_L g7513 ( 
.A(n_6495),
.Y(n_7513)
);

OAI21x1_ASAP7_75t_L g7514 ( 
.A1(n_6986),
.A2(n_5956),
.B(n_5949),
.Y(n_7514)
);

BUFx4f_ASAP7_75t_SL g7515 ( 
.A(n_6942),
.Y(n_7515)
);

INVx2_ASAP7_75t_L g7516 ( 
.A(n_7279),
.Y(n_7516)
);

AOI22xp33_ASAP7_75t_L g7517 ( 
.A1(n_6611),
.A2(n_5677),
.B1(n_5573),
.B2(n_5719),
.Y(n_7517)
);

INVx1_ASAP7_75t_L g7518 ( 
.A(n_6495),
.Y(n_7518)
);

AOI22xp33_ASAP7_75t_L g7519 ( 
.A1(n_6611),
.A2(n_5677),
.B1(n_5573),
.B2(n_5719),
.Y(n_7519)
);

BUFx6f_ASAP7_75t_SL g7520 ( 
.A(n_6574),
.Y(n_7520)
);

BUFx12f_ASAP7_75t_L g7521 ( 
.A(n_6799),
.Y(n_7521)
);

HB1xp67_ASAP7_75t_L g7522 ( 
.A(n_6489),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_6498),
.Y(n_7523)
);

AOI22xp33_ASAP7_75t_L g7524 ( 
.A1(n_6608),
.A2(n_5677),
.B1(n_5573),
.B2(n_5719),
.Y(n_7524)
);

BUFx2_ASAP7_75t_L g7525 ( 
.A(n_6521),
.Y(n_7525)
);

INVx3_ASAP7_75t_L g7526 ( 
.A(n_6855),
.Y(n_7526)
);

INVx2_ASAP7_75t_L g7527 ( 
.A(n_7279),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_6498),
.Y(n_7528)
);

BUFx6f_ASAP7_75t_L g7529 ( 
.A(n_6574),
.Y(n_7529)
);

INVx1_ASAP7_75t_L g7530 ( 
.A(n_6512),
.Y(n_7530)
);

INVx2_ASAP7_75t_L g7531 ( 
.A(n_7279),
.Y(n_7531)
);

INVx3_ASAP7_75t_L g7532 ( 
.A(n_7178),
.Y(n_7532)
);

HB1xp67_ASAP7_75t_L g7533 ( 
.A(n_6494),
.Y(n_7533)
);

BUFx6f_ASAP7_75t_L g7534 ( 
.A(n_6574),
.Y(n_7534)
);

INVx2_ASAP7_75t_SL g7535 ( 
.A(n_7376),
.Y(n_7535)
);

AOI22xp33_ASAP7_75t_L g7536 ( 
.A1(n_6608),
.A2(n_5677),
.B1(n_5573),
.B2(n_5719),
.Y(n_7536)
);

INVx2_ASAP7_75t_L g7537 ( 
.A(n_7279),
.Y(n_7537)
);

AOI21x1_ASAP7_75t_L g7538 ( 
.A1(n_7324),
.A2(n_6131),
.B(n_6112),
.Y(n_7538)
);

INVx1_ASAP7_75t_L g7539 ( 
.A(n_6512),
.Y(n_7539)
);

HB1xp67_ASAP7_75t_L g7540 ( 
.A(n_6494),
.Y(n_7540)
);

INVx1_ASAP7_75t_SL g7541 ( 
.A(n_6942),
.Y(n_7541)
);

OR2x2_ASAP7_75t_L g7542 ( 
.A(n_6585),
.B(n_6123),
.Y(n_7542)
);

BUFx2_ASAP7_75t_L g7543 ( 
.A(n_6521),
.Y(n_7543)
);

BUFx4f_ASAP7_75t_SL g7544 ( 
.A(n_6891),
.Y(n_7544)
);

BUFx2_ASAP7_75t_SL g7545 ( 
.A(n_7306),
.Y(n_7545)
);

INVx2_ASAP7_75t_L g7546 ( 
.A(n_7296),
.Y(n_7546)
);

INVx1_ASAP7_75t_L g7547 ( 
.A(n_6517),
.Y(n_7547)
);

INVx2_ASAP7_75t_L g7548 ( 
.A(n_7296),
.Y(n_7548)
);

INVx3_ASAP7_75t_L g7549 ( 
.A(n_7178),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_6517),
.Y(n_7550)
);

AOI22xp33_ASAP7_75t_L g7551 ( 
.A1(n_6595),
.A2(n_5677),
.B1(n_5798),
.B2(n_5719),
.Y(n_7551)
);

CKINVDCx20_ASAP7_75t_R g7552 ( 
.A(n_6851),
.Y(n_7552)
);

INVx2_ASAP7_75t_SL g7553 ( 
.A(n_6519),
.Y(n_7553)
);

AOI22xp33_ASAP7_75t_L g7554 ( 
.A1(n_6595),
.A2(n_5677),
.B1(n_5798),
.B2(n_5719),
.Y(n_7554)
);

INVx2_ASAP7_75t_L g7555 ( 
.A(n_7296),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_6518),
.Y(n_7556)
);

AOI21x1_ASAP7_75t_L g7557 ( 
.A1(n_7324),
.A2(n_6151),
.B(n_6131),
.Y(n_7557)
);

INVx2_ASAP7_75t_L g7558 ( 
.A(n_7296),
.Y(n_7558)
);

INVx1_ASAP7_75t_SL g7559 ( 
.A(n_6851),
.Y(n_7559)
);

BUFx2_ASAP7_75t_L g7560 ( 
.A(n_6521),
.Y(n_7560)
);

INVx1_ASAP7_75t_L g7561 ( 
.A(n_6518),
.Y(n_7561)
);

INVx2_ASAP7_75t_L g7562 ( 
.A(n_7296),
.Y(n_7562)
);

AND2x2_ASAP7_75t_L g7563 ( 
.A(n_7403),
.B(n_7295),
.Y(n_7563)
);

OR2x2_ASAP7_75t_L g7564 ( 
.A(n_6585),
.B(n_6123),
.Y(n_7564)
);

INVx1_ASAP7_75t_L g7565 ( 
.A(n_6548),
.Y(n_7565)
);

OA21x2_ASAP7_75t_L g7566 ( 
.A1(n_6702),
.A2(n_6445),
.B(n_6444),
.Y(n_7566)
);

INVx2_ASAP7_75t_L g7567 ( 
.A(n_7357),
.Y(n_7567)
);

INVx3_ASAP7_75t_L g7568 ( 
.A(n_7178),
.Y(n_7568)
);

OAI22xp5_ASAP7_75t_L g7569 ( 
.A1(n_6549),
.A2(n_5916),
.B1(n_5895),
.B2(n_6320),
.Y(n_7569)
);

CKINVDCx20_ASAP7_75t_R g7570 ( 
.A(n_6879),
.Y(n_7570)
);

BUFx2_ASAP7_75t_R g7571 ( 
.A(n_6926),
.Y(n_7571)
);

INVx1_ASAP7_75t_L g7572 ( 
.A(n_6548),
.Y(n_7572)
);

AND2x2_ASAP7_75t_L g7573 ( 
.A(n_7295),
.B(n_6892),
.Y(n_7573)
);

INVx1_ASAP7_75t_L g7574 ( 
.A(n_6554),
.Y(n_7574)
);

INVxp67_ASAP7_75t_L g7575 ( 
.A(n_7098),
.Y(n_7575)
);

AOI22xp33_ASAP7_75t_L g7576 ( 
.A1(n_6635),
.A2(n_5677),
.B1(n_5798),
.B2(n_5719),
.Y(n_7576)
);

INVxp67_ASAP7_75t_L g7577 ( 
.A(n_7098),
.Y(n_7577)
);

AND2x4_ASAP7_75t_L g7578 ( 
.A(n_6506),
.B(n_6167),
.Y(n_7578)
);

CKINVDCx5p33_ASAP7_75t_R g7579 ( 
.A(n_6879),
.Y(n_7579)
);

INVx1_ASAP7_75t_L g7580 ( 
.A(n_6554),
.Y(n_7580)
);

OR2x2_ASAP7_75t_L g7581 ( 
.A(n_7099),
.B(n_5987),
.Y(n_7581)
);

OAI22xp5_ASAP7_75t_L g7582 ( 
.A1(n_6586),
.A2(n_5916),
.B1(n_6011),
.B2(n_5638),
.Y(n_7582)
);

INVx1_ASAP7_75t_L g7583 ( 
.A(n_6555),
.Y(n_7583)
);

INVx3_ASAP7_75t_L g7584 ( 
.A(n_7178),
.Y(n_7584)
);

INVx2_ASAP7_75t_SL g7585 ( 
.A(n_6519),
.Y(n_7585)
);

HB1xp67_ASAP7_75t_L g7586 ( 
.A(n_6542),
.Y(n_7586)
);

INVx2_ASAP7_75t_L g7587 ( 
.A(n_6894),
.Y(n_7587)
);

INVx6_ASAP7_75t_L g7588 ( 
.A(n_6774),
.Y(n_7588)
);

INVx1_ASAP7_75t_L g7589 ( 
.A(n_6555),
.Y(n_7589)
);

INVx1_ASAP7_75t_L g7590 ( 
.A(n_6560),
.Y(n_7590)
);

INVx2_ASAP7_75t_L g7591 ( 
.A(n_6743),
.Y(n_7591)
);

NAND2xp5_ASAP7_75t_L g7592 ( 
.A(n_7077),
.B(n_6214),
.Y(n_7592)
);

INVx1_ASAP7_75t_L g7593 ( 
.A(n_6560),
.Y(n_7593)
);

INVx2_ASAP7_75t_L g7594 ( 
.A(n_7357),
.Y(n_7594)
);

HB1xp67_ASAP7_75t_L g7595 ( 
.A(n_6542),
.Y(n_7595)
);

AND2x4_ASAP7_75t_L g7596 ( 
.A(n_6506),
.B(n_6167),
.Y(n_7596)
);

AND2x2_ASAP7_75t_L g7597 ( 
.A(n_6892),
.B(n_6238),
.Y(n_7597)
);

INVx1_ASAP7_75t_L g7598 ( 
.A(n_6575),
.Y(n_7598)
);

AOI22xp33_ASAP7_75t_L g7599 ( 
.A1(n_6635),
.A2(n_5677),
.B1(n_5863),
.B2(n_5798),
.Y(n_7599)
);

BUFx3_ASAP7_75t_L g7600 ( 
.A(n_7306),
.Y(n_7600)
);

INVx2_ASAP7_75t_L g7601 ( 
.A(n_7357),
.Y(n_7601)
);

INVx1_ASAP7_75t_L g7602 ( 
.A(n_6575),
.Y(n_7602)
);

INVx1_ASAP7_75t_L g7603 ( 
.A(n_6576),
.Y(n_7603)
);

INVx2_ASAP7_75t_L g7604 ( 
.A(n_7357),
.Y(n_7604)
);

NAND2x1p5_ASAP7_75t_L g7605 ( 
.A(n_7198),
.B(n_5880),
.Y(n_7605)
);

AND2x4_ASAP7_75t_L g7606 ( 
.A(n_6506),
.B(n_6167),
.Y(n_7606)
);

BUFx4f_ASAP7_75t_L g7607 ( 
.A(n_7382),
.Y(n_7607)
);

OAI22xp5_ASAP7_75t_L g7608 ( 
.A1(n_6586),
.A2(n_5916),
.B1(n_6011),
.B2(n_5638),
.Y(n_7608)
);

NAND2xp5_ASAP7_75t_L g7609 ( 
.A(n_6645),
.B(n_6214),
.Y(n_7609)
);

INVx1_ASAP7_75t_L g7610 ( 
.A(n_6576),
.Y(n_7610)
);

INVx1_ASAP7_75t_L g7611 ( 
.A(n_6590),
.Y(n_7611)
);

NAND2x1p5_ASAP7_75t_L g7612 ( 
.A(n_7198),
.B(n_5880),
.Y(n_7612)
);

INVx1_ASAP7_75t_L g7613 ( 
.A(n_6590),
.Y(n_7613)
);

INVx2_ASAP7_75t_L g7614 ( 
.A(n_7357),
.Y(n_7614)
);

INVx1_ASAP7_75t_L g7615 ( 
.A(n_6597),
.Y(n_7615)
);

INVx2_ASAP7_75t_SL g7616 ( 
.A(n_6519),
.Y(n_7616)
);

INVx1_ASAP7_75t_L g7617 ( 
.A(n_6597),
.Y(n_7617)
);

AO21x1_ASAP7_75t_L g7618 ( 
.A1(n_7135),
.A2(n_5800),
.B(n_5799),
.Y(n_7618)
);

CKINVDCx20_ASAP7_75t_R g7619 ( 
.A(n_7224),
.Y(n_7619)
);

AND2x2_ASAP7_75t_L g7620 ( 
.A(n_6892),
.B(n_6907),
.Y(n_7620)
);

OAI22xp5_ASAP7_75t_L g7621 ( 
.A1(n_6586),
.A2(n_6011),
.B1(n_5638),
.B2(n_5992),
.Y(n_7621)
);

INVx2_ASAP7_75t_L g7622 ( 
.A(n_7367),
.Y(n_7622)
);

INVx3_ASAP7_75t_L g7623 ( 
.A(n_7178),
.Y(n_7623)
);

INVx2_ASAP7_75t_L g7624 ( 
.A(n_7367),
.Y(n_7624)
);

HB1xp67_ASAP7_75t_L g7625 ( 
.A(n_6553),
.Y(n_7625)
);

AND2x4_ASAP7_75t_L g7626 ( 
.A(n_6506),
.B(n_6167),
.Y(n_7626)
);

AND2x4_ASAP7_75t_L g7627 ( 
.A(n_6506),
.B(n_6193),
.Y(n_7627)
);

OAI22xp5_ASAP7_75t_L g7628 ( 
.A1(n_6461),
.A2(n_6011),
.B1(n_5638),
.B2(n_5992),
.Y(n_7628)
);

AOI22xp33_ASAP7_75t_SL g7629 ( 
.A1(n_6716),
.A2(n_5677),
.B1(n_5861),
.B2(n_6193),
.Y(n_7629)
);

AO21x1_ASAP7_75t_SL g7630 ( 
.A1(n_6551),
.A2(n_6092),
.B(n_6078),
.Y(n_7630)
);

HB1xp67_ASAP7_75t_L g7631 ( 
.A(n_6553),
.Y(n_7631)
);

AOI21x1_ASAP7_75t_L g7632 ( 
.A1(n_6516),
.A2(n_6151),
.B(n_6131),
.Y(n_7632)
);

AND2x4_ASAP7_75t_L g7633 ( 
.A(n_6930),
.B(n_6193),
.Y(n_7633)
);

OA21x2_ASAP7_75t_L g7634 ( 
.A1(n_6702),
.A2(n_6054),
.B(n_6045),
.Y(n_7634)
);

INVx3_ASAP7_75t_L g7635 ( 
.A(n_7022),
.Y(n_7635)
);

OAI21x1_ASAP7_75t_L g7636 ( 
.A1(n_6476),
.A2(n_5983),
.B(n_5956),
.Y(n_7636)
);

AOI22xp33_ASAP7_75t_L g7637 ( 
.A1(n_6551),
.A2(n_5863),
.B1(n_5981),
.B2(n_5798),
.Y(n_7637)
);

INVx2_ASAP7_75t_L g7638 ( 
.A(n_7367),
.Y(n_7638)
);

INVx1_ASAP7_75t_L g7639 ( 
.A(n_6612),
.Y(n_7639)
);

INVx3_ASAP7_75t_L g7640 ( 
.A(n_7022),
.Y(n_7640)
);

AO21x1_ASAP7_75t_SL g7641 ( 
.A1(n_6742),
.A2(n_6108),
.B(n_6096),
.Y(n_7641)
);

OAI22xp5_ASAP7_75t_L g7642 ( 
.A1(n_6461),
.A2(n_6234),
.B1(n_6341),
.B2(n_5876),
.Y(n_7642)
);

HB1xp67_ASAP7_75t_L g7643 ( 
.A(n_6582),
.Y(n_7643)
);

INVx3_ASAP7_75t_L g7644 ( 
.A(n_7022),
.Y(n_7644)
);

BUFx2_ASAP7_75t_L g7645 ( 
.A(n_6521),
.Y(n_7645)
);

OAI22xp5_ASAP7_75t_L g7646 ( 
.A1(n_6492),
.A2(n_6234),
.B1(n_6341),
.B2(n_5876),
.Y(n_7646)
);

INVx8_ASAP7_75t_L g7647 ( 
.A(n_6824),
.Y(n_7647)
);

AOI22xp33_ASAP7_75t_SL g7648 ( 
.A1(n_6716),
.A2(n_5861),
.B1(n_6225),
.B2(n_6193),
.Y(n_7648)
);

INVx1_ASAP7_75t_L g7649 ( 
.A(n_6612),
.Y(n_7649)
);

AOI22xp33_ASAP7_75t_L g7650 ( 
.A1(n_6862),
.A2(n_5863),
.B1(n_5981),
.B2(n_5798),
.Y(n_7650)
);

AOI22xp33_ASAP7_75t_L g7651 ( 
.A1(n_6862),
.A2(n_6736),
.B1(n_6727),
.B2(n_6909),
.Y(n_7651)
);

AND2x2_ASAP7_75t_L g7652 ( 
.A(n_6907),
.B(n_6238),
.Y(n_7652)
);

INVx1_ASAP7_75t_L g7653 ( 
.A(n_6615),
.Y(n_7653)
);

INVx2_ASAP7_75t_L g7654 ( 
.A(n_7367),
.Y(n_7654)
);

INVx3_ASAP7_75t_L g7655 ( 
.A(n_7022),
.Y(n_7655)
);

INVx2_ASAP7_75t_L g7656 ( 
.A(n_7367),
.Y(n_7656)
);

BUFx2_ASAP7_75t_L g7657 ( 
.A(n_6521),
.Y(n_7657)
);

NAND2xp5_ASAP7_75t_L g7658 ( 
.A(n_6645),
.B(n_6330),
.Y(n_7658)
);

INVx1_ASAP7_75t_L g7659 ( 
.A(n_6615),
.Y(n_7659)
);

INVx1_ASAP7_75t_L g7660 ( 
.A(n_6621),
.Y(n_7660)
);

AOI22xp33_ASAP7_75t_L g7661 ( 
.A1(n_6862),
.A2(n_5863),
.B1(n_5981),
.B2(n_5798),
.Y(n_7661)
);

INVx1_ASAP7_75t_SL g7662 ( 
.A(n_7224),
.Y(n_7662)
);

AOI22xp33_ASAP7_75t_L g7663 ( 
.A1(n_6727),
.A2(n_5981),
.B1(n_6192),
.B2(n_5863),
.Y(n_7663)
);

INVx2_ASAP7_75t_L g7664 ( 
.A(n_7400),
.Y(n_7664)
);

HB1xp67_ASAP7_75t_L g7665 ( 
.A(n_6582),
.Y(n_7665)
);

HB1xp67_ASAP7_75t_L g7666 ( 
.A(n_6592),
.Y(n_7666)
);

INVx1_ASAP7_75t_L g7667 ( 
.A(n_6621),
.Y(n_7667)
);

BUFx3_ASAP7_75t_L g7668 ( 
.A(n_6799),
.Y(n_7668)
);

OAI21x1_ASAP7_75t_L g7669 ( 
.A1(n_6476),
.A2(n_5983),
.B(n_5956),
.Y(n_7669)
);

BUFx4f_ASAP7_75t_SL g7670 ( 
.A(n_6891),
.Y(n_7670)
);

INVx1_ASAP7_75t_L g7671 ( 
.A(n_6624),
.Y(n_7671)
);

AND2x2_ASAP7_75t_L g7672 ( 
.A(n_6907),
.B(n_6268),
.Y(n_7672)
);

BUFx2_ASAP7_75t_L g7673 ( 
.A(n_6521),
.Y(n_7673)
);

NAND2x1p5_ASAP7_75t_L g7674 ( 
.A(n_7198),
.B(n_5880),
.Y(n_7674)
);

INVx1_ASAP7_75t_L g7675 ( 
.A(n_6624),
.Y(n_7675)
);

OA21x2_ASAP7_75t_L g7676 ( 
.A1(n_6444),
.A2(n_6164),
.B(n_6054),
.Y(n_7676)
);

INVx1_ASAP7_75t_L g7677 ( 
.A(n_6633),
.Y(n_7677)
);

AO21x1_ASAP7_75t_SL g7678 ( 
.A1(n_6742),
.A2(n_6108),
.B(n_6096),
.Y(n_7678)
);

INVx2_ASAP7_75t_L g7679 ( 
.A(n_7400),
.Y(n_7679)
);

AOI22xp5_ASAP7_75t_L g7680 ( 
.A1(n_6505),
.A2(n_5674),
.B1(n_5962),
.B2(n_5988),
.Y(n_7680)
);

OAI22xp5_ASAP7_75t_L g7681 ( 
.A1(n_6492),
.A2(n_5876),
.B1(n_5859),
.B2(n_6285),
.Y(n_7681)
);

BUFx3_ASAP7_75t_L g7682 ( 
.A(n_6799),
.Y(n_7682)
);

INVx1_ASAP7_75t_L g7683 ( 
.A(n_6633),
.Y(n_7683)
);

BUFx8_ASAP7_75t_SL g7684 ( 
.A(n_6891),
.Y(n_7684)
);

BUFx6f_ASAP7_75t_L g7685 ( 
.A(n_6622),
.Y(n_7685)
);

AOI22xp33_ASAP7_75t_SL g7686 ( 
.A1(n_6915),
.A2(n_6235),
.B1(n_6270),
.B2(n_6225),
.Y(n_7686)
);

OR2x2_ASAP7_75t_L g7687 ( 
.A(n_7099),
.B(n_6533),
.Y(n_7687)
);

OAI22xp5_ASAP7_75t_L g7688 ( 
.A1(n_6909),
.A2(n_5859),
.B1(n_6424),
.B2(n_6285),
.Y(n_7688)
);

AO21x1_ASAP7_75t_L g7689 ( 
.A1(n_7135),
.A2(n_5800),
.B(n_5799),
.Y(n_7689)
);

INVx2_ASAP7_75t_L g7690 ( 
.A(n_7400),
.Y(n_7690)
);

INVx2_ASAP7_75t_L g7691 ( 
.A(n_7400),
.Y(n_7691)
);

INVx2_ASAP7_75t_L g7692 ( 
.A(n_7400),
.Y(n_7692)
);

OR2x6_ASAP7_75t_L g7693 ( 
.A(n_6606),
.B(n_5863),
.Y(n_7693)
);

NOR2xp33_ASAP7_75t_L g7694 ( 
.A(n_7215),
.B(n_5823),
.Y(n_7694)
);

INVx2_ASAP7_75t_L g7695 ( 
.A(n_7406),
.Y(n_7695)
);

CKINVDCx20_ASAP7_75t_R g7696 ( 
.A(n_7017),
.Y(n_7696)
);

INVx8_ASAP7_75t_L g7697 ( 
.A(n_6824),
.Y(n_7697)
);

OAI22xp5_ASAP7_75t_L g7698 ( 
.A1(n_6484),
.A2(n_5859),
.B1(n_6424),
.B2(n_6285),
.Y(n_7698)
);

OA21x2_ASAP7_75t_L g7699 ( 
.A1(n_6444),
.A2(n_6321),
.B(n_6164),
.Y(n_7699)
);

OR2x6_ASAP7_75t_L g7700 ( 
.A(n_6606),
.B(n_5981),
.Y(n_7700)
);

INVx2_ASAP7_75t_L g7701 ( 
.A(n_7406),
.Y(n_7701)
);

BUFx4f_ASAP7_75t_L g7702 ( 
.A(n_7382),
.Y(n_7702)
);

AOI22xp33_ASAP7_75t_L g7703 ( 
.A1(n_6736),
.A2(n_5981),
.B1(n_6192),
.B2(n_5863),
.Y(n_7703)
);

AOI22xp5_ASAP7_75t_L g7704 ( 
.A1(n_6505),
.A2(n_5674),
.B1(n_5962),
.B2(n_5988),
.Y(n_7704)
);

INVx1_ASAP7_75t_L g7705 ( 
.A(n_6636),
.Y(n_7705)
);

INVx2_ASAP7_75t_L g7706 ( 
.A(n_7406),
.Y(n_7706)
);

INVx2_ASAP7_75t_L g7707 ( 
.A(n_7406),
.Y(n_7707)
);

INVx2_ASAP7_75t_L g7708 ( 
.A(n_7406),
.Y(n_7708)
);

AND2x4_ASAP7_75t_L g7709 ( 
.A(n_6930),
.B(n_6225),
.Y(n_7709)
);

NAND2xp5_ASAP7_75t_L g7710 ( 
.A(n_6655),
.B(n_6330),
.Y(n_7710)
);

BUFx2_ASAP7_75t_L g7711 ( 
.A(n_7346),
.Y(n_7711)
);

AND2x2_ASAP7_75t_L g7712 ( 
.A(n_6914),
.B(n_6268),
.Y(n_7712)
);

AO21x1_ASAP7_75t_L g7713 ( 
.A1(n_6915),
.A2(n_5808),
.B(n_5807),
.Y(n_7713)
);

INVx1_ASAP7_75t_L g7714 ( 
.A(n_6636),
.Y(n_7714)
);

AOI22xp33_ASAP7_75t_L g7715 ( 
.A1(n_6787),
.A2(n_6192),
.B1(n_5981),
.B2(n_6242),
.Y(n_7715)
);

INVx1_ASAP7_75t_L g7716 ( 
.A(n_6643),
.Y(n_7716)
);

AOI22xp33_ASAP7_75t_L g7717 ( 
.A1(n_6787),
.A2(n_6192),
.B1(n_6319),
.B2(n_6242),
.Y(n_7717)
);

INVx2_ASAP7_75t_L g7718 ( 
.A(n_6743),
.Y(n_7718)
);

INVx2_ASAP7_75t_L g7719 ( 
.A(n_6743),
.Y(n_7719)
);

OAI21x1_ASAP7_75t_L g7720 ( 
.A1(n_6899),
.A2(n_5989),
.B(n_5983),
.Y(n_7720)
);

CKINVDCx5p33_ASAP7_75t_R g7721 ( 
.A(n_6887),
.Y(n_7721)
);

INVx1_ASAP7_75t_L g7722 ( 
.A(n_6643),
.Y(n_7722)
);

AOI22xp33_ASAP7_75t_L g7723 ( 
.A1(n_6563),
.A2(n_6192),
.B1(n_6319),
.B2(n_6242),
.Y(n_7723)
);

HB1xp67_ASAP7_75t_L g7724 ( 
.A(n_6592),
.Y(n_7724)
);

AOI22xp33_ASAP7_75t_L g7725 ( 
.A1(n_6563),
.A2(n_6956),
.B1(n_7018),
.B2(n_6699),
.Y(n_7725)
);

NAND2xp5_ASAP7_75t_L g7726 ( 
.A(n_6655),
.B(n_5965),
.Y(n_7726)
);

AOI22xp33_ASAP7_75t_L g7727 ( 
.A1(n_6956),
.A2(n_6192),
.B1(n_6319),
.B2(n_6242),
.Y(n_7727)
);

INVx1_ASAP7_75t_L g7728 ( 
.A(n_6658),
.Y(n_7728)
);

INVx2_ASAP7_75t_L g7729 ( 
.A(n_6743),
.Y(n_7729)
);

HB1xp67_ASAP7_75t_L g7730 ( 
.A(n_6674),
.Y(n_7730)
);

OAI22xp5_ASAP7_75t_L g7731 ( 
.A1(n_6484),
.A2(n_6424),
.B1(n_5957),
.B2(n_5736),
.Y(n_7731)
);

AND2x2_ASAP7_75t_L g7732 ( 
.A(n_6914),
.B(n_6268),
.Y(n_7732)
);

BUFx2_ASAP7_75t_R g7733 ( 
.A(n_7028),
.Y(n_7733)
);

INVx1_ASAP7_75t_L g7734 ( 
.A(n_6658),
.Y(n_7734)
);

OAI22xp33_ASAP7_75t_L g7735 ( 
.A1(n_6566),
.A2(n_6543),
.B1(n_6710),
.B2(n_6533),
.Y(n_7735)
);

OAI21x1_ASAP7_75t_SL g7736 ( 
.A1(n_6801),
.A2(n_6130),
.B(n_6122),
.Y(n_7736)
);

INVx1_ASAP7_75t_L g7737 ( 
.A(n_6677),
.Y(n_7737)
);

INVx11_ASAP7_75t_L g7738 ( 
.A(n_6887),
.Y(n_7738)
);

INVx2_ASAP7_75t_L g7739 ( 
.A(n_6743),
.Y(n_7739)
);

CKINVDCx11_ASAP7_75t_R g7740 ( 
.A(n_6967),
.Y(n_7740)
);

INVx3_ASAP7_75t_L g7741 ( 
.A(n_7022),
.Y(n_7741)
);

CKINVDCx9p33_ASAP7_75t_R g7742 ( 
.A(n_7215),
.Y(n_7742)
);

NAND2x1p5_ASAP7_75t_L g7743 ( 
.A(n_7198),
.B(n_5880),
.Y(n_7743)
);

INVx1_ASAP7_75t_L g7744 ( 
.A(n_6677),
.Y(n_7744)
);

INVx1_ASAP7_75t_L g7745 ( 
.A(n_6681),
.Y(n_7745)
);

INVx1_ASAP7_75t_L g7746 ( 
.A(n_6681),
.Y(n_7746)
);

INVx2_ASAP7_75t_L g7747 ( 
.A(n_7059),
.Y(n_7747)
);

BUFx3_ASAP7_75t_L g7748 ( 
.A(n_6887),
.Y(n_7748)
);

NAND2x1p5_ASAP7_75t_L g7749 ( 
.A(n_7198),
.B(n_5882),
.Y(n_7749)
);

AOI22xp33_ASAP7_75t_L g7750 ( 
.A1(n_7018),
.A2(n_6192),
.B1(n_6319),
.B2(n_6242),
.Y(n_7750)
);

AOI22xp5_ASAP7_75t_SL g7751 ( 
.A1(n_6587),
.A2(n_6152),
.B1(n_6169),
.B2(n_6098),
.Y(n_7751)
);

OR2x2_ASAP7_75t_L g7752 ( 
.A(n_7099),
.B(n_5987),
.Y(n_7752)
);

INVx6_ASAP7_75t_L g7753 ( 
.A(n_6774),
.Y(n_7753)
);

INVx2_ASAP7_75t_L g7754 ( 
.A(n_7059),
.Y(n_7754)
);

INVx1_ASAP7_75t_L g7755 ( 
.A(n_6689),
.Y(n_7755)
);

INVx2_ASAP7_75t_L g7756 ( 
.A(n_7059),
.Y(n_7756)
);

AOI22xp33_ASAP7_75t_SL g7757 ( 
.A1(n_7014),
.A2(n_6235),
.B1(n_6270),
.B2(n_6225),
.Y(n_7757)
);

INVx3_ASAP7_75t_L g7758 ( 
.A(n_7102),
.Y(n_7758)
);

NAND2x1p5_ASAP7_75t_L g7759 ( 
.A(n_7198),
.B(n_7008),
.Y(n_7759)
);

INVx1_ASAP7_75t_L g7760 ( 
.A(n_6689),
.Y(n_7760)
);

AND2x4_ASAP7_75t_L g7761 ( 
.A(n_6930),
.B(n_6235),
.Y(n_7761)
);

BUFx6f_ASAP7_75t_L g7762 ( 
.A(n_6622),
.Y(n_7762)
);

INVx1_ASAP7_75t_L g7763 ( 
.A(n_6706),
.Y(n_7763)
);

INVx1_ASAP7_75t_L g7764 ( 
.A(n_6706),
.Y(n_7764)
);

BUFx4f_ASAP7_75t_SL g7765 ( 
.A(n_6967),
.Y(n_7765)
);

INVx3_ASAP7_75t_L g7766 ( 
.A(n_7102),
.Y(n_7766)
);

INVx1_ASAP7_75t_L g7767 ( 
.A(n_6707),
.Y(n_7767)
);

OAI22xp33_ASAP7_75t_L g7768 ( 
.A1(n_6566),
.A2(n_6230),
.B1(n_6013),
.B2(n_5750),
.Y(n_7768)
);

CKINVDCx5p33_ASAP7_75t_R g7769 ( 
.A(n_6967),
.Y(n_7769)
);

AND2x4_ASAP7_75t_L g7770 ( 
.A(n_6930),
.B(n_6235),
.Y(n_7770)
);

BUFx4f_ASAP7_75t_SL g7771 ( 
.A(n_7382),
.Y(n_7771)
);

AND2x2_ASAP7_75t_L g7772 ( 
.A(n_6914),
.B(n_6268),
.Y(n_7772)
);

INVx2_ASAP7_75t_L g7773 ( 
.A(n_7059),
.Y(n_7773)
);

BUFx3_ASAP7_75t_L g7774 ( 
.A(n_6680),
.Y(n_7774)
);

INVx1_ASAP7_75t_L g7775 ( 
.A(n_6707),
.Y(n_7775)
);

INVx1_ASAP7_75t_L g7776 ( 
.A(n_6712),
.Y(n_7776)
);

INVx2_ASAP7_75t_L g7777 ( 
.A(n_7059),
.Y(n_7777)
);

AOI22xp33_ASAP7_75t_L g7778 ( 
.A1(n_7018),
.A2(n_6319),
.B1(n_6242),
.B2(n_5559),
.Y(n_7778)
);

INVx1_ASAP7_75t_L g7779 ( 
.A(n_6712),
.Y(n_7779)
);

INVx1_ASAP7_75t_L g7780 ( 
.A(n_6724),
.Y(n_7780)
);

BUFx2_ASAP7_75t_L g7781 ( 
.A(n_7346),
.Y(n_7781)
);

BUFx2_ASAP7_75t_L g7782 ( 
.A(n_6680),
.Y(n_7782)
);

OAI21x1_ASAP7_75t_L g7783 ( 
.A1(n_6899),
.A2(n_5989),
.B(n_5983),
.Y(n_7783)
);

AND2x4_ASAP7_75t_L g7784 ( 
.A(n_6930),
.B(n_6270),
.Y(n_7784)
);

BUFx6f_ASAP7_75t_L g7785 ( 
.A(n_6622),
.Y(n_7785)
);

INVx3_ASAP7_75t_L g7786 ( 
.A(n_7102),
.Y(n_7786)
);

INVx1_ASAP7_75t_L g7787 ( 
.A(n_6724),
.Y(n_7787)
);

HB1xp67_ASAP7_75t_L g7788 ( 
.A(n_6674),
.Y(n_7788)
);

INVx2_ASAP7_75t_SL g7789 ( 
.A(n_6520),
.Y(n_7789)
);

AOI22xp33_ASAP7_75t_L g7790 ( 
.A1(n_7018),
.A2(n_6319),
.B1(n_6242),
.B2(n_5559),
.Y(n_7790)
);

HB1xp67_ASAP7_75t_L g7791 ( 
.A(n_6826),
.Y(n_7791)
);

INVx1_ASAP7_75t_SL g7792 ( 
.A(n_7017),
.Y(n_7792)
);

INVx2_ASAP7_75t_L g7793 ( 
.A(n_7065),
.Y(n_7793)
);

INVx1_ASAP7_75t_L g7794 ( 
.A(n_6739),
.Y(n_7794)
);

NOR2xp33_ASAP7_75t_L g7795 ( 
.A(n_7142),
.B(n_5907),
.Y(n_7795)
);

INVx1_ASAP7_75t_L g7796 ( 
.A(n_6739),
.Y(n_7796)
);

INVx2_ASAP7_75t_L g7797 ( 
.A(n_7065),
.Y(n_7797)
);

BUFx2_ASAP7_75t_R g7798 ( 
.A(n_7163),
.Y(n_7798)
);

NAND2x1p5_ASAP7_75t_L g7799 ( 
.A(n_7008),
.B(n_5882),
.Y(n_7799)
);

BUFx4f_ASAP7_75t_SL g7800 ( 
.A(n_6680),
.Y(n_7800)
);

OAI22xp5_ASAP7_75t_L g7801 ( 
.A1(n_6514),
.A2(n_6583),
.B1(n_6710),
.B2(n_7348),
.Y(n_7801)
);

NOR2xp33_ASAP7_75t_SL g7802 ( 
.A(n_6954),
.B(n_6001),
.Y(n_7802)
);

BUFx2_ASAP7_75t_L g7803 ( 
.A(n_6954),
.Y(n_7803)
);

INVx1_ASAP7_75t_L g7804 ( 
.A(n_6753),
.Y(n_7804)
);

AOI21x1_ASAP7_75t_L g7805 ( 
.A1(n_6516),
.A2(n_6177),
.B(n_6151),
.Y(n_7805)
);

INVx2_ASAP7_75t_L g7806 ( 
.A(n_7065),
.Y(n_7806)
);

AOI22xp33_ASAP7_75t_SL g7807 ( 
.A1(n_7014),
.A2(n_6276),
.B1(n_6297),
.B2(n_6270),
.Y(n_7807)
);

NAND2x1p5_ASAP7_75t_L g7808 ( 
.A(n_7008),
.B(n_5882),
.Y(n_7808)
);

INVx1_ASAP7_75t_L g7809 ( 
.A(n_6753),
.Y(n_7809)
);

OAI22xp33_ASAP7_75t_L g7810 ( 
.A1(n_6543),
.A2(n_5750),
.B1(n_6070),
.B2(n_6049),
.Y(n_7810)
);

INVx1_ASAP7_75t_L g7811 ( 
.A(n_6763),
.Y(n_7811)
);

INVx1_ASAP7_75t_L g7812 ( 
.A(n_6763),
.Y(n_7812)
);

HB1xp67_ASAP7_75t_L g7813 ( 
.A(n_6826),
.Y(n_7813)
);

AO21x1_ASAP7_75t_SL g7814 ( 
.A1(n_6857),
.A2(n_6115),
.B(n_6135),
.Y(n_7814)
);

OR2x2_ASAP7_75t_L g7815 ( 
.A(n_6649),
.B(n_6453),
.Y(n_7815)
);

INVx1_ASAP7_75t_L g7816 ( 
.A(n_6766),
.Y(n_7816)
);

INVx2_ASAP7_75t_L g7817 ( 
.A(n_7065),
.Y(n_7817)
);

INVx2_ASAP7_75t_L g7818 ( 
.A(n_7080),
.Y(n_7818)
);

OA21x2_ASAP7_75t_L g7819 ( 
.A1(n_6463),
.A2(n_6321),
.B(n_5603),
.Y(n_7819)
);

OAI21x1_ASAP7_75t_L g7820 ( 
.A1(n_6928),
.A2(n_5989),
.B(n_5983),
.Y(n_7820)
);

INVx1_ASAP7_75t_L g7821 ( 
.A(n_6766),
.Y(n_7821)
);

INVx1_ASAP7_75t_L g7822 ( 
.A(n_6779),
.Y(n_7822)
);

INVx1_ASAP7_75t_L g7823 ( 
.A(n_6779),
.Y(n_7823)
);

NAND2x1p5_ASAP7_75t_L g7824 ( 
.A(n_7008),
.B(n_7061),
.Y(n_7824)
);

AO21x1_ASAP7_75t_L g7825 ( 
.A1(n_7243),
.A2(n_6507),
.B(n_6469),
.Y(n_7825)
);

INVx1_ASAP7_75t_L g7826 ( 
.A(n_6782),
.Y(n_7826)
);

OAI21xp5_ASAP7_75t_L g7827 ( 
.A1(n_7243),
.A2(n_5547),
.B(n_5702),
.Y(n_7827)
);

INVx8_ASAP7_75t_L g7828 ( 
.A(n_6824),
.Y(n_7828)
);

BUFx3_ASAP7_75t_L g7829 ( 
.A(n_6774),
.Y(n_7829)
);

BUFx2_ASAP7_75t_R g7830 ( 
.A(n_7302),
.Y(n_7830)
);

OAI21xp33_ASAP7_75t_L g7831 ( 
.A1(n_7130),
.A2(n_6153),
.B(n_6148),
.Y(n_7831)
);

INVx1_ASAP7_75t_L g7832 ( 
.A(n_6782),
.Y(n_7832)
);

OAI21x1_ASAP7_75t_L g7833 ( 
.A1(n_6928),
.A2(n_5994),
.B(n_5989),
.Y(n_7833)
);

INVx2_ASAP7_75t_L g7834 ( 
.A(n_7080),
.Y(n_7834)
);

AND2x4_ASAP7_75t_L g7835 ( 
.A(n_6930),
.B(n_6276),
.Y(n_7835)
);

AOI22xp33_ASAP7_75t_SL g7836 ( 
.A1(n_7207),
.A2(n_6297),
.B1(n_6301),
.B2(n_6276),
.Y(n_7836)
);

INVx1_ASAP7_75t_L g7837 ( 
.A(n_6790),
.Y(n_7837)
);

BUFx2_ASAP7_75t_L g7838 ( 
.A(n_6632),
.Y(n_7838)
);

AND2x4_ASAP7_75t_L g7839 ( 
.A(n_6951),
.B(n_6276),
.Y(n_7839)
);

OA21x2_ASAP7_75t_L g7840 ( 
.A1(n_6463),
.A2(n_6194),
.B(n_6177),
.Y(n_7840)
);

NAND2xp5_ASAP7_75t_L g7841 ( 
.A(n_6695),
.B(n_5965),
.Y(n_7841)
);

INVx2_ASAP7_75t_L g7842 ( 
.A(n_7080),
.Y(n_7842)
);

NAND2xp5_ASAP7_75t_L g7843 ( 
.A(n_6695),
.B(n_6027),
.Y(n_7843)
);

AOI21x1_ASAP7_75t_L g7844 ( 
.A1(n_6456),
.A2(n_6194),
.B(n_6177),
.Y(n_7844)
);

INVx2_ASAP7_75t_SL g7845 ( 
.A(n_6520),
.Y(n_7845)
);

CKINVDCx11_ASAP7_75t_R g7846 ( 
.A(n_7179),
.Y(n_7846)
);

INVx2_ASAP7_75t_L g7847 ( 
.A(n_7080),
.Y(n_7847)
);

INVx2_ASAP7_75t_L g7848 ( 
.A(n_7093),
.Y(n_7848)
);

INVx1_ASAP7_75t_L g7849 ( 
.A(n_6790),
.Y(n_7849)
);

AOI22xp33_ASAP7_75t_L g7850 ( 
.A1(n_6699),
.A2(n_6319),
.B1(n_5720),
.B2(n_5765),
.Y(n_7850)
);

AND2x2_ASAP7_75t_L g7851 ( 
.A(n_6448),
.B(n_6268),
.Y(n_7851)
);

AOI22xp33_ASAP7_75t_L g7852 ( 
.A1(n_6698),
.A2(n_5720),
.B1(n_5765),
.B2(n_5883),
.Y(n_7852)
);

AOI22xp33_ASAP7_75t_L g7853 ( 
.A1(n_6698),
.A2(n_5720),
.B1(n_5765),
.B2(n_5883),
.Y(n_7853)
);

INVx1_ASAP7_75t_L g7854 ( 
.A(n_6804),
.Y(n_7854)
);

NAND2x1p5_ASAP7_75t_L g7855 ( 
.A(n_7008),
.B(n_5882),
.Y(n_7855)
);

INVx2_ASAP7_75t_L g7856 ( 
.A(n_7093),
.Y(n_7856)
);

AOI22xp33_ASAP7_75t_L g7857 ( 
.A1(n_6613),
.A2(n_5720),
.B1(n_5765),
.B2(n_6007),
.Y(n_7857)
);

AOI22xp33_ASAP7_75t_L g7858 ( 
.A1(n_6613),
.A2(n_5720),
.B1(n_5765),
.B2(n_6239),
.Y(n_7858)
);

INVx1_ASAP7_75t_L g7859 ( 
.A(n_6804),
.Y(n_7859)
);

INVx6_ASAP7_75t_L g7860 ( 
.A(n_6774),
.Y(n_7860)
);

AND2x4_ASAP7_75t_L g7861 ( 
.A(n_6951),
.B(n_6297),
.Y(n_7861)
);

INVx1_ASAP7_75t_L g7862 ( 
.A(n_6810),
.Y(n_7862)
);

BUFx12f_ASAP7_75t_L g7863 ( 
.A(n_6539),
.Y(n_7863)
);

NAND2x1p5_ASAP7_75t_L g7864 ( 
.A(n_7008),
.B(n_5882),
.Y(n_7864)
);

AND2x4_ASAP7_75t_L g7865 ( 
.A(n_6951),
.B(n_6297),
.Y(n_7865)
);

AOI21x1_ASAP7_75t_L g7866 ( 
.A1(n_6456),
.A2(n_6218),
.B(n_6194),
.Y(n_7866)
);

INVx2_ASAP7_75t_L g7867 ( 
.A(n_7093),
.Y(n_7867)
);

INVx2_ASAP7_75t_L g7868 ( 
.A(n_7093),
.Y(n_7868)
);

INVx2_ASAP7_75t_L g7869 ( 
.A(n_7114),
.Y(n_7869)
);

OR2x2_ASAP7_75t_L g7870 ( 
.A(n_6649),
.B(n_5987),
.Y(n_7870)
);

AND2x2_ASAP7_75t_L g7871 ( 
.A(n_6448),
.B(n_6487),
.Y(n_7871)
);

HB1xp67_ASAP7_75t_L g7872 ( 
.A(n_6828),
.Y(n_7872)
);

AOI22xp33_ASAP7_75t_L g7873 ( 
.A1(n_7130),
.A2(n_5720),
.B1(n_5765),
.B2(n_6239),
.Y(n_7873)
);

INVx5_ASAP7_75t_L g7874 ( 
.A(n_6539),
.Y(n_7874)
);

INVx1_ASAP7_75t_L g7875 ( 
.A(n_6810),
.Y(n_7875)
);

AOI22xp33_ASAP7_75t_L g7876 ( 
.A1(n_7137),
.A2(n_6301),
.B1(n_6356),
.B2(n_6307),
.Y(n_7876)
);

INVx1_ASAP7_75t_SL g7877 ( 
.A(n_7179),
.Y(n_7877)
);

NOR2xp33_ASAP7_75t_L g7878 ( 
.A(n_7142),
.B(n_5907),
.Y(n_7878)
);

AOI22xp33_ASAP7_75t_L g7879 ( 
.A1(n_7137),
.A2(n_6301),
.B1(n_6356),
.B2(n_6307),
.Y(n_7879)
);

INVx1_ASAP7_75t_L g7880 ( 
.A(n_6832),
.Y(n_7880)
);

INVx1_ASAP7_75t_L g7881 ( 
.A(n_6832),
.Y(n_7881)
);

INVx2_ASAP7_75t_L g7882 ( 
.A(n_7114),
.Y(n_7882)
);

CKINVDCx20_ASAP7_75t_R g7883 ( 
.A(n_7120),
.Y(n_7883)
);

BUFx2_ASAP7_75t_L g7884 ( 
.A(n_6632),
.Y(n_7884)
);

INVx4_ASAP7_75t_L g7885 ( 
.A(n_6824),
.Y(n_7885)
);

OAI22xp5_ASAP7_75t_L g7886 ( 
.A1(n_6514),
.A2(n_5957),
.B1(n_5736),
.B2(n_6059),
.Y(n_7886)
);

OAI21x1_ASAP7_75t_L g7887 ( 
.A1(n_6504),
.A2(n_5994),
.B(n_5989),
.Y(n_7887)
);

INVx1_ASAP7_75t_L g7888 ( 
.A(n_6835),
.Y(n_7888)
);

INVx1_ASAP7_75t_L g7889 ( 
.A(n_6835),
.Y(n_7889)
);

OAI22xp33_ASAP7_75t_L g7890 ( 
.A1(n_6884),
.A2(n_6070),
.B1(n_6049),
.B2(n_5888),
.Y(n_7890)
);

AOI22xp33_ASAP7_75t_L g7891 ( 
.A1(n_6648),
.A2(n_6301),
.B1(n_6356),
.B2(n_6307),
.Y(n_7891)
);

HB1xp67_ASAP7_75t_L g7892 ( 
.A(n_6828),
.Y(n_7892)
);

AOI21xp5_ASAP7_75t_L g7893 ( 
.A1(n_6515),
.A2(n_6158),
.B(n_6386),
.Y(n_7893)
);

BUFx6f_ASAP7_75t_L g7894 ( 
.A(n_6520),
.Y(n_7894)
);

INVx3_ASAP7_75t_L g7895 ( 
.A(n_7102),
.Y(n_7895)
);

AO21x1_ASAP7_75t_L g7896 ( 
.A1(n_6469),
.A2(n_6507),
.B(n_6890),
.Y(n_7896)
);

INVx2_ASAP7_75t_L g7897 ( 
.A(n_7114),
.Y(n_7897)
);

OAI21x1_ASAP7_75t_L g7898 ( 
.A1(n_6504),
.A2(n_6000),
.B(n_5994),
.Y(n_7898)
);

BUFx12f_ASAP7_75t_L g7899 ( 
.A(n_6539),
.Y(n_7899)
);

AOI22xp33_ASAP7_75t_L g7900 ( 
.A1(n_6648),
.A2(n_7348),
.B1(n_7271),
.B2(n_7207),
.Y(n_7900)
);

AOI22xp33_ASAP7_75t_L g7901 ( 
.A1(n_7271),
.A2(n_6307),
.B1(n_6413),
.B2(n_6356),
.Y(n_7901)
);

OA21x2_ASAP7_75t_L g7902 ( 
.A1(n_6450),
.A2(n_6255),
.B(n_6218),
.Y(n_7902)
);

INVx2_ASAP7_75t_SL g7903 ( 
.A(n_6534),
.Y(n_7903)
);

AO21x2_ASAP7_75t_L g7904 ( 
.A1(n_6450),
.A2(n_5722),
.B(n_5702),
.Y(n_7904)
);

AND2x4_ASAP7_75t_L g7905 ( 
.A(n_6951),
.B(n_6413),
.Y(n_7905)
);

OAI21x1_ASAP7_75t_L g7906 ( 
.A1(n_6504),
.A2(n_6000),
.B(n_5994),
.Y(n_7906)
);

HB1xp67_ASAP7_75t_L g7907 ( 
.A(n_6829),
.Y(n_7907)
);

INVx6_ASAP7_75t_L g7908 ( 
.A(n_6774),
.Y(n_7908)
);

INVx1_ASAP7_75t_L g7909 ( 
.A(n_6845),
.Y(n_7909)
);

INVx1_ASAP7_75t_L g7910 ( 
.A(n_6845),
.Y(n_7910)
);

INVx1_ASAP7_75t_L g7911 ( 
.A(n_6848),
.Y(n_7911)
);

INVx2_ASAP7_75t_L g7912 ( 
.A(n_7114),
.Y(n_7912)
);

OAI21x1_ASAP7_75t_L g7913 ( 
.A1(n_6997),
.A2(n_6000),
.B(n_5994),
.Y(n_7913)
);

BUFx3_ASAP7_75t_L g7914 ( 
.A(n_7004),
.Y(n_7914)
);

INVx1_ASAP7_75t_L g7915 ( 
.A(n_6848),
.Y(n_7915)
);

INVx3_ASAP7_75t_L g7916 ( 
.A(n_7102),
.Y(n_7916)
);

AOI22xp33_ASAP7_75t_L g7917 ( 
.A1(n_7207),
.A2(n_6413),
.B1(n_6433),
.B2(n_5927),
.Y(n_7917)
);

AOI22xp5_ASAP7_75t_L g7918 ( 
.A1(n_6731),
.A2(n_5888),
.B1(n_5917),
.B2(n_6059),
.Y(n_7918)
);

INVx1_ASAP7_75t_L g7919 ( 
.A(n_6865),
.Y(n_7919)
);

INVx2_ASAP7_75t_SL g7920 ( 
.A(n_6534),
.Y(n_7920)
);

NAND2xp5_ASAP7_75t_L g7921 ( 
.A(n_6731),
.B(n_6027),
.Y(n_7921)
);

INVx1_ASAP7_75t_L g7922 ( 
.A(n_6865),
.Y(n_7922)
);

INVx1_ASAP7_75t_L g7923 ( 
.A(n_6868),
.Y(n_7923)
);

INVx1_ASAP7_75t_SL g7924 ( 
.A(n_6593),
.Y(n_7924)
);

AOI21x1_ASAP7_75t_L g7925 ( 
.A1(n_6456),
.A2(n_6255),
.B(n_6218),
.Y(n_7925)
);

INVx1_ASAP7_75t_L g7926 ( 
.A(n_6868),
.Y(n_7926)
);

OAI22xp5_ASAP7_75t_L g7927 ( 
.A1(n_6583),
.A2(n_5957),
.B1(n_6381),
.B2(n_6317),
.Y(n_7927)
);

AND2x2_ASAP7_75t_L g7928 ( 
.A(n_6448),
.B(n_6487),
.Y(n_7928)
);

BUFx2_ASAP7_75t_R g7929 ( 
.A(n_6502),
.Y(n_7929)
);

OA21x2_ASAP7_75t_L g7930 ( 
.A1(n_6450),
.A2(n_6260),
.B(n_6255),
.Y(n_7930)
);

INVx6_ASAP7_75t_L g7931 ( 
.A(n_7004),
.Y(n_7931)
);

CKINVDCx11_ASAP7_75t_R g7932 ( 
.A(n_6593),
.Y(n_7932)
);

INVx1_ASAP7_75t_L g7933 ( 
.A(n_6880),
.Y(n_7933)
);

INVx3_ASAP7_75t_L g7934 ( 
.A(n_7115),
.Y(n_7934)
);

INVx1_ASAP7_75t_L g7935 ( 
.A(n_6880),
.Y(n_7935)
);

BUFx2_ASAP7_75t_SL g7936 ( 
.A(n_6632),
.Y(n_7936)
);

AOI22xp33_ASAP7_75t_L g7937 ( 
.A1(n_7207),
.A2(n_6601),
.B1(n_7037),
.B2(n_6805),
.Y(n_7937)
);

CKINVDCx5p33_ASAP7_75t_R g7938 ( 
.A(n_6663),
.Y(n_7938)
);

NAND2xp5_ASAP7_75t_L g7939 ( 
.A(n_6874),
.B(n_6109),
.Y(n_7939)
);

NAND2x1p5_ASAP7_75t_L g7940 ( 
.A(n_7008),
.B(n_5882),
.Y(n_7940)
);

AOI22xp33_ASAP7_75t_L g7941 ( 
.A1(n_7207),
.A2(n_6413),
.B1(n_6433),
.B2(n_5927),
.Y(n_7941)
);

INVx1_ASAP7_75t_L g7942 ( 
.A(n_6886),
.Y(n_7942)
);

INVx2_ASAP7_75t_L g7943 ( 
.A(n_7146),
.Y(n_7943)
);

INVx1_ASAP7_75t_SL g7944 ( 
.A(n_6690),
.Y(n_7944)
);

INVx2_ASAP7_75t_L g7945 ( 
.A(n_7146),
.Y(n_7945)
);

NAND2xp5_ASAP7_75t_L g7946 ( 
.A(n_6874),
.B(n_6109),
.Y(n_7946)
);

OAI22xp5_ASAP7_75t_L g7947 ( 
.A1(n_7207),
.A2(n_6325),
.B1(n_6381),
.B2(n_6317),
.Y(n_7947)
);

AOI22xp33_ASAP7_75t_L g7948 ( 
.A1(n_6601),
.A2(n_7037),
.B1(n_6805),
.B2(n_6673),
.Y(n_7948)
);

INVx2_ASAP7_75t_L g7949 ( 
.A(n_7146),
.Y(n_7949)
);

BUFx6f_ASAP7_75t_L g7950 ( 
.A(n_6534),
.Y(n_7950)
);

INVx1_ASAP7_75t_L g7951 ( 
.A(n_6886),
.Y(n_7951)
);

INVx1_ASAP7_75t_SL g7952 ( 
.A(n_6690),
.Y(n_7952)
);

INVx2_ASAP7_75t_L g7953 ( 
.A(n_7146),
.Y(n_7953)
);

INVx2_ASAP7_75t_L g7954 ( 
.A(n_7146),
.Y(n_7954)
);

AND2x4_ASAP7_75t_L g7955 ( 
.A(n_6951),
.B(n_6433),
.Y(n_7955)
);

OR2x2_ASAP7_75t_L g7956 ( 
.A(n_6453),
.B(n_6030),
.Y(n_7956)
);

INVx2_ASAP7_75t_L g7957 ( 
.A(n_6897),
.Y(n_7957)
);

AOI22xp5_ASAP7_75t_L g7958 ( 
.A1(n_6678),
.A2(n_5917),
.B1(n_6229),
.B2(n_5595),
.Y(n_7958)
);

BUFx2_ASAP7_75t_SL g7959 ( 
.A(n_6632),
.Y(n_7959)
);

BUFx2_ASAP7_75t_SL g7960 ( 
.A(n_6632),
.Y(n_7960)
);

INVx2_ASAP7_75t_L g7961 ( 
.A(n_6897),
.Y(n_7961)
);

NAND2xp5_ASAP7_75t_L g7962 ( 
.A(n_6878),
.B(n_6110),
.Y(n_7962)
);

BUFx6f_ASAP7_75t_L g7963 ( 
.A(n_6544),
.Y(n_7963)
);

AO21x2_ASAP7_75t_L g7964 ( 
.A1(n_6460),
.A2(n_5722),
.B(n_5782),
.Y(n_7964)
);

AOI22xp33_ASAP7_75t_SL g7965 ( 
.A1(n_6881),
.A2(n_6433),
.B1(n_5545),
.B2(n_6264),
.Y(n_7965)
);

INVx1_ASAP7_75t_L g7966 ( 
.A(n_6900),
.Y(n_7966)
);

INVx2_ASAP7_75t_L g7967 ( 
.A(n_6897),
.Y(n_7967)
);

INVx3_ASAP7_75t_L g7968 ( 
.A(n_7115),
.Y(n_7968)
);

BUFx2_ASAP7_75t_R g7969 ( 
.A(n_6704),
.Y(n_7969)
);

INVx1_ASAP7_75t_L g7970 ( 
.A(n_6900),
.Y(n_7970)
);

INVx1_ASAP7_75t_L g7971 ( 
.A(n_6905),
.Y(n_7971)
);

INVx1_ASAP7_75t_L g7972 ( 
.A(n_6905),
.Y(n_7972)
);

INVx2_ASAP7_75t_L g7973 ( 
.A(n_6897),
.Y(n_7973)
);

INVx2_ASAP7_75t_L g7974 ( 
.A(n_7362),
.Y(n_7974)
);

AOI22xp33_ASAP7_75t_L g7975 ( 
.A1(n_7037),
.A2(n_6673),
.B1(n_6570),
.B2(n_6493),
.Y(n_7975)
);

INVx1_ASAP7_75t_SL g7976 ( 
.A(n_6729),
.Y(n_7976)
);

INVx2_ASAP7_75t_L g7977 ( 
.A(n_6895),
.Y(n_7977)
);

INVx3_ASAP7_75t_L g7978 ( 
.A(n_7115),
.Y(n_7978)
);

AOI22xp33_ASAP7_75t_L g7979 ( 
.A1(n_7037),
.A2(n_6570),
.B1(n_6493),
.B2(n_6470),
.Y(n_7979)
);

INVx1_ASAP7_75t_L g7980 ( 
.A(n_6934),
.Y(n_7980)
);

AO21x1_ASAP7_75t_L g7981 ( 
.A1(n_6890),
.A2(n_5808),
.B(n_5807),
.Y(n_7981)
);

INVx1_ASAP7_75t_L g7982 ( 
.A(n_6934),
.Y(n_7982)
);

INVx2_ASAP7_75t_L g7983 ( 
.A(n_6895),
.Y(n_7983)
);

AND2x2_ASAP7_75t_L g7984 ( 
.A(n_6487),
.B(n_5933),
.Y(n_7984)
);

CKINVDCx11_ASAP7_75t_R g7985 ( 
.A(n_6729),
.Y(n_7985)
);

AOI21xp33_ASAP7_75t_L g7986 ( 
.A1(n_6767),
.A2(n_6333),
.B(n_6207),
.Y(n_7986)
);

OAI22xp33_ASAP7_75t_L g7987 ( 
.A1(n_6884),
.A2(n_6236),
.B1(n_6264),
.B2(n_5781),
.Y(n_7987)
);

INVx6_ASAP7_75t_L g7988 ( 
.A(n_7004),
.Y(n_7988)
);

OA21x2_ASAP7_75t_L g7989 ( 
.A1(n_6460),
.A2(n_6289),
.B(n_6260),
.Y(n_7989)
);

HB1xp67_ASAP7_75t_L g7990 ( 
.A(n_6829),
.Y(n_7990)
);

OAI22xp5_ASAP7_75t_L g7991 ( 
.A1(n_6587),
.A2(n_6325),
.B1(n_6381),
.B2(n_6317),
.Y(n_7991)
);

INVx1_ASAP7_75t_L g7992 ( 
.A(n_6958),
.Y(n_7992)
);

INVx2_ASAP7_75t_SL g7993 ( 
.A(n_6544),
.Y(n_7993)
);

INVx2_ASAP7_75t_L g7994 ( 
.A(n_6895),
.Y(n_7994)
);

INVx1_ASAP7_75t_L g7995 ( 
.A(n_6958),
.Y(n_7995)
);

INVx2_ASAP7_75t_L g7996 ( 
.A(n_6895),
.Y(n_7996)
);

HB1xp67_ASAP7_75t_L g7997 ( 
.A(n_6902),
.Y(n_7997)
);

AOI22xp33_ASAP7_75t_L g7998 ( 
.A1(n_7037),
.A2(n_5927),
.B1(n_5781),
.B2(n_4740),
.Y(n_7998)
);

INVx1_ASAP7_75t_L g7999 ( 
.A(n_6970),
.Y(n_7999)
);

OA21x2_ASAP7_75t_L g8000 ( 
.A1(n_6460),
.A2(n_6289),
.B(n_6260),
.Y(n_8000)
);

INVx2_ASAP7_75t_SL g8001 ( 
.A(n_6544),
.Y(n_8001)
);

NAND2xp5_ASAP7_75t_L g8002 ( 
.A(n_6878),
.B(n_6110),
.Y(n_8002)
);

INVx2_ASAP7_75t_L g8003 ( 
.A(n_6895),
.Y(n_8003)
);

HB1xp67_ASAP7_75t_L g8004 ( 
.A(n_6902),
.Y(n_8004)
);

CKINVDCx5p33_ASAP7_75t_R g8005 ( 
.A(n_6836),
.Y(n_8005)
);

NAND2x1p5_ASAP7_75t_L g8006 ( 
.A(n_7008),
.B(n_5882),
.Y(n_8006)
);

INVxp67_ASAP7_75t_L g8007 ( 
.A(n_7013),
.Y(n_8007)
);

INVx1_ASAP7_75t_L g8008 ( 
.A(n_6970),
.Y(n_8008)
);

INVx2_ASAP7_75t_L g8009 ( 
.A(n_7362),
.Y(n_8009)
);

HB1xp67_ASAP7_75t_L g8010 ( 
.A(n_7085),
.Y(n_8010)
);

INVx1_ASAP7_75t_L g8011 ( 
.A(n_6973),
.Y(n_8011)
);

BUFx6f_ASAP7_75t_L g8012 ( 
.A(n_6641),
.Y(n_8012)
);

INVx4_ASAP7_75t_L g8013 ( 
.A(n_6824),
.Y(n_8013)
);

BUFx2_ASAP7_75t_R g8014 ( 
.A(n_6883),
.Y(n_8014)
);

OAI22xp5_ASAP7_75t_L g8015 ( 
.A1(n_7308),
.A2(n_6325),
.B1(n_6317),
.B2(n_6381),
.Y(n_8015)
);

NAND2x1p5_ASAP7_75t_L g8016 ( 
.A(n_7061),
.B(n_5882),
.Y(n_8016)
);

OAI21x1_ASAP7_75t_L g8017 ( 
.A1(n_6997),
.A2(n_6016),
.B(n_6000),
.Y(n_8017)
);

INVx1_ASAP7_75t_L g8018 ( 
.A(n_6973),
.Y(n_8018)
);

INVx2_ASAP7_75t_L g8019 ( 
.A(n_7362),
.Y(n_8019)
);

AOI22xp33_ASAP7_75t_L g8020 ( 
.A1(n_6470),
.A2(n_5927),
.B1(n_5781),
.B2(n_4740),
.Y(n_8020)
);

AOI22xp33_ASAP7_75t_L g8021 ( 
.A1(n_6470),
.A2(n_5927),
.B1(n_5781),
.B2(n_4740),
.Y(n_8021)
);

BUFx12f_ASAP7_75t_L g8022 ( 
.A(n_6539),
.Y(n_8022)
);

INVx1_ASAP7_75t_L g8023 ( 
.A(n_6985),
.Y(n_8023)
);

AND2x2_ASAP7_75t_L g8024 ( 
.A(n_6509),
.B(n_5933),
.Y(n_8024)
);

CKINVDCx11_ASAP7_75t_R g8025 ( 
.A(n_6962),
.Y(n_8025)
);

AOI21x1_ASAP7_75t_L g8026 ( 
.A1(n_6457),
.A2(n_6332),
.B(n_6289),
.Y(n_8026)
);

INVx1_ASAP7_75t_L g8027 ( 
.A(n_6985),
.Y(n_8027)
);

AO21x1_ASAP7_75t_SL g8028 ( 
.A1(n_6857),
.A2(n_6115),
.B(n_6135),
.Y(n_8028)
);

INVx2_ASAP7_75t_L g8029 ( 
.A(n_7362),
.Y(n_8029)
);

HB1xp67_ASAP7_75t_L g8030 ( 
.A(n_7085),
.Y(n_8030)
);

INVx6_ASAP7_75t_L g8031 ( 
.A(n_7004),
.Y(n_8031)
);

OAI22xp5_ASAP7_75t_L g8032 ( 
.A1(n_7308),
.A2(n_6325),
.B1(n_6237),
.B2(n_6229),
.Y(n_8032)
);

INVx1_ASAP7_75t_L g8033 ( 
.A(n_6987),
.Y(n_8033)
);

AOI22xp33_ASAP7_75t_SL g8034 ( 
.A1(n_6881),
.A2(n_5545),
.B1(n_6264),
.B2(n_6236),
.Y(n_8034)
);

INVx1_ASAP7_75t_L g8035 ( 
.A(n_6987),
.Y(n_8035)
);

INVx1_ASAP7_75t_L g8036 ( 
.A(n_6989),
.Y(n_8036)
);

CKINVDCx20_ASAP7_75t_R g8037 ( 
.A(n_6921),
.Y(n_8037)
);

NAND2xp5_ASAP7_75t_L g8038 ( 
.A(n_6918),
.B(n_6114),
.Y(n_8038)
);

INVx2_ASAP7_75t_L g8039 ( 
.A(n_7260),
.Y(n_8039)
);

INVx2_ASAP7_75t_L g8040 ( 
.A(n_7260),
.Y(n_8040)
);

NOR2xp33_ASAP7_75t_L g8041 ( 
.A(n_6962),
.B(n_5907),
.Y(n_8041)
);

INVx2_ASAP7_75t_L g8042 ( 
.A(n_7260),
.Y(n_8042)
);

INVx2_ASAP7_75t_L g8043 ( 
.A(n_7260),
.Y(n_8043)
);

AOI22xp33_ASAP7_75t_L g8044 ( 
.A1(n_6470),
.A2(n_5781),
.B1(n_4740),
.B2(n_5694),
.Y(n_8044)
);

CKINVDCx20_ASAP7_75t_R g8045 ( 
.A(n_6962),
.Y(n_8045)
);

OAI22xp5_ASAP7_75t_L g8046 ( 
.A1(n_6619),
.A2(n_6237),
.B1(n_6122),
.B2(n_6156),
.Y(n_8046)
);

INVx1_ASAP7_75t_L g8047 ( 
.A(n_6989),
.Y(n_8047)
);

INVx1_ASAP7_75t_L g8048 ( 
.A(n_6998),
.Y(n_8048)
);

AND2x2_ASAP7_75t_L g8049 ( 
.A(n_6509),
.B(n_6545),
.Y(n_8049)
);

INVx2_ASAP7_75t_L g8050 ( 
.A(n_7274),
.Y(n_8050)
);

AND2x2_ASAP7_75t_SL g8051 ( 
.A(n_7390),
.B(n_6332),
.Y(n_8051)
);

OAI21x1_ASAP7_75t_L g8052 ( 
.A1(n_6997),
.A2(n_6016),
.B(n_6000),
.Y(n_8052)
);

INVx1_ASAP7_75t_L g8053 ( 
.A(n_6998),
.Y(n_8053)
);

BUFx8_ASAP7_75t_L g8054 ( 
.A(n_6641),
.Y(n_8054)
);

INVx1_ASAP7_75t_L g8055 ( 
.A(n_6999),
.Y(n_8055)
);

INVx1_ASAP7_75t_L g8056 ( 
.A(n_6999),
.Y(n_8056)
);

NOR2xp33_ASAP7_75t_L g8057 ( 
.A(n_7211),
.B(n_5907),
.Y(n_8057)
);

OAI22xp5_ASAP7_75t_L g8058 ( 
.A1(n_6619),
.A2(n_6140),
.B1(n_6191),
.B2(n_6156),
.Y(n_8058)
);

AND2x2_ASAP7_75t_L g8059 ( 
.A(n_6509),
.B(n_5933),
.Y(n_8059)
);

INVx1_ASAP7_75t_L g8060 ( 
.A(n_7009),
.Y(n_8060)
);

INVx2_ASAP7_75t_L g8061 ( 
.A(n_6944),
.Y(n_8061)
);

INVx2_ASAP7_75t_L g8062 ( 
.A(n_6944),
.Y(n_8062)
);

INVx4_ASAP7_75t_SL g8063 ( 
.A(n_6660),
.Y(n_8063)
);

NAND2xp5_ASAP7_75t_L g8064 ( 
.A(n_6918),
.B(n_6974),
.Y(n_8064)
);

INVx2_ASAP7_75t_L g8065 ( 
.A(n_6944),
.Y(n_8065)
);

INVx2_ASAP7_75t_L g8066 ( 
.A(n_6944),
.Y(n_8066)
);

INVx1_ASAP7_75t_L g8067 ( 
.A(n_7009),
.Y(n_8067)
);

INVx6_ASAP7_75t_L g8068 ( 
.A(n_7004),
.Y(n_8068)
);

INVx2_ASAP7_75t_L g8069 ( 
.A(n_6944),
.Y(n_8069)
);

CKINVDCx5p33_ASAP7_75t_R g8070 ( 
.A(n_6971),
.Y(n_8070)
);

CKINVDCx6p67_ASAP7_75t_R g8071 ( 
.A(n_6824),
.Y(n_8071)
);

CKINVDCx5p33_ASAP7_75t_R g8072 ( 
.A(n_6971),
.Y(n_8072)
);

BUFx2_ASAP7_75t_SL g8073 ( 
.A(n_6640),
.Y(n_8073)
);

AOI22xp33_ASAP7_75t_L g8074 ( 
.A1(n_6493),
.A2(n_5781),
.B1(n_5582),
.B2(n_5729),
.Y(n_8074)
);

INVx1_ASAP7_75t_SL g8075 ( 
.A(n_7211),
.Y(n_8075)
);

HB1xp67_ASAP7_75t_L g8076 ( 
.A(n_7182),
.Y(n_8076)
);

INVx3_ASAP7_75t_L g8077 ( 
.A(n_7115),
.Y(n_8077)
);

NAND3xp33_ASAP7_75t_SL g8078 ( 
.A(n_6837),
.B(n_6133),
.C(n_6114),
.Y(n_8078)
);

AOI22xp5_ASAP7_75t_L g8079 ( 
.A1(n_6678),
.A2(n_5595),
.B1(n_6333),
.B2(n_6293),
.Y(n_8079)
);

INVx1_ASAP7_75t_SL g8080 ( 
.A(n_7176),
.Y(n_8080)
);

NAND2xp5_ASAP7_75t_L g8081 ( 
.A(n_6974),
.B(n_6133),
.Y(n_8081)
);

INVx1_ASAP7_75t_L g8082 ( 
.A(n_7011),
.Y(n_8082)
);

OAI21x1_ASAP7_75t_L g8083 ( 
.A1(n_6572),
.A2(n_6019),
.B(n_6016),
.Y(n_8083)
);

INVx1_ASAP7_75t_L g8084 ( 
.A(n_7011),
.Y(n_8084)
);

INVx3_ASAP7_75t_L g8085 ( 
.A(n_7115),
.Y(n_8085)
);

AND2x2_ASAP7_75t_L g8086 ( 
.A(n_6545),
.B(n_5933),
.Y(n_8086)
);

INVx2_ASAP7_75t_L g8087 ( 
.A(n_6944),
.Y(n_8087)
);

INVx1_ASAP7_75t_L g8088 ( 
.A(n_7027),
.Y(n_8088)
);

BUFx6f_ASAP7_75t_L g8089 ( 
.A(n_6641),
.Y(n_8089)
);

INVx1_ASAP7_75t_L g8090 ( 
.A(n_7027),
.Y(n_8090)
);

INVx2_ASAP7_75t_L g8091 ( 
.A(n_6944),
.Y(n_8091)
);

INVx2_ASAP7_75t_L g8092 ( 
.A(n_6992),
.Y(n_8092)
);

INVx1_ASAP7_75t_L g8093 ( 
.A(n_7035),
.Y(n_8093)
);

BUFx2_ASAP7_75t_L g8094 ( 
.A(n_6640),
.Y(n_8094)
);

OAI22xp5_ASAP7_75t_L g8095 ( 
.A1(n_7317),
.A2(n_6140),
.B1(n_6199),
.B2(n_6191),
.Y(n_8095)
);

INVx6_ASAP7_75t_L g8096 ( 
.A(n_6539),
.Y(n_8096)
);

BUFx8_ASAP7_75t_L g8097 ( 
.A(n_6661),
.Y(n_8097)
);

AOI22xp5_ASAP7_75t_L g8098 ( 
.A1(n_7317),
.A2(n_6397),
.B1(n_6293),
.B2(n_6418),
.Y(n_8098)
);

OR2x2_ASAP7_75t_L g8099 ( 
.A(n_6453),
.B(n_6475),
.Y(n_8099)
);

AOI22xp33_ASAP7_75t_SL g8100 ( 
.A1(n_6881),
.A2(n_5545),
.B1(n_6264),
.B2(n_6236),
.Y(n_8100)
);

CKINVDCx11_ASAP7_75t_R g8101 ( 
.A(n_6640),
.Y(n_8101)
);

OAI21xp5_ASAP7_75t_L g8102 ( 
.A1(n_6837),
.A2(n_6162),
.B(n_6148),
.Y(n_8102)
);

INVx1_ASAP7_75t_L g8103 ( 
.A(n_7035),
.Y(n_8103)
);

OAI22xp5_ASAP7_75t_L g8104 ( 
.A1(n_6769),
.A2(n_6140),
.B1(n_6199),
.B2(n_6191),
.Y(n_8104)
);

BUFx6f_ASAP7_75t_L g8105 ( 
.A(n_6661),
.Y(n_8105)
);

INVx2_ASAP7_75t_L g8106 ( 
.A(n_7274),
.Y(n_8106)
);

HB1xp67_ASAP7_75t_L g8107 ( 
.A(n_7182),
.Y(n_8107)
);

INVx2_ASAP7_75t_L g8108 ( 
.A(n_7274),
.Y(n_8108)
);

AOI22xp33_ASAP7_75t_L g8109 ( 
.A1(n_6493),
.A2(n_5781),
.B1(n_5582),
.B2(n_5729),
.Y(n_8109)
);

OAI21xp5_ASAP7_75t_L g8110 ( 
.A1(n_7001),
.A2(n_6162),
.B(n_6332),
.Y(n_8110)
);

BUFx12f_ASAP7_75t_L g8111 ( 
.A(n_6640),
.Y(n_8111)
);

OA21x2_ASAP7_75t_L g8112 ( 
.A1(n_6532),
.A2(n_6342),
.B(n_6339),
.Y(n_8112)
);

BUFx6f_ASAP7_75t_L g8113 ( 
.A(n_6661),
.Y(n_8113)
);

INVxp67_ASAP7_75t_SL g8114 ( 
.A(n_6911),
.Y(n_8114)
);

OR2x2_ASAP7_75t_L g8115 ( 
.A(n_6475),
.B(n_6030),
.Y(n_8115)
);

INVx3_ASAP7_75t_L g8116 ( 
.A(n_7152),
.Y(n_8116)
);

HB1xp67_ASAP7_75t_L g8117 ( 
.A(n_7236),
.Y(n_8117)
);

INVx1_ASAP7_75t_L g8118 ( 
.A(n_7043),
.Y(n_8118)
);

OAI22xp33_ASAP7_75t_L g8119 ( 
.A1(n_6744),
.A2(n_6236),
.B1(n_5550),
.B2(n_5694),
.Y(n_8119)
);

INVxp67_ASAP7_75t_SL g8120 ( 
.A(n_6911),
.Y(n_8120)
);

AOI22xp33_ASAP7_75t_SL g8121 ( 
.A1(n_6881),
.A2(n_5545),
.B1(n_5699),
.B2(n_5666),
.Y(n_8121)
);

INVx2_ASAP7_75t_L g8122 ( 
.A(n_7274),
.Y(n_8122)
);

INVx6_ASAP7_75t_L g8123 ( 
.A(n_6640),
.Y(n_8123)
);

INVxp67_ASAP7_75t_SL g8124 ( 
.A(n_6912),
.Y(n_8124)
);

AOI22xp33_ASAP7_75t_L g8125 ( 
.A1(n_7044),
.A2(n_5582),
.B1(n_5729),
.B2(n_5694),
.Y(n_8125)
);

AND2x2_ASAP7_75t_L g8126 ( 
.A(n_6545),
.B(n_5933),
.Y(n_8126)
);

INVx2_ASAP7_75t_L g8127 ( 
.A(n_7280),
.Y(n_8127)
);

HB1xp67_ASAP7_75t_L g8128 ( 
.A(n_7236),
.Y(n_8128)
);

AOI21x1_ASAP7_75t_L g8129 ( 
.A1(n_6457),
.A2(n_6342),
.B(n_6339),
.Y(n_8129)
);

NOR2xp33_ASAP7_75t_L g8130 ( 
.A(n_6931),
.B(n_6077),
.Y(n_8130)
);

INVx2_ASAP7_75t_L g8131 ( 
.A(n_7280),
.Y(n_8131)
);

INVx2_ASAP7_75t_L g8132 ( 
.A(n_7280),
.Y(n_8132)
);

AND2x4_ASAP7_75t_L g8133 ( 
.A(n_6951),
.B(n_5858),
.Y(n_8133)
);

OR2x2_ASAP7_75t_L g8134 ( 
.A(n_6475),
.B(n_6030),
.Y(n_8134)
);

AOI22xp33_ASAP7_75t_L g8135 ( 
.A1(n_7044),
.A2(n_5582),
.B1(n_5729),
.B2(n_5694),
.Y(n_8135)
);

OA21x2_ASAP7_75t_L g8136 ( 
.A1(n_6532),
.A2(n_6342),
.B(n_6339),
.Y(n_8136)
);

INVx2_ASAP7_75t_L g8137 ( 
.A(n_7280),
.Y(n_8137)
);

NAND2x1p5_ASAP7_75t_L g8138 ( 
.A(n_7061),
.B(n_5882),
.Y(n_8138)
);

INVx2_ASAP7_75t_L g8139 ( 
.A(n_6992),
.Y(n_8139)
);

BUFx2_ASAP7_75t_L g8140 ( 
.A(n_6931),
.Y(n_8140)
);

INVx1_ASAP7_75t_L g8141 ( 
.A(n_7043),
.Y(n_8141)
);

AOI21x1_ASAP7_75t_L g8142 ( 
.A1(n_6457),
.A2(n_6382),
.B(n_6346),
.Y(n_8142)
);

INVx6_ASAP7_75t_L g8143 ( 
.A(n_6931),
.Y(n_8143)
);

AOI22xp33_ASAP7_75t_SL g8144 ( 
.A1(n_6881),
.A2(n_5545),
.B1(n_5699),
.B2(n_5666),
.Y(n_8144)
);

BUFx3_ASAP7_75t_L g8145 ( 
.A(n_7169),
.Y(n_8145)
);

INVx2_ASAP7_75t_L g8146 ( 
.A(n_7287),
.Y(n_8146)
);

OAI22xp5_ASAP7_75t_SL g8147 ( 
.A1(n_6660),
.A2(n_6397),
.B1(n_6198),
.B2(n_6274),
.Y(n_8147)
);

OAI21x1_ASAP7_75t_L g8148 ( 
.A1(n_6572),
.A2(n_6019),
.B(n_6016),
.Y(n_8148)
);

INVx2_ASAP7_75t_SL g8149 ( 
.A(n_7169),
.Y(n_8149)
);

INVx2_ASAP7_75t_L g8150 ( 
.A(n_6992),
.Y(n_8150)
);

BUFx6f_ASAP7_75t_L g8151 ( 
.A(n_6683),
.Y(n_8151)
);

INVx2_ASAP7_75t_L g8152 ( 
.A(n_6992),
.Y(n_8152)
);

HB1xp67_ASAP7_75t_L g8153 ( 
.A(n_7242),
.Y(n_8153)
);

INVx1_ASAP7_75t_L g8154 ( 
.A(n_7058),
.Y(n_8154)
);

NAND2xp5_ASAP7_75t_L g8155 ( 
.A(n_6963),
.B(n_6541),
.Y(n_8155)
);

AOI21x1_ASAP7_75t_L g8156 ( 
.A1(n_6481),
.A2(n_6382),
.B(n_6346),
.Y(n_8156)
);

INVx1_ASAP7_75t_L g8157 ( 
.A(n_7058),
.Y(n_8157)
);

INVx1_ASAP7_75t_L g8158 ( 
.A(n_7070),
.Y(n_8158)
);

INVx1_ASAP7_75t_L g8159 ( 
.A(n_7070),
.Y(n_8159)
);

INVx2_ASAP7_75t_L g8160 ( 
.A(n_7287),
.Y(n_8160)
);

INVx1_ASAP7_75t_L g8161 ( 
.A(n_7071),
.Y(n_8161)
);

NAND2xp5_ASAP7_75t_L g8162 ( 
.A(n_6963),
.B(n_6160),
.Y(n_8162)
);

INVx2_ASAP7_75t_L g8163 ( 
.A(n_6992),
.Y(n_8163)
);

NAND2x1p5_ASAP7_75t_L g8164 ( 
.A(n_7061),
.B(n_7237),
.Y(n_8164)
);

INVx6_ASAP7_75t_L g8165 ( 
.A(n_6931),
.Y(n_8165)
);

INVx1_ASAP7_75t_L g8166 ( 
.A(n_7071),
.Y(n_8166)
);

NAND2x1p5_ASAP7_75t_L g8167 ( 
.A(n_7061),
.B(n_5884),
.Y(n_8167)
);

OAI22xp5_ASAP7_75t_L g8168 ( 
.A1(n_6769),
.A2(n_6199),
.B1(n_6282),
.B2(n_6256),
.Y(n_8168)
);

INVx1_ASAP7_75t_L g8169 ( 
.A(n_7078),
.Y(n_8169)
);

INVx1_ASAP7_75t_L g8170 ( 
.A(n_7078),
.Y(n_8170)
);

AOI21x1_ASAP7_75t_L g8171 ( 
.A1(n_6481),
.A2(n_6382),
.B(n_6346),
.Y(n_8171)
);

NAND2x1_ASAP7_75t_L g8172 ( 
.A(n_7106),
.B(n_7126),
.Y(n_8172)
);

INVx1_ASAP7_75t_L g8173 ( 
.A(n_7083),
.Y(n_8173)
);

AO21x2_ASAP7_75t_L g8174 ( 
.A1(n_7157),
.A2(n_5796),
.B(n_5782),
.Y(n_8174)
);

AND2x2_ASAP7_75t_L g8175 ( 
.A(n_6591),
.B(n_6004),
.Y(n_8175)
);

AOI21x1_ASAP7_75t_L g8176 ( 
.A1(n_6481),
.A2(n_6400),
.B(n_6392),
.Y(n_8176)
);

INVx1_ASAP7_75t_L g8177 ( 
.A(n_7083),
.Y(n_8177)
);

BUFx4f_ASAP7_75t_L g8178 ( 
.A(n_7169),
.Y(n_8178)
);

INVx1_ASAP7_75t_L g8179 ( 
.A(n_7087),
.Y(n_8179)
);

INVx1_ASAP7_75t_L g8180 ( 
.A(n_7087),
.Y(n_8180)
);

BUFx2_ASAP7_75t_L g8181 ( 
.A(n_6931),
.Y(n_8181)
);

INVx2_ASAP7_75t_SL g8182 ( 
.A(n_7169),
.Y(n_8182)
);

INVx1_ASAP7_75t_L g8183 ( 
.A(n_7089),
.Y(n_8183)
);

BUFx2_ASAP7_75t_L g8184 ( 
.A(n_7350),
.Y(n_8184)
);

INVx2_ASAP7_75t_SL g8185 ( 
.A(n_7169),
.Y(n_8185)
);

AOI22xp33_ASAP7_75t_L g8186 ( 
.A1(n_6465),
.A2(n_5582),
.B1(n_5729),
.B2(n_5694),
.Y(n_8186)
);

INVx1_ASAP7_75t_L g8187 ( 
.A(n_7089),
.Y(n_8187)
);

INVx3_ASAP7_75t_L g8188 ( 
.A(n_7152),
.Y(n_8188)
);

BUFx2_ASAP7_75t_L g8189 ( 
.A(n_7350),
.Y(n_8189)
);

OAI21x1_ASAP7_75t_SL g8190 ( 
.A1(n_6803),
.A2(n_6282),
.B(n_6256),
.Y(n_8190)
);

AOI22xp33_ASAP7_75t_L g8191 ( 
.A1(n_6465),
.A2(n_5792),
.B1(n_5928),
.B2(n_5875),
.Y(n_8191)
);

INVx1_ASAP7_75t_L g8192 ( 
.A(n_7092),
.Y(n_8192)
);

HB1xp67_ASAP7_75t_L g8193 ( 
.A(n_7242),
.Y(n_8193)
);

INVx1_ASAP7_75t_L g8194 ( 
.A(n_7092),
.Y(n_8194)
);

AOI22xp33_ASAP7_75t_L g8195 ( 
.A1(n_6465),
.A2(n_5792),
.B1(n_5928),
.B2(n_5875),
.Y(n_8195)
);

AOI22xp33_ASAP7_75t_L g8196 ( 
.A1(n_6465),
.A2(n_5792),
.B1(n_5928),
.B2(n_5875),
.Y(n_8196)
);

INVx2_ASAP7_75t_L g8197 ( 
.A(n_7287),
.Y(n_8197)
);

NAND2xp5_ASAP7_75t_L g8198 ( 
.A(n_6541),
.B(n_6160),
.Y(n_8198)
);

BUFx4f_ASAP7_75t_SL g8199 ( 
.A(n_6683),
.Y(n_8199)
);

HB1xp67_ASAP7_75t_L g8200 ( 
.A(n_7318),
.Y(n_8200)
);

INVx4_ASAP7_75t_L g8201 ( 
.A(n_7169),
.Y(n_8201)
);

INVx1_ASAP7_75t_L g8202 ( 
.A(n_7100),
.Y(n_8202)
);

INVx2_ASAP7_75t_L g8203 ( 
.A(n_7287),
.Y(n_8203)
);

INVx1_ASAP7_75t_L g8204 ( 
.A(n_7100),
.Y(n_8204)
);

HB1xp67_ASAP7_75t_L g8205 ( 
.A(n_7318),
.Y(n_8205)
);

BUFx6f_ASAP7_75t_L g8206 ( 
.A(n_6683),
.Y(n_8206)
);

INVx2_ASAP7_75t_L g8207 ( 
.A(n_7305),
.Y(n_8207)
);

INVx2_ASAP7_75t_L g8208 ( 
.A(n_7305),
.Y(n_8208)
);

OA21x2_ASAP7_75t_L g8209 ( 
.A1(n_6532),
.A2(n_6400),
.B(n_6392),
.Y(n_8209)
);

BUFx6f_ASAP7_75t_L g8210 ( 
.A(n_6854),
.Y(n_8210)
);

OAI22xp33_ASAP7_75t_L g8211 ( 
.A1(n_6744),
.A2(n_5550),
.B1(n_5998),
.B2(n_5950),
.Y(n_8211)
);

OAI21x1_ASAP7_75t_L g8212 ( 
.A1(n_6572),
.A2(n_6019),
.B(n_6016),
.Y(n_8212)
);

INVx1_ASAP7_75t_L g8213 ( 
.A(n_7116),
.Y(n_8213)
);

BUFx2_ASAP7_75t_SL g8214 ( 
.A(n_7110),
.Y(n_8214)
);

BUFx6f_ASAP7_75t_L g8215 ( 
.A(n_6854),
.Y(n_8215)
);

INVx1_ASAP7_75t_L g8216 ( 
.A(n_7116),
.Y(n_8216)
);

AOI22xp33_ASAP7_75t_SL g8217 ( 
.A1(n_6500),
.A2(n_5666),
.B1(n_5699),
.B2(n_5706),
.Y(n_8217)
);

BUFx12f_ASAP7_75t_L g8218 ( 
.A(n_7057),
.Y(n_8218)
);

AND2x2_ASAP7_75t_L g8219 ( 
.A(n_6591),
.B(n_6004),
.Y(n_8219)
);

INVxp67_ASAP7_75t_L g8220 ( 
.A(n_7013),
.Y(n_8220)
);

CKINVDCx8_ASAP7_75t_R g8221 ( 
.A(n_7313),
.Y(n_8221)
);

INVx2_ASAP7_75t_L g8222 ( 
.A(n_6992),
.Y(n_8222)
);

INVx2_ASAP7_75t_L g8223 ( 
.A(n_6992),
.Y(n_8223)
);

BUFx6f_ASAP7_75t_L g8224 ( 
.A(n_6854),
.Y(n_8224)
);

OAI22xp5_ASAP7_75t_L g8225 ( 
.A1(n_6789),
.A2(n_6256),
.B1(n_6303),
.B2(n_6282),
.Y(n_8225)
);

OAI21x1_ASAP7_75t_L g8226 ( 
.A1(n_6579),
.A2(n_6021),
.B(n_6019),
.Y(n_8226)
);

INVx2_ASAP7_75t_L g8227 ( 
.A(n_7131),
.Y(n_8227)
);

BUFx2_ASAP7_75t_R g8228 ( 
.A(n_7196),
.Y(n_8228)
);

HB1xp67_ASAP7_75t_L g8229 ( 
.A(n_7360),
.Y(n_8229)
);

INVx1_ASAP7_75t_L g8230 ( 
.A(n_7133),
.Y(n_8230)
);

AND2x2_ASAP7_75t_L g8231 ( 
.A(n_6591),
.B(n_6004),
.Y(n_8231)
);

BUFx3_ASAP7_75t_L g8232 ( 
.A(n_7313),
.Y(n_8232)
);

AOI22xp33_ASAP7_75t_L g8233 ( 
.A1(n_6465),
.A2(n_5792),
.B1(n_5928),
.B2(n_5875),
.Y(n_8233)
);

BUFx2_ASAP7_75t_L g8234 ( 
.A(n_7270),
.Y(n_8234)
);

AOI22xp33_ASAP7_75t_L g8235 ( 
.A1(n_7157),
.A2(n_5792),
.B1(n_5928),
.B2(n_5875),
.Y(n_8235)
);

INVx2_ASAP7_75t_L g8236 ( 
.A(n_7131),
.Y(n_8236)
);

INVx3_ASAP7_75t_L g8237 ( 
.A(n_7152),
.Y(n_8237)
);

AOI22xp33_ASAP7_75t_L g8238 ( 
.A1(n_7157),
.A2(n_5792),
.B1(n_5928),
.B2(n_5875),
.Y(n_8238)
);

OAI22xp5_ASAP7_75t_L g8239 ( 
.A1(n_6789),
.A2(n_6802),
.B1(n_6599),
.B2(n_6830),
.Y(n_8239)
);

OAI22xp5_ASAP7_75t_L g8240 ( 
.A1(n_6802),
.A2(n_6303),
.B1(n_6373),
.B2(n_6313),
.Y(n_8240)
);

INVx1_ASAP7_75t_L g8241 ( 
.A(n_7133),
.Y(n_8241)
);

INVx1_ASAP7_75t_L g8242 ( 
.A(n_7134),
.Y(n_8242)
);

NOR2xp33_ASAP7_75t_L g8243 ( 
.A(n_7019),
.B(n_6077),
.Y(n_8243)
);

INVx2_ASAP7_75t_L g8244 ( 
.A(n_7131),
.Y(n_8244)
);

BUFx2_ASAP7_75t_L g8245 ( 
.A(n_7270),
.Y(n_8245)
);

OA21x2_ASAP7_75t_L g8246 ( 
.A1(n_6474),
.A2(n_6400),
.B(n_6392),
.Y(n_8246)
);

INVx6_ASAP7_75t_L g8247 ( 
.A(n_6665),
.Y(n_8247)
);

INVx4_ASAP7_75t_L g8248 ( 
.A(n_7313),
.Y(n_8248)
);

AND2x2_ASAP7_75t_L g8249 ( 
.A(n_6620),
.B(n_6004),
.Y(n_8249)
);

INVx3_ASAP7_75t_L g8250 ( 
.A(n_7152),
.Y(n_8250)
);

INVx2_ASAP7_75t_L g8251 ( 
.A(n_7305),
.Y(n_8251)
);

INVx1_ASAP7_75t_L g8252 ( 
.A(n_7134),
.Y(n_8252)
);

BUFx10_ASAP7_75t_L g8253 ( 
.A(n_6513),
.Y(n_8253)
);

INVx5_ASAP7_75t_L g8254 ( 
.A(n_6513),
.Y(n_8254)
);

INVx4_ASAP7_75t_L g8255 ( 
.A(n_7313),
.Y(n_8255)
);

BUFx3_ASAP7_75t_L g8256 ( 
.A(n_7313),
.Y(n_8256)
);

INVx1_ASAP7_75t_L g8257 ( 
.A(n_7141),
.Y(n_8257)
);

INVx1_ASAP7_75t_L g8258 ( 
.A(n_7141),
.Y(n_8258)
);

INVx11_ASAP7_75t_L g8259 ( 
.A(n_7313),
.Y(n_8259)
);

HB1xp67_ASAP7_75t_L g8260 ( 
.A(n_7360),
.Y(n_8260)
);

BUFx2_ASAP7_75t_SL g8261 ( 
.A(n_7110),
.Y(n_8261)
);

OR2x2_ASAP7_75t_L g8262 ( 
.A(n_7054),
.B(n_6034),
.Y(n_8262)
);

AOI22xp33_ASAP7_75t_L g8263 ( 
.A1(n_7157),
.A2(n_5792),
.B1(n_5928),
.B2(n_5875),
.Y(n_8263)
);

INVx2_ASAP7_75t_L g8264 ( 
.A(n_7131),
.Y(n_8264)
);

NAND2x1p5_ASAP7_75t_L g8265 ( 
.A(n_7061),
.B(n_5884),
.Y(n_8265)
);

BUFx3_ASAP7_75t_L g8266 ( 
.A(n_7000),
.Y(n_8266)
);

INVx1_ASAP7_75t_L g8267 ( 
.A(n_7147),
.Y(n_8267)
);

OA21x2_ASAP7_75t_L g8268 ( 
.A1(n_6474),
.A2(n_6411),
.B(n_6409),
.Y(n_8268)
);

INVx2_ASAP7_75t_L g8269 ( 
.A(n_7305),
.Y(n_8269)
);

INVx1_ASAP7_75t_L g8270 ( 
.A(n_7147),
.Y(n_8270)
);

INVx1_ASAP7_75t_L g8271 ( 
.A(n_7153),
.Y(n_8271)
);

INVx1_ASAP7_75t_L g8272 ( 
.A(n_7153),
.Y(n_8272)
);

INVx1_ASAP7_75t_L g8273 ( 
.A(n_7155),
.Y(n_8273)
);

INVx1_ASAP7_75t_L g8274 ( 
.A(n_7155),
.Y(n_8274)
);

INVx1_ASAP7_75t_L g8275 ( 
.A(n_7335),
.Y(n_8275)
);

INVx1_ASAP7_75t_L g8276 ( 
.A(n_7335),
.Y(n_8276)
);

NAND2xp5_ASAP7_75t_L g8277 ( 
.A(n_6767),
.B(n_6945),
.Y(n_8277)
);

INVx1_ASAP7_75t_L g8278 ( 
.A(n_7339),
.Y(n_8278)
);

OAI21x1_ASAP7_75t_L g8279 ( 
.A1(n_6579),
.A2(n_6021),
.B(n_6019),
.Y(n_8279)
);

HB1xp67_ASAP7_75t_L g8280 ( 
.A(n_7388),
.Y(n_8280)
);

INVx1_ASAP7_75t_SL g8281 ( 
.A(n_7176),
.Y(n_8281)
);

BUFx2_ASAP7_75t_L g8282 ( 
.A(n_7278),
.Y(n_8282)
);

NAND2xp5_ASAP7_75t_L g8283 ( 
.A(n_6945),
.B(n_6245),
.Y(n_8283)
);

INVx1_ASAP7_75t_L g8284 ( 
.A(n_7339),
.Y(n_8284)
);

INVx2_ASAP7_75t_L g8285 ( 
.A(n_7349),
.Y(n_8285)
);

OAI21x1_ASAP7_75t_L g8286 ( 
.A1(n_6579),
.A2(n_6983),
.B(n_7154),
.Y(n_8286)
);

BUFx6f_ASAP7_75t_L g8287 ( 
.A(n_7000),
.Y(n_8287)
);

INVx1_ASAP7_75t_L g8288 ( 
.A(n_7340),
.Y(n_8288)
);

AOI22xp33_ASAP7_75t_SL g8289 ( 
.A1(n_6500),
.A2(n_5699),
.B1(n_5747),
.B2(n_5706),
.Y(n_8289)
);

AOI22xp33_ASAP7_75t_L g8290 ( 
.A1(n_6686),
.A2(n_5995),
.B1(n_6087),
.B2(n_4865),
.Y(n_8290)
);

BUFx3_ASAP7_75t_L g8291 ( 
.A(n_7000),
.Y(n_8291)
);

AOI22xp33_ASAP7_75t_L g8292 ( 
.A1(n_6686),
.A2(n_5995),
.B1(n_6087),
.B2(n_4865),
.Y(n_8292)
);

OAI21x1_ASAP7_75t_L g8293 ( 
.A1(n_6983),
.A2(n_6040),
.B(n_6021),
.Y(n_8293)
);

NAND2x1p5_ASAP7_75t_L g8294 ( 
.A(n_7061),
.B(n_5884),
.Y(n_8294)
);

AOI21xp33_ASAP7_75t_SL g8295 ( 
.A1(n_6705),
.A2(n_5952),
.B(n_5897),
.Y(n_8295)
);

NOR2xp33_ASAP7_75t_L g8296 ( 
.A(n_7019),
.B(n_6077),
.Y(n_8296)
);

INVx1_ASAP7_75t_L g8297 ( 
.A(n_7340),
.Y(n_8297)
);

INVx1_ASAP7_75t_L g8298 ( 
.A(n_7353),
.Y(n_8298)
);

BUFx2_ASAP7_75t_L g8299 ( 
.A(n_7278),
.Y(n_8299)
);

HB1xp67_ASAP7_75t_L g8300 ( 
.A(n_7388),
.Y(n_8300)
);

INVx2_ASAP7_75t_L g8301 ( 
.A(n_7131),
.Y(n_8301)
);

INVx2_ASAP7_75t_SL g8302 ( 
.A(n_7042),
.Y(n_8302)
);

INVx1_ASAP7_75t_L g8303 ( 
.A(n_7353),
.Y(n_8303)
);

CKINVDCx11_ASAP7_75t_R g8304 ( 
.A(n_7042),
.Y(n_8304)
);

INVx2_ASAP7_75t_L g8305 ( 
.A(n_7131),
.Y(n_8305)
);

INVx1_ASAP7_75t_SL g8306 ( 
.A(n_7191),
.Y(n_8306)
);

AOI22xp33_ASAP7_75t_L g8307 ( 
.A1(n_6877),
.A2(n_5995),
.B1(n_6087),
.B2(n_4865),
.Y(n_8307)
);

INVx1_ASAP7_75t_L g8308 ( 
.A(n_7369),
.Y(n_8308)
);

INVx1_ASAP7_75t_L g8309 ( 
.A(n_7369),
.Y(n_8309)
);

INVx1_ASAP7_75t_L g8310 ( 
.A(n_7380),
.Y(n_8310)
);

AND2x2_ASAP7_75t_L g8311 ( 
.A(n_6620),
.B(n_6639),
.Y(n_8311)
);

INVx1_ASAP7_75t_L g8312 ( 
.A(n_7380),
.Y(n_8312)
);

INVx1_ASAP7_75t_L g8313 ( 
.A(n_7383),
.Y(n_8313)
);

OAI21x1_ASAP7_75t_L g8314 ( 
.A1(n_6983),
.A2(n_6040),
.B(n_6021),
.Y(n_8314)
);

OAI21x1_ASAP7_75t_L g8315 ( 
.A1(n_7154),
.A2(n_7180),
.B(n_7096),
.Y(n_8315)
);

INVx2_ASAP7_75t_L g8316 ( 
.A(n_7131),
.Y(n_8316)
);

INVx1_ASAP7_75t_L g8317 ( 
.A(n_7383),
.Y(n_8317)
);

INVx2_ASAP7_75t_L g8318 ( 
.A(n_7249),
.Y(n_8318)
);

AOI22xp33_ASAP7_75t_SL g8319 ( 
.A1(n_6500),
.A2(n_6510),
.B1(n_6825),
.B2(n_7061),
.Y(n_8319)
);

INVx1_ASAP7_75t_L g8320 ( 
.A(n_7391),
.Y(n_8320)
);

INVx1_ASAP7_75t_L g8321 ( 
.A(n_7391),
.Y(n_8321)
);

HB1xp67_ASAP7_75t_L g8322 ( 
.A(n_7372),
.Y(n_8322)
);

BUFx2_ASAP7_75t_L g8323 ( 
.A(n_7315),
.Y(n_8323)
);

INVx1_ASAP7_75t_L g8324 ( 
.A(n_7394),
.Y(n_8324)
);

INVx2_ASAP7_75t_L g8325 ( 
.A(n_7349),
.Y(n_8325)
);

INVx1_ASAP7_75t_L g8326 ( 
.A(n_7394),
.Y(n_8326)
);

INVx1_ASAP7_75t_L g8327 ( 
.A(n_7396),
.Y(n_8327)
);

OAI22xp5_ASAP7_75t_L g8328 ( 
.A1(n_6599),
.A2(n_6303),
.B1(n_6373),
.B2(n_6313),
.Y(n_8328)
);

AO21x2_ASAP7_75t_L g8329 ( 
.A1(n_6526),
.A2(n_6839),
.B(n_6474),
.Y(n_8329)
);

INVx1_ASAP7_75t_L g8330 ( 
.A(n_7396),
.Y(n_8330)
);

INVx1_ASAP7_75t_L g8331 ( 
.A(n_7405),
.Y(n_8331)
);

BUFx2_ASAP7_75t_R g8332 ( 
.A(n_7196),
.Y(n_8332)
);

NAND2x1p5_ASAP7_75t_L g8333 ( 
.A(n_7237),
.B(n_5884),
.Y(n_8333)
);

AOI21x1_ASAP7_75t_L g8334 ( 
.A1(n_7106),
.A2(n_6411),
.B(n_6409),
.Y(n_8334)
);

INVx1_ASAP7_75t_L g8335 ( 
.A(n_7405),
.Y(n_8335)
);

INVx1_ASAP7_75t_SL g8336 ( 
.A(n_7191),
.Y(n_8336)
);

AO21x2_ASAP7_75t_L g8337 ( 
.A1(n_6526),
.A2(n_5796),
.B(n_5782),
.Y(n_8337)
);

CKINVDCx20_ASAP7_75t_R g8338 ( 
.A(n_7381),
.Y(n_8338)
);

AOI22xp33_ASAP7_75t_L g8339 ( 
.A1(n_6877),
.A2(n_5995),
.B1(n_6087),
.B2(n_4865),
.Y(n_8339)
);

INVx2_ASAP7_75t_SL g8340 ( 
.A(n_7042),
.Y(n_8340)
);

BUFx2_ASAP7_75t_L g8341 ( 
.A(n_7315),
.Y(n_8341)
);

INVx1_ASAP7_75t_L g8342 ( 
.A(n_7160),
.Y(n_8342)
);

NOR2xp33_ASAP7_75t_L g8343 ( 
.A(n_7063),
.B(n_6198),
.Y(n_8343)
);

AOI21x1_ASAP7_75t_L g8344 ( 
.A1(n_7106),
.A2(n_6411),
.B(n_6409),
.Y(n_8344)
);

INVx1_ASAP7_75t_L g8345 ( 
.A(n_7160),
.Y(n_8345)
);

INVx1_ASAP7_75t_L g8346 ( 
.A(n_7173),
.Y(n_8346)
);

BUFx2_ASAP7_75t_R g8347 ( 
.A(n_7113),
.Y(n_8347)
);

INVx2_ASAP7_75t_L g8348 ( 
.A(n_7249),
.Y(n_8348)
);

AND2x2_ASAP7_75t_L g8349 ( 
.A(n_6620),
.B(n_6004),
.Y(n_8349)
);

INVx1_ASAP7_75t_L g8350 ( 
.A(n_7173),
.Y(n_8350)
);

BUFx2_ASAP7_75t_L g8351 ( 
.A(n_7126),
.Y(n_8351)
);

INVx1_ASAP7_75t_L g8352 ( 
.A(n_7174),
.Y(n_8352)
);

INVx1_ASAP7_75t_L g8353 ( 
.A(n_7174),
.Y(n_8353)
);

NAND2x1p5_ASAP7_75t_L g8354 ( 
.A(n_7371),
.B(n_5884),
.Y(n_8354)
);

AND2x2_ASAP7_75t_L g8355 ( 
.A(n_7433),
.B(n_6825),
.Y(n_8355)
);

OAI21x1_ASAP7_75t_L g8356 ( 
.A1(n_7423),
.A2(n_7180),
.B(n_6803),
.Y(n_8356)
);

HB1xp67_ASAP7_75t_L g8357 ( 
.A(n_7434),
.Y(n_8357)
);

INVx1_ASAP7_75t_L g8358 ( 
.A(n_7419),
.Y(n_8358)
);

BUFx4f_ASAP7_75t_L g8359 ( 
.A(n_7449),
.Y(n_8359)
);

INVx1_ASAP7_75t_L g8360 ( 
.A(n_7419),
.Y(n_8360)
);

AND2x2_ASAP7_75t_L g8361 ( 
.A(n_7433),
.B(n_6825),
.Y(n_8361)
);

INVx1_ASAP7_75t_L g8362 ( 
.A(n_7478),
.Y(n_8362)
);

INVx1_ASAP7_75t_L g8363 ( 
.A(n_7478),
.Y(n_8363)
);

INVx1_ASAP7_75t_L g8364 ( 
.A(n_7583),
.Y(n_8364)
);

OAI21x1_ASAP7_75t_L g8365 ( 
.A1(n_7423),
.A2(n_7489),
.B(n_7457),
.Y(n_8365)
);

AND2x2_ASAP7_75t_L g8366 ( 
.A(n_7463),
.B(n_6825),
.Y(n_8366)
);

OA21x2_ASAP7_75t_L g8367 ( 
.A1(n_7421),
.A2(n_7444),
.B(n_7979),
.Y(n_8367)
);

AOI221xp5_ASAP7_75t_L g8368 ( 
.A1(n_7416),
.A2(n_6567),
.B1(n_6664),
.B2(n_7167),
.C(n_7006),
.Y(n_8368)
);

AOI222xp33_ASAP7_75t_L g8369 ( 
.A1(n_7416),
.A2(n_7007),
.B1(n_7001),
.B2(n_7167),
.C1(n_6968),
.C2(n_6672),
.Y(n_8369)
);

INVx1_ASAP7_75t_L g8370 ( 
.A(n_7440),
.Y(n_8370)
);

AND2x2_ASAP7_75t_L g8371 ( 
.A(n_7463),
.B(n_6825),
.Y(n_8371)
);

INVx3_ASAP7_75t_L g8372 ( 
.A(n_7758),
.Y(n_8372)
);

INVx2_ASAP7_75t_L g8373 ( 
.A(n_7423),
.Y(n_8373)
);

INVx1_ASAP7_75t_L g8374 ( 
.A(n_7440),
.Y(n_8374)
);

INVx2_ASAP7_75t_L g8375 ( 
.A(n_7423),
.Y(n_8375)
);

HB1xp67_ASAP7_75t_L g8376 ( 
.A(n_7446),
.Y(n_8376)
);

INVxp67_ASAP7_75t_L g8377 ( 
.A(n_7803),
.Y(n_8377)
);

BUFx3_ASAP7_75t_L g8378 ( 
.A(n_7474),
.Y(n_8378)
);

OAI21x1_ASAP7_75t_L g8379 ( 
.A1(n_7457),
.A2(n_7510),
.B(n_7489),
.Y(n_8379)
);

INVx1_ASAP7_75t_L g8380 ( 
.A(n_7442),
.Y(n_8380)
);

CKINVDCx20_ASAP7_75t_R g8381 ( 
.A(n_7413),
.Y(n_8381)
);

INVx1_ASAP7_75t_L g8382 ( 
.A(n_7443),
.Y(n_8382)
);

BUFx3_ASAP7_75t_L g8383 ( 
.A(n_7474),
.Y(n_8383)
);

INVx2_ASAP7_75t_L g8384 ( 
.A(n_7457),
.Y(n_8384)
);

INVx2_ASAP7_75t_L g8385 ( 
.A(n_7457),
.Y(n_8385)
);

HB1xp67_ASAP7_75t_L g8386 ( 
.A(n_8080),
.Y(n_8386)
);

BUFx3_ASAP7_75t_L g8387 ( 
.A(n_7684),
.Y(n_8387)
);

INVx1_ASAP7_75t_L g8388 ( 
.A(n_7443),
.Y(n_8388)
);

NAND2xp5_ASAP7_75t_L g8389 ( 
.A(n_7618),
.B(n_6552),
.Y(n_8389)
);

INVx1_ASAP7_75t_L g8390 ( 
.A(n_7453),
.Y(n_8390)
);

INVx2_ASAP7_75t_L g8391 ( 
.A(n_7510),
.Y(n_8391)
);

AOI21x1_ASAP7_75t_L g8392 ( 
.A1(n_7469),
.A2(n_7202),
.B(n_7126),
.Y(n_8392)
);

INVx2_ASAP7_75t_SL g8393 ( 
.A(n_7449),
.Y(n_8393)
);

INVx1_ASAP7_75t_L g8394 ( 
.A(n_7453),
.Y(n_8394)
);

INVx1_ASAP7_75t_L g8395 ( 
.A(n_7530),
.Y(n_8395)
);

INVx1_ASAP7_75t_L g8396 ( 
.A(n_7530),
.Y(n_8396)
);

BUFx3_ASAP7_75t_L g8397 ( 
.A(n_7521),
.Y(n_8397)
);

INVx2_ASAP7_75t_L g8398 ( 
.A(n_7489),
.Y(n_8398)
);

OA21x2_ASAP7_75t_L g8399 ( 
.A1(n_7444),
.A2(n_6526),
.B(n_6486),
.Y(n_8399)
);

INVx2_ASAP7_75t_L g8400 ( 
.A(n_7489),
.Y(n_8400)
);

AND2x2_ASAP7_75t_L g8401 ( 
.A(n_7630),
.B(n_7202),
.Y(n_8401)
);

AOI22xp33_ASAP7_75t_L g8402 ( 
.A1(n_7472),
.A2(n_6567),
.B1(n_6500),
.B2(n_6510),
.Y(n_8402)
);

INVx1_ASAP7_75t_L g8403 ( 
.A(n_7465),
.Y(n_8403)
);

INVx1_ASAP7_75t_L g8404 ( 
.A(n_7465),
.Y(n_8404)
);

INVx1_ASAP7_75t_L g8405 ( 
.A(n_7484),
.Y(n_8405)
);

INVx1_ASAP7_75t_L g8406 ( 
.A(n_7484),
.Y(n_8406)
);

BUFx3_ASAP7_75t_L g8407 ( 
.A(n_7521),
.Y(n_8407)
);

AND2x2_ASAP7_75t_L g8408 ( 
.A(n_7630),
.B(n_7202),
.Y(n_8408)
);

INVx1_ASAP7_75t_L g8409 ( 
.A(n_7518),
.Y(n_8409)
);

INVx2_ASAP7_75t_L g8410 ( 
.A(n_7526),
.Y(n_8410)
);

OR2x6_ASAP7_75t_L g8411 ( 
.A(n_8164),
.B(n_7824),
.Y(n_8411)
);

INVx1_ASAP7_75t_L g8412 ( 
.A(n_7518),
.Y(n_8412)
);

INVx2_ASAP7_75t_L g8413 ( 
.A(n_7526),
.Y(n_8413)
);

OR2x2_ASAP7_75t_L g8414 ( 
.A(n_7687),
.B(n_7054),
.Y(n_8414)
);

INVx1_ASAP7_75t_L g8415 ( 
.A(n_7528),
.Y(n_8415)
);

AOI22xp33_ASAP7_75t_SL g8416 ( 
.A1(n_7472),
.A2(n_6510),
.B1(n_6500),
.B2(n_6443),
.Y(n_8416)
);

OAI22xp5_ASAP7_75t_L g8417 ( 
.A1(n_7435),
.A2(n_6927),
.B1(n_7309),
.B2(n_6830),
.Y(n_8417)
);

INVx1_ASAP7_75t_L g8418 ( 
.A(n_7456),
.Y(n_8418)
);

OAI21x1_ASAP7_75t_L g8419 ( 
.A1(n_7510),
.A2(n_7526),
.B(n_7758),
.Y(n_8419)
);

INVx2_ASAP7_75t_L g8420 ( 
.A(n_7510),
.Y(n_8420)
);

INVx2_ASAP7_75t_L g8421 ( 
.A(n_7526),
.Y(n_8421)
);

INVx2_ASAP7_75t_L g8422 ( 
.A(n_7635),
.Y(n_8422)
);

INVx2_ASAP7_75t_L g8423 ( 
.A(n_7635),
.Y(n_8423)
);

INVx1_ASAP7_75t_L g8424 ( 
.A(n_7456),
.Y(n_8424)
);

INVx2_ASAP7_75t_L g8425 ( 
.A(n_7635),
.Y(n_8425)
);

OAI22xp33_ASAP7_75t_L g8426 ( 
.A1(n_7509),
.A2(n_6596),
.B1(n_6715),
.B2(n_7007),
.Y(n_8426)
);

NAND2xp5_ASAP7_75t_L g8427 ( 
.A(n_7618),
.B(n_6552),
.Y(n_8427)
);

AND2x4_ASAP7_75t_L g8428 ( 
.A(n_8133),
.B(n_7164),
.Y(n_8428)
);

BUFx6f_ASAP7_75t_L g8429 ( 
.A(n_7412),
.Y(n_8429)
);

OAI22xp5_ASAP7_75t_L g8430 ( 
.A1(n_7506),
.A2(n_6927),
.B1(n_7309),
.B2(n_7159),
.Y(n_8430)
);

AND2x2_ASAP7_75t_L g8431 ( 
.A(n_7641),
.B(n_6639),
.Y(n_8431)
);

OR2x2_ASAP7_75t_L g8432 ( 
.A(n_7687),
.B(n_7054),
.Y(n_8432)
);

INVx1_ASAP7_75t_L g8433 ( 
.A(n_7583),
.Y(n_8433)
);

INVx1_ASAP7_75t_L g8434 ( 
.A(n_7716),
.Y(n_8434)
);

HB1xp67_ASAP7_75t_L g8435 ( 
.A(n_8281),
.Y(n_8435)
);

INVx1_ASAP7_75t_L g8436 ( 
.A(n_7716),
.Y(n_8436)
);

INVx1_ASAP7_75t_L g8437 ( 
.A(n_7821),
.Y(n_8437)
);

INVx1_ASAP7_75t_L g8438 ( 
.A(n_7821),
.Y(n_8438)
);

OAI21x1_ASAP7_75t_L g8439 ( 
.A1(n_7758),
.A2(n_6876),
.B(n_6656),
.Y(n_8439)
);

INVx1_ASAP7_75t_L g8440 ( 
.A(n_7822),
.Y(n_8440)
);

AOI22xp33_ASAP7_75t_L g8441 ( 
.A1(n_7509),
.A2(n_6510),
.B1(n_6839),
.B2(n_6596),
.Y(n_8441)
);

OAI22xp5_ASAP7_75t_L g8442 ( 
.A1(n_7525),
.A2(n_7159),
.B1(n_6657),
.B2(n_6949),
.Y(n_8442)
);

INVx2_ASAP7_75t_SL g8443 ( 
.A(n_7449),
.Y(n_8443)
);

INVx2_ASAP7_75t_L g8444 ( 
.A(n_7635),
.Y(n_8444)
);

INVx1_ASAP7_75t_L g8445 ( 
.A(n_7593),
.Y(n_8445)
);

AND2x2_ASAP7_75t_L g8446 ( 
.A(n_7641),
.B(n_6639),
.Y(n_8446)
);

OR2x6_ASAP7_75t_L g8447 ( 
.A(n_8164),
.B(n_7057),
.Y(n_8447)
);

NAND2xp5_ASAP7_75t_L g8448 ( 
.A(n_7689),
.B(n_6558),
.Y(n_8448)
);

INVx3_ASAP7_75t_L g8449 ( 
.A(n_7758),
.Y(n_8449)
);

HB1xp67_ASAP7_75t_L g8450 ( 
.A(n_8306),
.Y(n_8450)
);

AND2x2_ASAP7_75t_L g8451 ( 
.A(n_7678),
.B(n_7573),
.Y(n_8451)
);

BUFx2_ASAP7_75t_L g8452 ( 
.A(n_7803),
.Y(n_8452)
);

BUFx3_ASAP7_75t_L g8453 ( 
.A(n_7846),
.Y(n_8453)
);

HB1xp67_ASAP7_75t_L g8454 ( 
.A(n_8336),
.Y(n_8454)
);

BUFx3_ASAP7_75t_L g8455 ( 
.A(n_7740),
.Y(n_8455)
);

INVx3_ASAP7_75t_L g8456 ( 
.A(n_7766),
.Y(n_8456)
);

AO21x1_ASAP7_75t_L g8457 ( 
.A1(n_7735),
.A2(n_6664),
.B(n_7015),
.Y(n_8457)
);

INVx2_ASAP7_75t_L g8458 ( 
.A(n_7640),
.Y(n_8458)
);

INVx2_ASAP7_75t_L g8459 ( 
.A(n_7640),
.Y(n_8459)
);

AND2x2_ASAP7_75t_L g8460 ( 
.A(n_7678),
.B(n_6737),
.Y(n_8460)
);

BUFx2_ASAP7_75t_L g8461 ( 
.A(n_7412),
.Y(n_8461)
);

INVx2_ASAP7_75t_SL g8462 ( 
.A(n_7449),
.Y(n_8462)
);

INVx1_ASAP7_75t_L g8463 ( 
.A(n_7593),
.Y(n_8463)
);

INVx1_ASAP7_75t_L g8464 ( 
.A(n_7602),
.Y(n_8464)
);

NAND2xp5_ASAP7_75t_L g8465 ( 
.A(n_7689),
.B(n_6558),
.Y(n_8465)
);

INVx1_ASAP7_75t_L g8466 ( 
.A(n_7602),
.Y(n_8466)
);

INVx3_ASAP7_75t_L g8467 ( 
.A(n_7766),
.Y(n_8467)
);

INVx2_ASAP7_75t_L g8468 ( 
.A(n_7640),
.Y(n_8468)
);

INVx1_ASAP7_75t_L g8469 ( 
.A(n_7603),
.Y(n_8469)
);

CKINVDCx9p33_ASAP7_75t_R g8470 ( 
.A(n_7742),
.Y(n_8470)
);

AND2x2_ASAP7_75t_L g8471 ( 
.A(n_7573),
.B(n_6737),
.Y(n_8471)
);

INVx1_ASAP7_75t_L g8472 ( 
.A(n_7417),
.Y(n_8472)
);

INVx1_ASAP7_75t_L g8473 ( 
.A(n_7417),
.Y(n_8473)
);

INVx1_ASAP7_75t_L g8474 ( 
.A(n_7425),
.Y(n_8474)
);

INVx3_ASAP7_75t_L g8475 ( 
.A(n_7766),
.Y(n_8475)
);

HB1xp67_ASAP7_75t_L g8476 ( 
.A(n_8322),
.Y(n_8476)
);

OA21x2_ASAP7_75t_L g8477 ( 
.A1(n_7825),
.A2(n_6486),
.B(n_6483),
.Y(n_8477)
);

OAI21xp5_ASAP7_75t_L g8478 ( 
.A1(n_7801),
.A2(n_6772),
.B(n_6717),
.Y(n_8478)
);

OAI21x1_ASAP7_75t_L g8479 ( 
.A1(n_7766),
.A2(n_6876),
.B(n_6656),
.Y(n_8479)
);

OAI21x1_ASAP7_75t_L g8480 ( 
.A1(n_7786),
.A2(n_7129),
.B(n_6522),
.Y(n_8480)
);

OAI21x1_ASAP7_75t_L g8481 ( 
.A1(n_7786),
.A2(n_7129),
.B(n_6522),
.Y(n_8481)
);

BUFx12f_ASAP7_75t_L g8482 ( 
.A(n_7932),
.Y(n_8482)
);

INVx2_ASAP7_75t_SL g8483 ( 
.A(n_7449),
.Y(n_8483)
);

AND2x4_ASAP7_75t_L g8484 ( 
.A(n_8133),
.B(n_7164),
.Y(n_8484)
);

INVx1_ASAP7_75t_L g8485 ( 
.A(n_7425),
.Y(n_8485)
);

NOR2xp33_ASAP7_75t_L g8486 ( 
.A(n_7571),
.B(n_6001),
.Y(n_8486)
);

CKINVDCx9p33_ASAP7_75t_R g8487 ( 
.A(n_7694),
.Y(n_8487)
);

INVx1_ASAP7_75t_L g8488 ( 
.A(n_7580),
.Y(n_8488)
);

INVxp67_ASAP7_75t_L g8489 ( 
.A(n_8228),
.Y(n_8489)
);

INVx2_ASAP7_75t_L g8490 ( 
.A(n_7640),
.Y(n_8490)
);

BUFx3_ASAP7_75t_L g8491 ( 
.A(n_7696),
.Y(n_8491)
);

BUFx6f_ASAP7_75t_L g8492 ( 
.A(n_7412),
.Y(n_8492)
);

AOI221xp5_ASAP7_75t_L g8493 ( 
.A1(n_7525),
.A2(n_7006),
.B1(n_7015),
.B2(n_7026),
.C(n_6968),
.Y(n_8493)
);

INVx2_ASAP7_75t_L g8494 ( 
.A(n_7644),
.Y(n_8494)
);

OAI21xp33_ASAP7_75t_SL g8495 ( 
.A1(n_7937),
.A2(n_6947),
.B(n_6750),
.Y(n_8495)
);

AND2x2_ASAP7_75t_L g8496 ( 
.A(n_7468),
.B(n_6737),
.Y(n_8496)
);

INVx1_ASAP7_75t_L g8497 ( 
.A(n_7500),
.Y(n_8497)
);

INVx1_ASAP7_75t_L g8498 ( 
.A(n_7500),
.Y(n_8498)
);

INVx2_ASAP7_75t_L g8499 ( 
.A(n_7644),
.Y(n_8499)
);

INVx1_ASAP7_75t_L g8500 ( 
.A(n_7565),
.Y(n_8500)
);

INVx2_ASAP7_75t_L g8501 ( 
.A(n_7644),
.Y(n_8501)
);

INVx2_ASAP7_75t_L g8502 ( 
.A(n_7644),
.Y(n_8502)
);

INVx2_ASAP7_75t_L g8503 ( 
.A(n_7655),
.Y(n_8503)
);

INVx2_ASAP7_75t_L g8504 ( 
.A(n_7655),
.Y(n_8504)
);

NAND2x1_ASAP7_75t_L g8505 ( 
.A(n_7485),
.B(n_6573),
.Y(n_8505)
);

INVx1_ASAP7_75t_L g8506 ( 
.A(n_7565),
.Y(n_8506)
);

BUFx2_ASAP7_75t_L g8507 ( 
.A(n_7415),
.Y(n_8507)
);

AND2x4_ASAP7_75t_L g8508 ( 
.A(n_8133),
.B(n_7164),
.Y(n_8508)
);

INVx2_ASAP7_75t_L g8509 ( 
.A(n_7655),
.Y(n_8509)
);

AND2x2_ASAP7_75t_L g8510 ( 
.A(n_7468),
.B(n_6750),
.Y(n_8510)
);

INVx1_ASAP7_75t_L g8511 ( 
.A(n_7513),
.Y(n_8511)
);

INVx1_ASAP7_75t_L g8512 ( 
.A(n_7513),
.Y(n_8512)
);

NAND2xp5_ASAP7_75t_L g8513 ( 
.A(n_7445),
.B(n_6609),
.Y(n_8513)
);

BUFx4f_ASAP7_75t_SL g8514 ( 
.A(n_7619),
.Y(n_8514)
);

INVx1_ASAP7_75t_L g8515 ( 
.A(n_7451),
.Y(n_8515)
);

INVx3_ASAP7_75t_L g8516 ( 
.A(n_7786),
.Y(n_8516)
);

OR2x2_ASAP7_75t_L g8517 ( 
.A(n_7815),
.B(n_6666),
.Y(n_8517)
);

INVx1_ASAP7_75t_L g8518 ( 
.A(n_7451),
.Y(n_8518)
);

INVx2_ASAP7_75t_L g8519 ( 
.A(n_7655),
.Y(n_8519)
);

AND2x2_ASAP7_75t_L g8520 ( 
.A(n_7563),
.B(n_7424),
.Y(n_8520)
);

AO32x2_ASAP7_75t_L g8521 ( 
.A1(n_8239),
.A2(n_7002),
.A3(n_8095),
.B1(n_7553),
.B2(n_7616),
.Y(n_8521)
);

INVx1_ASAP7_75t_L g8522 ( 
.A(n_7528),
.Y(n_8522)
);

INVx2_ASAP7_75t_L g8523 ( 
.A(n_7741),
.Y(n_8523)
);

INVx3_ASAP7_75t_L g8524 ( 
.A(n_7786),
.Y(n_8524)
);

INVx2_ASAP7_75t_L g8525 ( 
.A(n_7741),
.Y(n_8525)
);

INVx1_ASAP7_75t_L g8526 ( 
.A(n_7572),
.Y(n_8526)
);

INVx1_ASAP7_75t_L g8527 ( 
.A(n_7572),
.Y(n_8527)
);

INVx1_ASAP7_75t_L g8528 ( 
.A(n_7574),
.Y(n_8528)
);

INVx1_ASAP7_75t_L g8529 ( 
.A(n_7574),
.Y(n_8529)
);

INVx2_ASAP7_75t_SL g8530 ( 
.A(n_7449),
.Y(n_8530)
);

INVx2_ASAP7_75t_L g8531 ( 
.A(n_7741),
.Y(n_8531)
);

INVx2_ASAP7_75t_SL g8532 ( 
.A(n_7738),
.Y(n_8532)
);

INVx2_ASAP7_75t_L g8533 ( 
.A(n_7741),
.Y(n_8533)
);

INVx1_ASAP7_75t_L g8534 ( 
.A(n_7539),
.Y(n_8534)
);

OA21x2_ASAP7_75t_L g8535 ( 
.A1(n_7825),
.A2(n_6486),
.B(n_6483),
.Y(n_8535)
);

AO21x2_ASAP7_75t_L g8536 ( 
.A1(n_8329),
.A2(n_6839),
.B(n_6550),
.Y(n_8536)
);

HB1xp67_ASAP7_75t_L g8537 ( 
.A(n_7499),
.Y(n_8537)
);

NAND2xp5_ASAP7_75t_L g8538 ( 
.A(n_8064),
.B(n_6609),
.Y(n_8538)
);

INVx2_ASAP7_75t_L g8539 ( 
.A(n_7895),
.Y(n_8539)
);

BUFx3_ASAP7_75t_L g8540 ( 
.A(n_7985),
.Y(n_8540)
);

OA21x2_ASAP7_75t_L g8541 ( 
.A1(n_7725),
.A2(n_6483),
.B(n_6527),
.Y(n_8541)
);

INVx2_ASAP7_75t_L g8542 ( 
.A(n_7895),
.Y(n_8542)
);

INVx2_ASAP7_75t_L g8543 ( 
.A(n_7895),
.Y(n_8543)
);

OAI22xp5_ASAP7_75t_L g8544 ( 
.A1(n_7543),
.A2(n_6657),
.B1(n_6949),
.B2(n_6756),
.Y(n_8544)
);

INVx2_ASAP7_75t_L g8545 ( 
.A(n_7895),
.Y(n_8545)
);

INVx1_ASAP7_75t_L g8546 ( 
.A(n_7556),
.Y(n_8546)
);

AOI22xp33_ASAP7_75t_SL g8547 ( 
.A1(n_7543),
.A2(n_6510),
.B1(n_6443),
.B2(n_6770),
.Y(n_8547)
);

INVx2_ASAP7_75t_L g8548 ( 
.A(n_7916),
.Y(n_8548)
);

INVx1_ASAP7_75t_L g8549 ( 
.A(n_7613),
.Y(n_8549)
);

INVx1_ASAP7_75t_L g8550 ( 
.A(n_7613),
.Y(n_8550)
);

OAI21x1_ASAP7_75t_L g8551 ( 
.A1(n_7916),
.A2(n_6522),
.B(n_6511),
.Y(n_8551)
);

INVx1_ASAP7_75t_L g8552 ( 
.A(n_7653),
.Y(n_8552)
);

NOR2xp33_ASAP7_75t_L g8553 ( 
.A(n_7733),
.B(n_6397),
.Y(n_8553)
);

INVx2_ASAP7_75t_L g8554 ( 
.A(n_7916),
.Y(n_8554)
);

INVx1_ASAP7_75t_L g8555 ( 
.A(n_7653),
.Y(n_8555)
);

OAI22xp5_ASAP7_75t_L g8556 ( 
.A1(n_7560),
.A2(n_6756),
.B1(n_6745),
.B2(n_6859),
.Y(n_8556)
);

INVx3_ASAP7_75t_L g8557 ( 
.A(n_7916),
.Y(n_8557)
);

NAND2x1p5_ASAP7_75t_L g8558 ( 
.A(n_7874),
.B(n_7057),
.Y(n_8558)
);

INVx1_ASAP7_75t_L g8559 ( 
.A(n_7671),
.Y(n_8559)
);

HB1xp67_ASAP7_75t_L g8560 ( 
.A(n_7522),
.Y(n_8560)
);

INVx3_ASAP7_75t_L g8561 ( 
.A(n_7934),
.Y(n_8561)
);

NAND2xp33_ASAP7_75t_SL g8562 ( 
.A(n_7560),
.B(n_7381),
.Y(n_8562)
);

OR2x6_ASAP7_75t_L g8563 ( 
.A(n_8164),
.B(n_7057),
.Y(n_8563)
);

INVx2_ASAP7_75t_L g8564 ( 
.A(n_7934),
.Y(n_8564)
);

INVx2_ASAP7_75t_L g8565 ( 
.A(n_7934),
.Y(n_8565)
);

BUFx6f_ASAP7_75t_L g8566 ( 
.A(n_7415),
.Y(n_8566)
);

INVx1_ASAP7_75t_SL g8567 ( 
.A(n_7515),
.Y(n_8567)
);

INVx2_ASAP7_75t_L g8568 ( 
.A(n_7934),
.Y(n_8568)
);

INVx1_ASAP7_75t_L g8569 ( 
.A(n_7590),
.Y(n_8569)
);

AND2x4_ASAP7_75t_L g8570 ( 
.A(n_8133),
.B(n_7164),
.Y(n_8570)
);

CKINVDCx6p67_ASAP7_75t_R g8571 ( 
.A(n_7415),
.Y(n_8571)
);

HB1xp67_ASAP7_75t_L g8572 ( 
.A(n_7533),
.Y(n_8572)
);

INVx1_ASAP7_75t_L g8573 ( 
.A(n_7523),
.Y(n_8573)
);

INVx3_ASAP7_75t_L g8574 ( 
.A(n_7968),
.Y(n_8574)
);

INVx1_ASAP7_75t_L g8575 ( 
.A(n_7523),
.Y(n_8575)
);

INVx2_ASAP7_75t_L g8576 ( 
.A(n_7968),
.Y(n_8576)
);

INVx2_ASAP7_75t_L g8577 ( 
.A(n_7968),
.Y(n_8577)
);

INVx2_ASAP7_75t_L g8578 ( 
.A(n_7968),
.Y(n_8578)
);

INVx2_ASAP7_75t_L g8579 ( 
.A(n_7978),
.Y(n_8579)
);

INVx3_ASAP7_75t_L g8580 ( 
.A(n_7978),
.Y(n_8580)
);

BUFx2_ASAP7_75t_L g8581 ( 
.A(n_7418),
.Y(n_8581)
);

INVx1_ASAP7_75t_L g8582 ( 
.A(n_7603),
.Y(n_8582)
);

INVx1_ASAP7_75t_L g8583 ( 
.A(n_7755),
.Y(n_8583)
);

INVx1_ASAP7_75t_L g8584 ( 
.A(n_7755),
.Y(n_8584)
);

OAI21x1_ASAP7_75t_L g8585 ( 
.A1(n_7978),
.A2(n_6511),
.B(n_6650),
.Y(n_8585)
);

A2O1A1Ixp33_ASAP7_75t_L g8586 ( 
.A1(n_7645),
.A2(n_7657),
.B(n_7673),
.C(n_8079),
.Y(n_8586)
);

OAI21x1_ASAP7_75t_L g8587 ( 
.A1(n_7978),
.A2(n_6511),
.B(n_6650),
.Y(n_8587)
);

OA21x2_ASAP7_75t_L g8588 ( 
.A1(n_7591),
.A2(n_7719),
.B(n_7718),
.Y(n_8588)
);

INVx2_ASAP7_75t_L g8589 ( 
.A(n_8077),
.Y(n_8589)
);

INVx2_ASAP7_75t_L g8590 ( 
.A(n_8077),
.Y(n_8590)
);

NOR2xp33_ASAP7_75t_L g8591 ( 
.A(n_7462),
.B(n_6397),
.Y(n_8591)
);

NAND2xp5_ASAP7_75t_L g8592 ( 
.A(n_7645),
.B(n_6637),
.Y(n_8592)
);

INVx1_ASAP7_75t_L g8593 ( 
.A(n_7671),
.Y(n_8593)
);

INVx2_ASAP7_75t_L g8594 ( 
.A(n_8077),
.Y(n_8594)
);

BUFx3_ASAP7_75t_L g8595 ( 
.A(n_7418),
.Y(n_8595)
);

INVx1_ASAP7_75t_L g8596 ( 
.A(n_7728),
.Y(n_8596)
);

INVx1_ASAP7_75t_L g8597 ( 
.A(n_7728),
.Y(n_8597)
);

NAND2xp5_ASAP7_75t_L g8598 ( 
.A(n_7657),
.B(n_6637),
.Y(n_8598)
);

INVx1_ASAP7_75t_L g8599 ( 
.A(n_7787),
.Y(n_8599)
);

AO31x2_ASAP7_75t_L g8600 ( 
.A1(n_7673),
.A2(n_6968),
.A3(n_6977),
.B(n_6672),
.Y(n_8600)
);

INVx1_ASAP7_75t_SL g8601 ( 
.A(n_7552),
.Y(n_8601)
);

AOI21x1_ASAP7_75t_L g8602 ( 
.A1(n_7469),
.A2(n_6977),
.B(n_6672),
.Y(n_8602)
);

AND2x4_ASAP7_75t_L g8603 ( 
.A(n_8063),
.B(n_7164),
.Y(n_8603)
);

INVx1_ASAP7_75t_L g8604 ( 
.A(n_7547),
.Y(n_8604)
);

AOI22xp5_ASAP7_75t_L g8605 ( 
.A1(n_7651),
.A2(n_6715),
.B1(n_7303),
.B2(n_6718),
.Y(n_8605)
);

INVx1_ASAP7_75t_L g8606 ( 
.A(n_7547),
.Y(n_8606)
);

INVx2_ASAP7_75t_L g8607 ( 
.A(n_8077),
.Y(n_8607)
);

OAI21x1_ASAP7_75t_L g8608 ( 
.A1(n_8085),
.A2(n_7329),
.B(n_7257),
.Y(n_8608)
);

INVx2_ASAP7_75t_L g8609 ( 
.A(n_8085),
.Y(n_8609)
);

NAND2xp5_ASAP7_75t_L g8610 ( 
.A(n_8155),
.B(n_7184),
.Y(n_8610)
);

INVx1_ASAP7_75t_L g8611 ( 
.A(n_7441),
.Y(n_8611)
);

INVx1_ASAP7_75t_L g8612 ( 
.A(n_7441),
.Y(n_8612)
);

INVx1_ASAP7_75t_L g8613 ( 
.A(n_7442),
.Y(n_8613)
);

INVx1_ASAP7_75t_L g8614 ( 
.A(n_7539),
.Y(n_8614)
);

HB1xp67_ASAP7_75t_L g8615 ( 
.A(n_7540),
.Y(n_8615)
);

INVx1_ASAP7_75t_L g8616 ( 
.A(n_7550),
.Y(n_8616)
);

INVx2_ASAP7_75t_SL g8617 ( 
.A(n_7738),
.Y(n_8617)
);

INVx1_ASAP7_75t_SL g8618 ( 
.A(n_7570),
.Y(n_8618)
);

BUFx3_ASAP7_75t_L g8619 ( 
.A(n_7418),
.Y(n_8619)
);

OA21x2_ASAP7_75t_L g8620 ( 
.A1(n_7591),
.A2(n_6527),
.B(n_6472),
.Y(n_8620)
);

BUFx6f_ASAP7_75t_L g8621 ( 
.A(n_7438),
.Y(n_8621)
);

OAI21x1_ASAP7_75t_L g8622 ( 
.A1(n_8085),
.A2(n_7329),
.B(n_7257),
.Y(n_8622)
);

AND2x2_ASAP7_75t_L g8623 ( 
.A(n_7563),
.B(n_6750),
.Y(n_8623)
);

HB1xp67_ASAP7_75t_L g8624 ( 
.A(n_7586),
.Y(n_8624)
);

INVx2_ASAP7_75t_SL g8625 ( 
.A(n_7438),
.Y(n_8625)
);

OR2x2_ASAP7_75t_L g8626 ( 
.A(n_7815),
.B(n_6666),
.Y(n_8626)
);

HB1xp67_ASAP7_75t_L g8627 ( 
.A(n_7595),
.Y(n_8627)
);

INVx1_ASAP7_75t_L g8628 ( 
.A(n_7598),
.Y(n_8628)
);

BUFx3_ASAP7_75t_L g8629 ( 
.A(n_7438),
.Y(n_8629)
);

INVx1_ASAP7_75t_L g8630 ( 
.A(n_7589),
.Y(n_8630)
);

INVx1_ASAP7_75t_L g8631 ( 
.A(n_7589),
.Y(n_8631)
);

INVx2_ASAP7_75t_SL g8632 ( 
.A(n_7458),
.Y(n_8632)
);

OR2x2_ASAP7_75t_L g8633 ( 
.A(n_7414),
.B(n_6697),
.Y(n_8633)
);

INVx2_ASAP7_75t_L g8634 ( 
.A(n_8085),
.Y(n_8634)
);

AND2x2_ASAP7_75t_L g8635 ( 
.A(n_7424),
.B(n_6925),
.Y(n_8635)
);

INVx2_ASAP7_75t_L g8636 ( 
.A(n_7943),
.Y(n_8636)
);

INVx3_ASAP7_75t_L g8637 ( 
.A(n_7479),
.Y(n_8637)
);

AND2x2_ASAP7_75t_L g8638 ( 
.A(n_7814),
.B(n_6925),
.Y(n_8638)
);

INVx2_ASAP7_75t_L g8639 ( 
.A(n_7943),
.Y(n_8639)
);

BUFx2_ASAP7_75t_L g8640 ( 
.A(n_7462),
.Y(n_8640)
);

INVx2_ASAP7_75t_L g8641 ( 
.A(n_7945),
.Y(n_8641)
);

BUFx6f_ASAP7_75t_L g8642 ( 
.A(n_7462),
.Y(n_8642)
);

INVx3_ASAP7_75t_L g8643 ( 
.A(n_7479),
.Y(n_8643)
);

OAI21xp5_ASAP7_75t_L g8644 ( 
.A1(n_8079),
.A2(n_6772),
.B(n_6717),
.Y(n_8644)
);

OR2x2_ASAP7_75t_L g8645 ( 
.A(n_7414),
.B(n_6697),
.Y(n_8645)
);

INVx1_ASAP7_75t_L g8646 ( 
.A(n_7714),
.Y(n_8646)
);

BUFx6f_ASAP7_75t_L g8647 ( 
.A(n_7462),
.Y(n_8647)
);

OR2x2_ASAP7_75t_L g8648 ( 
.A(n_8277),
.B(n_6762),
.Y(n_8648)
);

CKINVDCx20_ASAP7_75t_R g8649 ( 
.A(n_7883),
.Y(n_8649)
);

INVx1_ASAP7_75t_L g8650 ( 
.A(n_7550),
.Y(n_8650)
);

INVx1_ASAP7_75t_L g8651 ( 
.A(n_7561),
.Y(n_8651)
);

INVx2_ASAP7_75t_L g8652 ( 
.A(n_7945),
.Y(n_8652)
);

OAI21x1_ASAP7_75t_L g8653 ( 
.A1(n_7538),
.A2(n_7046),
.B(n_6838),
.Y(n_8653)
);

BUFx2_ASAP7_75t_L g8654 ( 
.A(n_7600),
.Y(n_8654)
);

INVx1_ASAP7_75t_L g8655 ( 
.A(n_7561),
.Y(n_8655)
);

OR2x6_ASAP7_75t_L g8656 ( 
.A(n_7824),
.B(n_8333),
.Y(n_8656)
);

INVx2_ASAP7_75t_L g8657 ( 
.A(n_7949),
.Y(n_8657)
);

INVx2_ASAP7_75t_L g8658 ( 
.A(n_7949),
.Y(n_8658)
);

INVx2_ASAP7_75t_L g8659 ( 
.A(n_7953),
.Y(n_8659)
);

INVx2_ASAP7_75t_SL g8660 ( 
.A(n_7458),
.Y(n_8660)
);

INVx2_ASAP7_75t_L g8661 ( 
.A(n_7953),
.Y(n_8661)
);

OA21x2_ASAP7_75t_L g8662 ( 
.A1(n_7591),
.A2(n_6527),
.B(n_6472),
.Y(n_8662)
);

AND2x2_ASAP7_75t_L g8663 ( 
.A(n_7814),
.B(n_6925),
.Y(n_8663)
);

INVx1_ASAP7_75t_L g8664 ( 
.A(n_7610),
.Y(n_8664)
);

AOI21xp5_ASAP7_75t_L g8665 ( 
.A1(n_7713),
.A2(n_6515),
.B(n_6796),
.Y(n_8665)
);

INVx1_ASAP7_75t_L g8666 ( 
.A(n_7610),
.Y(n_8666)
);

INVx1_ASAP7_75t_L g8667 ( 
.A(n_7611),
.Y(n_8667)
);

CKINVDCx11_ASAP7_75t_R g8668 ( 
.A(n_8037),
.Y(n_8668)
);

INVx2_ASAP7_75t_SL g8669 ( 
.A(n_7535),
.Y(n_8669)
);

BUFx3_ASAP7_75t_L g8670 ( 
.A(n_7544),
.Y(n_8670)
);

INVx1_ASAP7_75t_L g8671 ( 
.A(n_7590),
.Y(n_8671)
);

INVx2_ASAP7_75t_L g8672 ( 
.A(n_7954),
.Y(n_8672)
);

AND2x2_ASAP7_75t_L g8673 ( 
.A(n_8028),
.B(n_7620),
.Y(n_8673)
);

INVx1_ASAP7_75t_L g8674 ( 
.A(n_7714),
.Y(n_8674)
);

BUFx2_ASAP7_75t_L g8675 ( 
.A(n_7600),
.Y(n_8675)
);

BUFx3_ASAP7_75t_L g8676 ( 
.A(n_7670),
.Y(n_8676)
);

OR2x2_ASAP7_75t_L g8677 ( 
.A(n_7542),
.B(n_6762),
.Y(n_8677)
);

HB1xp67_ASAP7_75t_L g8678 ( 
.A(n_7625),
.Y(n_8678)
);

INVx2_ASAP7_75t_SL g8679 ( 
.A(n_7535),
.Y(n_8679)
);

AND2x4_ASAP7_75t_L g8680 ( 
.A(n_8063),
.B(n_7164),
.Y(n_8680)
);

OAI21xp5_ASAP7_75t_L g8681 ( 
.A1(n_7948),
.A2(n_6718),
.B(n_6796),
.Y(n_8681)
);

AND2x2_ASAP7_75t_L g8682 ( 
.A(n_8028),
.B(n_7620),
.Y(n_8682)
);

AND2x2_ASAP7_75t_L g8683 ( 
.A(n_7452),
.B(n_7455),
.Y(n_8683)
);

OR2x2_ASAP7_75t_L g8684 ( 
.A(n_7542),
.B(n_6798),
.Y(n_8684)
);

HB1xp67_ASAP7_75t_L g8685 ( 
.A(n_7631),
.Y(n_8685)
);

OR2x2_ASAP7_75t_L g8686 ( 
.A(n_7564),
.B(n_6798),
.Y(n_8686)
);

INVx1_ASAP7_75t_L g8687 ( 
.A(n_7556),
.Y(n_8687)
);

AOI21x1_ASAP7_75t_L g8688 ( 
.A1(n_7782),
.A2(n_8172),
.B(n_7557),
.Y(n_8688)
);

INVx1_ASAP7_75t_L g8689 ( 
.A(n_7617),
.Y(n_8689)
);

AND2x2_ASAP7_75t_L g8690 ( 
.A(n_7452),
.B(n_6846),
.Y(n_8690)
);

INVx1_ASAP7_75t_L g8691 ( 
.A(n_7598),
.Y(n_8691)
);

AOI21xp5_ASAP7_75t_L g8692 ( 
.A1(n_7713),
.A2(n_6776),
.B(n_6752),
.Y(n_8692)
);

INVx2_ASAP7_75t_L g8693 ( 
.A(n_7954),
.Y(n_8693)
);

INVx1_ASAP7_75t_L g8694 ( 
.A(n_7677),
.Y(n_8694)
);

INVx1_ASAP7_75t_L g8695 ( 
.A(n_7677),
.Y(n_8695)
);

INVx3_ASAP7_75t_L g8696 ( 
.A(n_7487),
.Y(n_8696)
);

INVx1_ASAP7_75t_L g8697 ( 
.A(n_7787),
.Y(n_8697)
);

INVx2_ASAP7_75t_L g8698 ( 
.A(n_8329),
.Y(n_8698)
);

INVx2_ASAP7_75t_SL g8699 ( 
.A(n_7600),
.Y(n_8699)
);

INVx1_ASAP7_75t_L g8700 ( 
.A(n_7611),
.Y(n_8700)
);

HB1xp67_ASAP7_75t_L g8701 ( 
.A(n_7643),
.Y(n_8701)
);

INVx2_ASAP7_75t_L g8702 ( 
.A(n_8329),
.Y(n_8702)
);

INVx1_ASAP7_75t_L g8703 ( 
.A(n_7649),
.Y(n_8703)
);

AO21x2_ASAP7_75t_L g8704 ( 
.A1(n_7896),
.A2(n_7480),
.B(n_7470),
.Y(n_8704)
);

INVx2_ASAP7_75t_L g8705 ( 
.A(n_7567),
.Y(n_8705)
);

INVx2_ASAP7_75t_L g8706 ( 
.A(n_7567),
.Y(n_8706)
);

AND2x2_ASAP7_75t_L g8707 ( 
.A(n_7455),
.B(n_6846),
.Y(n_8707)
);

HB1xp67_ASAP7_75t_L g8708 ( 
.A(n_7665),
.Y(n_8708)
);

NAND2xp5_ASAP7_75t_L g8709 ( 
.A(n_7658),
.B(n_7184),
.Y(n_8709)
);

INVx1_ASAP7_75t_L g8710 ( 
.A(n_7615),
.Y(n_8710)
);

INVx1_ASAP7_75t_L g8711 ( 
.A(n_7615),
.Y(n_8711)
);

NAND2xp5_ASAP7_75t_L g8712 ( 
.A(n_7710),
.B(n_7188),
.Y(n_8712)
);

OR2x2_ASAP7_75t_L g8713 ( 
.A(n_7564),
.B(n_6833),
.Y(n_8713)
);

HB1xp67_ASAP7_75t_L g8714 ( 
.A(n_7666),
.Y(n_8714)
);

INVx1_ASAP7_75t_L g8715 ( 
.A(n_7617),
.Y(n_8715)
);

INVx2_ASAP7_75t_L g8716 ( 
.A(n_7594),
.Y(n_8716)
);

INVx4_ASAP7_75t_L g8717 ( 
.A(n_7607),
.Y(n_8717)
);

INVx2_ASAP7_75t_L g8718 ( 
.A(n_7594),
.Y(n_8718)
);

INVx2_ASAP7_75t_L g8719 ( 
.A(n_7601),
.Y(n_8719)
);

OR2x2_ASAP7_75t_L g8720 ( 
.A(n_7870),
.B(n_8099),
.Y(n_8720)
);

INVxp67_ASAP7_75t_L g8721 ( 
.A(n_8332),
.Y(n_8721)
);

AOI21x1_ASAP7_75t_L g8722 ( 
.A1(n_7782),
.A2(n_6977),
.B(n_7046),
.Y(n_8722)
);

NAND2xp33_ASAP7_75t_R g8723 ( 
.A(n_7711),
.B(n_5758),
.Y(n_8723)
);

HB1xp67_ASAP7_75t_L g8724 ( 
.A(n_7724),
.Y(n_8724)
);

INVx1_ASAP7_75t_L g8725 ( 
.A(n_7660),
.Y(n_8725)
);

AND2x2_ASAP7_75t_L g8726 ( 
.A(n_7597),
.B(n_7652),
.Y(n_8726)
);

INVx1_ASAP7_75t_L g8727 ( 
.A(n_7660),
.Y(n_8727)
);

INVx2_ASAP7_75t_L g8728 ( 
.A(n_7601),
.Y(n_8728)
);

BUFx2_ASAP7_75t_L g8729 ( 
.A(n_8063),
.Y(n_8729)
);

CKINVDCx5p33_ASAP7_75t_R g8730 ( 
.A(n_7938),
.Y(n_8730)
);

AND2x2_ASAP7_75t_L g8731 ( 
.A(n_7597),
.B(n_7652),
.Y(n_8731)
);

INVx3_ASAP7_75t_L g8732 ( 
.A(n_7487),
.Y(n_8732)
);

NAND2xp5_ASAP7_75t_L g8733 ( 
.A(n_7981),
.B(n_7188),
.Y(n_8733)
);

BUFx6f_ASAP7_75t_L g8734 ( 
.A(n_7607),
.Y(n_8734)
);

NAND2xp5_ASAP7_75t_L g8735 ( 
.A(n_7981),
.B(n_7002),
.Y(n_8735)
);

HB1xp67_ASAP7_75t_L g8736 ( 
.A(n_7730),
.Y(n_8736)
);

INVx1_ASAP7_75t_L g8737 ( 
.A(n_7649),
.Y(n_8737)
);

OR2x2_ASAP7_75t_L g8738 ( 
.A(n_7870),
.B(n_6833),
.Y(n_8738)
);

NAND2xp5_ASAP7_75t_L g8739 ( 
.A(n_7609),
.B(n_7026),
.Y(n_8739)
);

AND2x4_ASAP7_75t_L g8740 ( 
.A(n_8063),
.B(n_7195),
.Y(n_8740)
);

NAND2xp5_ASAP7_75t_L g8741 ( 
.A(n_7921),
.B(n_7060),
.Y(n_8741)
);

OR2x6_ASAP7_75t_L g8742 ( 
.A(n_7824),
.B(n_7057),
.Y(n_8742)
);

OA21x2_ASAP7_75t_L g8743 ( 
.A1(n_7718),
.A2(n_6472),
.B(n_6638),
.Y(n_8743)
);

OR2x2_ASAP7_75t_L g8744 ( 
.A(n_8099),
.B(n_7168),
.Y(n_8744)
);

INVx2_ASAP7_75t_L g8745 ( 
.A(n_7604),
.Y(n_8745)
);

AND2x2_ASAP7_75t_L g8746 ( 
.A(n_7672),
.B(n_6846),
.Y(n_8746)
);

OAI21x1_ASAP7_75t_L g8747 ( 
.A1(n_7538),
.A2(n_7557),
.B(n_7632),
.Y(n_8747)
);

INVx2_ASAP7_75t_L g8748 ( 
.A(n_7604),
.Y(n_8748)
);

INVx2_ASAP7_75t_L g8749 ( 
.A(n_7614),
.Y(n_8749)
);

INVx2_ASAP7_75t_L g8750 ( 
.A(n_7614),
.Y(n_8750)
);

INVx2_ASAP7_75t_L g8751 ( 
.A(n_7477),
.Y(n_8751)
);

HB1xp67_ASAP7_75t_L g8752 ( 
.A(n_7788),
.Y(n_8752)
);

OAI21xp5_ASAP7_75t_L g8753 ( 
.A1(n_7975),
.A2(n_7190),
.B(n_6676),
.Y(n_8753)
);

INVx2_ASAP7_75t_L g8754 ( 
.A(n_7477),
.Y(n_8754)
);

INVx1_ASAP7_75t_L g8755 ( 
.A(n_7745),
.Y(n_8755)
);

INVx2_ASAP7_75t_L g8756 ( 
.A(n_7516),
.Y(n_8756)
);

INVx5_ASAP7_75t_SL g8757 ( 
.A(n_8259),
.Y(n_8757)
);

BUFx3_ASAP7_75t_L g8758 ( 
.A(n_7765),
.Y(n_8758)
);

INVx2_ASAP7_75t_L g8759 ( 
.A(n_7516),
.Y(n_8759)
);

INVx3_ASAP7_75t_L g8760 ( 
.A(n_7634),
.Y(n_8760)
);

NOR2xp33_ASAP7_75t_L g8761 ( 
.A(n_7798),
.B(n_6198),
.Y(n_8761)
);

INVx1_ASAP7_75t_L g8762 ( 
.A(n_7746),
.Y(n_8762)
);

INVx1_ASAP7_75t_L g8763 ( 
.A(n_7746),
.Y(n_8763)
);

NOR2xp33_ASAP7_75t_L g8764 ( 
.A(n_7830),
.B(n_6198),
.Y(n_8764)
);

INVx2_ASAP7_75t_L g8765 ( 
.A(n_7527),
.Y(n_8765)
);

INVx1_ASAP7_75t_L g8766 ( 
.A(n_7767),
.Y(n_8766)
);

NAND2xp5_ASAP7_75t_L g8767 ( 
.A(n_7831),
.B(n_7592),
.Y(n_8767)
);

INVx1_ASAP7_75t_L g8768 ( 
.A(n_7667),
.Y(n_8768)
);

AO21x2_ASAP7_75t_L g8769 ( 
.A1(n_7896),
.A2(n_6839),
.B(n_6550),
.Y(n_8769)
);

INVx1_ASAP7_75t_L g8770 ( 
.A(n_7667),
.Y(n_8770)
);

INVx2_ASAP7_75t_SL g8771 ( 
.A(n_7607),
.Y(n_8771)
);

AOI21x1_ASAP7_75t_L g8772 ( 
.A1(n_8172),
.A2(n_6940),
.B(n_6935),
.Y(n_8772)
);

INVx2_ASAP7_75t_L g8773 ( 
.A(n_7527),
.Y(n_8773)
);

HB1xp67_ASAP7_75t_SL g8774 ( 
.A(n_7929),
.Y(n_8774)
);

INVx1_ASAP7_75t_L g8775 ( 
.A(n_7683),
.Y(n_8775)
);

INVx1_ASAP7_75t_L g8776 ( 
.A(n_7683),
.Y(n_8776)
);

AND2x2_ASAP7_75t_L g8777 ( 
.A(n_7672),
.B(n_6846),
.Y(n_8777)
);

INVx3_ASAP7_75t_L g8778 ( 
.A(n_7487),
.Y(n_8778)
);

INVx2_ASAP7_75t_L g8779 ( 
.A(n_7531),
.Y(n_8779)
);

INVx1_ASAP7_75t_L g8780 ( 
.A(n_7744),
.Y(n_8780)
);

OAI21x1_ASAP7_75t_L g8781 ( 
.A1(n_7632),
.A2(n_6838),
.B(n_7190),
.Y(n_8781)
);

INVx1_ASAP7_75t_L g8782 ( 
.A(n_7639),
.Y(n_8782)
);

BUFx2_ASAP7_75t_L g8783 ( 
.A(n_8063),
.Y(n_8783)
);

INVx1_ASAP7_75t_L g8784 ( 
.A(n_7639),
.Y(n_8784)
);

HB1xp67_ASAP7_75t_L g8785 ( 
.A(n_7791),
.Y(n_8785)
);

INVx1_ASAP7_75t_L g8786 ( 
.A(n_7767),
.Y(n_8786)
);

INVx1_ASAP7_75t_L g8787 ( 
.A(n_7776),
.Y(n_8787)
);

INVx1_ASAP7_75t_L g8788 ( 
.A(n_7776),
.Y(n_8788)
);

INVx1_ASAP7_75t_L g8789 ( 
.A(n_7809),
.Y(n_8789)
);

INVx1_ASAP7_75t_L g8790 ( 
.A(n_7809),
.Y(n_8790)
);

HB1xp67_ASAP7_75t_L g8791 ( 
.A(n_7813),
.Y(n_8791)
);

AOI21xp5_ASAP7_75t_L g8792 ( 
.A1(n_7490),
.A2(n_6776),
.B(n_6752),
.Y(n_8792)
);

HB1xp67_ASAP7_75t_L g8793 ( 
.A(n_7872),
.Y(n_8793)
);

AOI21x1_ASAP7_75t_L g8794 ( 
.A1(n_7805),
.A2(n_6940),
.B(n_6935),
.Y(n_8794)
);

NAND2x1p5_ASAP7_75t_L g8795 ( 
.A(n_7874),
.B(n_7291),
.Y(n_8795)
);

AND2x6_ASAP7_75t_SL g8796 ( 
.A(n_8057),
.B(n_5899),
.Y(n_8796)
);

INVx2_ASAP7_75t_L g8797 ( 
.A(n_7531),
.Y(n_8797)
);

INVx3_ASAP7_75t_L g8798 ( 
.A(n_7487),
.Y(n_8798)
);

INVx1_ASAP7_75t_L g8799 ( 
.A(n_7737),
.Y(n_8799)
);

AND2x2_ASAP7_75t_L g8800 ( 
.A(n_7712),
.B(n_6846),
.Y(n_8800)
);

AO21x2_ASAP7_75t_L g8801 ( 
.A1(n_7470),
.A2(n_6550),
.B(n_6559),
.Y(n_8801)
);

INVx1_ASAP7_75t_SL g8802 ( 
.A(n_7969),
.Y(n_8802)
);

INVx1_ASAP7_75t_L g8803 ( 
.A(n_7737),
.Y(n_8803)
);

INVx1_ASAP7_75t_L g8804 ( 
.A(n_7794),
.Y(n_8804)
);

INVx2_ASAP7_75t_L g8805 ( 
.A(n_7537),
.Y(n_8805)
);

INVx2_ASAP7_75t_L g8806 ( 
.A(n_7537),
.Y(n_8806)
);

INVx2_ASAP7_75t_L g8807 ( 
.A(n_7546),
.Y(n_8807)
);

INVxp33_ASAP7_75t_L g8808 ( 
.A(n_7505),
.Y(n_8808)
);

OA21x2_ASAP7_75t_L g8809 ( 
.A1(n_7718),
.A2(n_6638),
.B(n_6501),
.Y(n_8809)
);

INVx2_ASAP7_75t_L g8810 ( 
.A(n_7546),
.Y(n_8810)
);

INVx1_ASAP7_75t_L g8811 ( 
.A(n_7580),
.Y(n_8811)
);

INVx3_ASAP7_75t_L g8812 ( 
.A(n_7634),
.Y(n_8812)
);

AND2x2_ASAP7_75t_L g8813 ( 
.A(n_7712),
.B(n_6933),
.Y(n_8813)
);

INVx1_ASAP7_75t_L g8814 ( 
.A(n_7811),
.Y(n_8814)
);

BUFx3_ASAP7_75t_L g8815 ( 
.A(n_8045),
.Y(n_8815)
);

INVx1_ASAP7_75t_L g8816 ( 
.A(n_7811),
.Y(n_8816)
);

BUFx2_ASAP7_75t_L g8817 ( 
.A(n_7774),
.Y(n_8817)
);

INVx2_ASAP7_75t_L g8818 ( 
.A(n_7548),
.Y(n_8818)
);

INVx2_ASAP7_75t_L g8819 ( 
.A(n_7548),
.Y(n_8819)
);

INVx2_ASAP7_75t_L g8820 ( 
.A(n_7555),
.Y(n_8820)
);

INVx2_ASAP7_75t_SL g8821 ( 
.A(n_7702),
.Y(n_8821)
);

INVx2_ASAP7_75t_L g8822 ( 
.A(n_7555),
.Y(n_8822)
);

INVx1_ASAP7_75t_L g8823 ( 
.A(n_7722),
.Y(n_8823)
);

OAI21x1_ASAP7_75t_L g8824 ( 
.A1(n_7805),
.A2(n_6838),
.B(n_7275),
.Y(n_8824)
);

INVx2_ASAP7_75t_L g8825 ( 
.A(n_7558),
.Y(n_8825)
);

INVx2_ASAP7_75t_L g8826 ( 
.A(n_7558),
.Y(n_8826)
);

INVx2_ASAP7_75t_L g8827 ( 
.A(n_7562),
.Y(n_8827)
);

INVx2_ASAP7_75t_L g8828 ( 
.A(n_7562),
.Y(n_8828)
);

INVx2_ASAP7_75t_L g8829 ( 
.A(n_7622),
.Y(n_8829)
);

INVx8_ASAP7_75t_L g8830 ( 
.A(n_7647),
.Y(n_8830)
);

OAI21x1_ASAP7_75t_L g8831 ( 
.A1(n_8334),
.A2(n_7275),
.B(n_6946),
.Y(n_8831)
);

INVx2_ASAP7_75t_L g8832 ( 
.A(n_7622),
.Y(n_8832)
);

AOI21x1_ASAP7_75t_L g8833 ( 
.A1(n_7431),
.A2(n_6946),
.B(n_6912),
.Y(n_8833)
);

INVx3_ASAP7_75t_L g8834 ( 
.A(n_7634),
.Y(n_8834)
);

INVx3_ASAP7_75t_L g8835 ( 
.A(n_7634),
.Y(n_8835)
);

AND2x4_ASAP7_75t_L g8836 ( 
.A(n_7874),
.B(n_7195),
.Y(n_8836)
);

BUFx6f_ASAP7_75t_L g8837 ( 
.A(n_7702),
.Y(n_8837)
);

INVx1_ASAP7_75t_L g8838 ( 
.A(n_7745),
.Y(n_8838)
);

INVx2_ASAP7_75t_L g8839 ( 
.A(n_7624),
.Y(n_8839)
);

INVx2_ASAP7_75t_SL g8840 ( 
.A(n_7702),
.Y(n_8840)
);

INVx1_ASAP7_75t_L g8841 ( 
.A(n_7705),
.Y(n_8841)
);

INVx1_ASAP7_75t_L g8842 ( 
.A(n_7705),
.Y(n_8842)
);

INVx1_ASAP7_75t_L g8843 ( 
.A(n_7779),
.Y(n_8843)
);

AND2x2_ASAP7_75t_L g8844 ( 
.A(n_7732),
.B(n_6933),
.Y(n_8844)
);

INVx2_ASAP7_75t_SL g8845 ( 
.A(n_7800),
.Y(n_8845)
);

NAND2xp5_ASAP7_75t_L g8846 ( 
.A(n_7831),
.B(n_7060),
.Y(n_8846)
);

INVx1_ASAP7_75t_L g8847 ( 
.A(n_7779),
.Y(n_8847)
);

BUFx8_ASAP7_75t_SL g8848 ( 
.A(n_7769),
.Y(n_8848)
);

OAI21x1_ASAP7_75t_L g8849 ( 
.A1(n_8334),
.A2(n_6525),
.B(n_6523),
.Y(n_8849)
);

OA21x2_ASAP7_75t_L g8850 ( 
.A1(n_7719),
.A2(n_6638),
.B(n_6501),
.Y(n_8850)
);

AO21x2_ASAP7_75t_L g8851 ( 
.A1(n_7470),
.A2(n_6550),
.B(n_6559),
.Y(n_8851)
);

BUFx2_ASAP7_75t_L g8852 ( 
.A(n_7774),
.Y(n_8852)
);

INVx2_ASAP7_75t_L g8853 ( 
.A(n_7624),
.Y(n_8853)
);

INVx1_ASAP7_75t_L g8854 ( 
.A(n_7722),
.Y(n_8854)
);

INVx2_ASAP7_75t_L g8855 ( 
.A(n_7638),
.Y(n_8855)
);

INVx2_ASAP7_75t_SL g8856 ( 
.A(n_7774),
.Y(n_8856)
);

INVx1_ASAP7_75t_L g8857 ( 
.A(n_7775),
.Y(n_8857)
);

AOI21x1_ASAP7_75t_L g8858 ( 
.A1(n_7431),
.A2(n_6452),
.B(n_6447),
.Y(n_8858)
);

OAI22xp33_ASAP7_75t_L g8859 ( 
.A1(n_7918),
.A2(n_7025),
.B1(n_6709),
.B2(n_6693),
.Y(n_8859)
);

OAI22xp5_ASAP7_75t_L g8860 ( 
.A1(n_7464),
.A2(n_6745),
.B1(n_6859),
.B2(n_7390),
.Y(n_8860)
);

INVx1_ASAP7_75t_L g8861 ( 
.A(n_7744),
.Y(n_8861)
);

OR2x2_ASAP7_75t_L g8862 ( 
.A(n_7581),
.B(n_7168),
.Y(n_8862)
);

NAND2xp5_ASAP7_75t_L g8863 ( 
.A(n_8114),
.B(n_8120),
.Y(n_8863)
);

INVx1_ASAP7_75t_L g8864 ( 
.A(n_7780),
.Y(n_8864)
);

BUFx2_ASAP7_75t_L g8865 ( 
.A(n_7711),
.Y(n_8865)
);

INVx1_ASAP7_75t_L g8866 ( 
.A(n_7794),
.Y(n_8866)
);

INVx2_ASAP7_75t_L g8867 ( 
.A(n_7638),
.Y(n_8867)
);

INVx1_ASAP7_75t_L g8868 ( 
.A(n_7796),
.Y(n_8868)
);

INVx2_ASAP7_75t_L g8869 ( 
.A(n_7654),
.Y(n_8869)
);

INVx1_ASAP7_75t_L g8870 ( 
.A(n_7796),
.Y(n_8870)
);

BUFx2_ASAP7_75t_L g8871 ( 
.A(n_7781),
.Y(n_8871)
);

INVx1_ASAP7_75t_L g8872 ( 
.A(n_7812),
.Y(n_8872)
);

INVx2_ASAP7_75t_L g8873 ( 
.A(n_7654),
.Y(n_8873)
);

OAI21x1_ASAP7_75t_L g8874 ( 
.A1(n_8344),
.A2(n_6525),
.B(n_6523),
.Y(n_8874)
);

INVx1_ASAP7_75t_L g8875 ( 
.A(n_7760),
.Y(n_8875)
);

INVx2_ASAP7_75t_L g8876 ( 
.A(n_7656),
.Y(n_8876)
);

NAND2x1p5_ASAP7_75t_L g8877 ( 
.A(n_7874),
.B(n_7291),
.Y(n_8877)
);

INVx2_ASAP7_75t_L g8878 ( 
.A(n_7656),
.Y(n_8878)
);

BUFx4f_ASAP7_75t_SL g8879 ( 
.A(n_7437),
.Y(n_8879)
);

INVx2_ASAP7_75t_L g8880 ( 
.A(n_7664),
.Y(n_8880)
);

BUFx12f_ASAP7_75t_L g8881 ( 
.A(n_8025),
.Y(n_8881)
);

INVx1_ASAP7_75t_L g8882 ( 
.A(n_7775),
.Y(n_8882)
);

INVx1_ASAP7_75t_L g8883 ( 
.A(n_7832),
.Y(n_8883)
);

INVx1_ASAP7_75t_L g8884 ( 
.A(n_7832),
.Y(n_8884)
);

INVx2_ASAP7_75t_L g8885 ( 
.A(n_7664),
.Y(n_8885)
);

INVx2_ASAP7_75t_L g8886 ( 
.A(n_7679),
.Y(n_8886)
);

OAI22xp5_ASAP7_75t_L g8887 ( 
.A1(n_7411),
.A2(n_6758),
.B1(n_7288),
.B2(n_7272),
.Y(n_8887)
);

INVx1_ASAP7_75t_L g8888 ( 
.A(n_7764),
.Y(n_8888)
);

AOI21x1_ASAP7_75t_L g8889 ( 
.A1(n_7436),
.A2(n_6452),
.B(n_6447),
.Y(n_8889)
);

INVx2_ASAP7_75t_SL g8890 ( 
.A(n_8123),
.Y(n_8890)
);

INVx1_ASAP7_75t_L g8891 ( 
.A(n_7764),
.Y(n_8891)
);

INVx1_ASAP7_75t_L g8892 ( 
.A(n_7823),
.Y(n_8892)
);

INVx1_ASAP7_75t_L g8893 ( 
.A(n_7823),
.Y(n_8893)
);

INVx3_ASAP7_75t_L g8894 ( 
.A(n_7532),
.Y(n_8894)
);

AND2x4_ASAP7_75t_L g8895 ( 
.A(n_7874),
.B(n_7195),
.Y(n_8895)
);

INVx1_ASAP7_75t_L g8896 ( 
.A(n_7826),
.Y(n_8896)
);

INVx2_ASAP7_75t_L g8897 ( 
.A(n_7679),
.Y(n_8897)
);

INVx2_ASAP7_75t_L g8898 ( 
.A(n_7690),
.Y(n_8898)
);

AO21x2_ASAP7_75t_L g8899 ( 
.A1(n_7480),
.A2(n_6550),
.B(n_6559),
.Y(n_8899)
);

HB1xp67_ASAP7_75t_L g8900 ( 
.A(n_7892),
.Y(n_8900)
);

INVx3_ASAP7_75t_L g8901 ( 
.A(n_7532),
.Y(n_8901)
);

AND2x2_ASAP7_75t_L g8902 ( 
.A(n_7732),
.B(n_6933),
.Y(n_8902)
);

BUFx2_ASAP7_75t_L g8903 ( 
.A(n_7781),
.Y(n_8903)
);

OAI21x1_ASAP7_75t_L g8904 ( 
.A1(n_8344),
.A2(n_6525),
.B(n_6523),
.Y(n_8904)
);

INVx1_ASAP7_75t_L g8905 ( 
.A(n_7849),
.Y(n_8905)
);

AND2x2_ASAP7_75t_L g8906 ( 
.A(n_7772),
.B(n_6933),
.Y(n_8906)
);

INVx1_ASAP7_75t_L g8907 ( 
.A(n_7849),
.Y(n_8907)
);

A2O1A1Ixp33_ASAP7_75t_L g8908 ( 
.A1(n_7900),
.A2(n_8098),
.B(n_7918),
.C(n_7569),
.Y(n_8908)
);

INVx2_ASAP7_75t_L g8909 ( 
.A(n_7690),
.Y(n_8909)
);

AOI22xp5_ASAP7_75t_L g8910 ( 
.A1(n_7511),
.A2(n_7303),
.B1(n_7249),
.B2(n_6840),
.Y(n_8910)
);

AND2x4_ASAP7_75t_L g8911 ( 
.A(n_7874),
.B(n_7195),
.Y(n_8911)
);

INVx3_ASAP7_75t_L g8912 ( 
.A(n_7532),
.Y(n_8912)
);

INVx2_ASAP7_75t_L g8913 ( 
.A(n_7691),
.Y(n_8913)
);

AND2x2_ASAP7_75t_L g8914 ( 
.A(n_7772),
.B(n_6933),
.Y(n_8914)
);

INVx2_ASAP7_75t_L g8915 ( 
.A(n_7691),
.Y(n_8915)
);

INVx1_ASAP7_75t_SL g8916 ( 
.A(n_8014),
.Y(n_8916)
);

INVx2_ASAP7_75t_L g8917 ( 
.A(n_7692),
.Y(n_8917)
);

OAI21x1_ASAP7_75t_L g8918 ( 
.A1(n_7532),
.A2(n_7568),
.B(n_7549),
.Y(n_8918)
);

HB1xp67_ASAP7_75t_L g8919 ( 
.A(n_7907),
.Y(n_8919)
);

INVx2_ASAP7_75t_L g8920 ( 
.A(n_7692),
.Y(n_8920)
);

BUFx3_ASAP7_75t_L g8921 ( 
.A(n_7668),
.Y(n_8921)
);

INVx1_ASAP7_75t_L g8922 ( 
.A(n_7816),
.Y(n_8922)
);

BUFx2_ASAP7_75t_L g8923 ( 
.A(n_8111),
.Y(n_8923)
);

INVx2_ASAP7_75t_L g8924 ( 
.A(n_7695),
.Y(n_8924)
);

INVx2_ASAP7_75t_L g8925 ( 
.A(n_7695),
.Y(n_8925)
);

BUFx3_ASAP7_75t_L g8926 ( 
.A(n_7668),
.Y(n_8926)
);

INVx2_ASAP7_75t_L g8927 ( 
.A(n_7701),
.Y(n_8927)
);

AOI22xp33_ASAP7_75t_L g8928 ( 
.A1(n_7663),
.A2(n_6443),
.B1(n_7249),
.B2(n_6653),
.Y(n_8928)
);

INVx2_ASAP7_75t_L g8929 ( 
.A(n_7701),
.Y(n_8929)
);

NAND2x1p5_ASAP7_75t_L g8930 ( 
.A(n_8178),
.B(n_7291),
.Y(n_8930)
);

AND2x2_ASAP7_75t_SL g8931 ( 
.A(n_8323),
.B(n_7208),
.Y(n_8931)
);

INVx1_ASAP7_75t_L g8932 ( 
.A(n_7888),
.Y(n_8932)
);

INVx3_ASAP7_75t_L g8933 ( 
.A(n_7549),
.Y(n_8933)
);

INVx2_ASAP7_75t_L g8934 ( 
.A(n_7706),
.Y(n_8934)
);

BUFx2_ASAP7_75t_L g8935 ( 
.A(n_8111),
.Y(n_8935)
);

AND2x2_ASAP7_75t_L g8936 ( 
.A(n_7871),
.B(n_7928),
.Y(n_8936)
);

INVx1_ASAP7_75t_L g8937 ( 
.A(n_7888),
.Y(n_8937)
);

INVx2_ASAP7_75t_L g8938 ( 
.A(n_7706),
.Y(n_8938)
);

INVx1_ASAP7_75t_L g8939 ( 
.A(n_7760),
.Y(n_8939)
);

INVx2_ASAP7_75t_L g8940 ( 
.A(n_7707),
.Y(n_8940)
);

INVx2_ASAP7_75t_L g8941 ( 
.A(n_7707),
.Y(n_8941)
);

INVx1_ASAP7_75t_L g8942 ( 
.A(n_7734),
.Y(n_8942)
);

OAI21x1_ASAP7_75t_L g8943 ( 
.A1(n_7549),
.A2(n_6594),
.B(n_6588),
.Y(n_8943)
);

INVx2_ASAP7_75t_SL g8944 ( 
.A(n_8123),
.Y(n_8944)
);

OAI22xp33_ASAP7_75t_L g8945 ( 
.A1(n_7958),
.A2(n_7025),
.B1(n_6709),
.B2(n_6693),
.Y(n_8945)
);

INVx1_ASAP7_75t_L g8946 ( 
.A(n_7734),
.Y(n_8946)
);

INVx3_ASAP7_75t_L g8947 ( 
.A(n_7549),
.Y(n_8947)
);

HB1xp67_ASAP7_75t_L g8948 ( 
.A(n_7990),
.Y(n_8948)
);

OAI21x1_ASAP7_75t_L g8949 ( 
.A1(n_7568),
.A2(n_6594),
.B(n_6588),
.Y(n_8949)
);

INVx1_ASAP7_75t_L g8950 ( 
.A(n_7816),
.Y(n_8950)
);

INVx2_ASAP7_75t_L g8951 ( 
.A(n_7708),
.Y(n_8951)
);

INVx1_ASAP7_75t_L g8952 ( 
.A(n_7972),
.Y(n_8952)
);

INVx2_ASAP7_75t_L g8953 ( 
.A(n_7708),
.Y(n_8953)
);

INVx1_ASAP7_75t_L g8954 ( 
.A(n_7859),
.Y(n_8954)
);

OAI22xp33_ASAP7_75t_L g8955 ( 
.A1(n_7958),
.A2(n_6709),
.B1(n_6693),
.B2(n_6843),
.Y(n_8955)
);

OAI21x1_ASAP7_75t_L g8956 ( 
.A1(n_7568),
.A2(n_6594),
.B(n_6588),
.Y(n_8956)
);

INVx3_ASAP7_75t_L g8957 ( 
.A(n_7568),
.Y(n_8957)
);

INVx2_ASAP7_75t_SL g8958 ( 
.A(n_8123),
.Y(n_8958)
);

INVx1_ASAP7_75t_L g8959 ( 
.A(n_7804),
.Y(n_8959)
);

INVx1_ASAP7_75t_L g8960 ( 
.A(n_7804),
.Y(n_8960)
);

INVx1_ASAP7_75t_L g8961 ( 
.A(n_7880),
.Y(n_8961)
);

INVx2_ASAP7_75t_L g8962 ( 
.A(n_7448),
.Y(n_8962)
);

INVx3_ASAP7_75t_L g8963 ( 
.A(n_7584),
.Y(n_8963)
);

INVx1_ASAP7_75t_L g8964 ( 
.A(n_7880),
.Y(n_8964)
);

INVx3_ASAP7_75t_L g8965 ( 
.A(n_7584),
.Y(n_8965)
);

INVx1_ASAP7_75t_L g8966 ( 
.A(n_7881),
.Y(n_8966)
);

INVx1_ASAP7_75t_L g8967 ( 
.A(n_7881),
.Y(n_8967)
);

OAI21x1_ASAP7_75t_L g8968 ( 
.A1(n_7584),
.A2(n_6700),
.B(n_6792),
.Y(n_8968)
);

AND2x2_ASAP7_75t_L g8969 ( 
.A(n_7871),
.B(n_6508),
.Y(n_8969)
);

INVx1_ASAP7_75t_SL g8970 ( 
.A(n_7579),
.Y(n_8970)
);

INVx1_ASAP7_75t_L g8971 ( 
.A(n_7822),
.Y(n_8971)
);

NAND2xp5_ASAP7_75t_L g8972 ( 
.A(n_8124),
.B(n_7393),
.Y(n_8972)
);

INVx2_ASAP7_75t_SL g8973 ( 
.A(n_8123),
.Y(n_8973)
);

INVx2_ASAP7_75t_L g8974 ( 
.A(n_7448),
.Y(n_8974)
);

INVx2_ASAP7_75t_SL g8975 ( 
.A(n_8143),
.Y(n_8975)
);

NAND2xp5_ASAP7_75t_L g8976 ( 
.A(n_7841),
.B(n_7393),
.Y(n_8976)
);

INVx1_ASAP7_75t_L g8977 ( 
.A(n_7889),
.Y(n_8977)
);

INVx2_ASAP7_75t_L g8978 ( 
.A(n_7454),
.Y(n_8978)
);

HB1xp67_ASAP7_75t_L g8979 ( 
.A(n_7997),
.Y(n_8979)
);

AO21x1_ASAP7_75t_SL g8980 ( 
.A1(n_8098),
.A2(n_6938),
.B(n_6870),
.Y(n_8980)
);

AOI21x1_ASAP7_75t_L g8981 ( 
.A1(n_7436),
.A2(n_6981),
.B(n_6875),
.Y(n_8981)
);

INVx2_ASAP7_75t_L g8982 ( 
.A(n_7454),
.Y(n_8982)
);

INVx1_ASAP7_75t_L g8983 ( 
.A(n_7780),
.Y(n_8983)
);

INVx1_ASAP7_75t_L g8984 ( 
.A(n_7659),
.Y(n_8984)
);

AOI22xp33_ASAP7_75t_L g8985 ( 
.A1(n_7703),
.A2(n_7420),
.B1(n_8046),
.B2(n_7790),
.Y(n_8985)
);

NAND2xp5_ASAP7_75t_L g8986 ( 
.A(n_7843),
.B(n_7326),
.Y(n_8986)
);

INVx2_ASAP7_75t_SL g8987 ( 
.A(n_8143),
.Y(n_8987)
);

BUFx3_ASAP7_75t_L g8988 ( 
.A(n_7668),
.Y(n_8988)
);

AND2x2_ASAP7_75t_L g8989 ( 
.A(n_7928),
.B(n_6508),
.Y(n_8989)
);

AND2x2_ASAP7_75t_L g8990 ( 
.A(n_8049),
.B(n_6508),
.Y(n_8990)
);

INVx1_ASAP7_75t_L g8991 ( 
.A(n_7659),
.Y(n_8991)
);

NOR2xp33_ASAP7_75t_L g8992 ( 
.A(n_7802),
.B(n_6274),
.Y(n_8992)
);

INVx1_ASAP7_75t_L g8993 ( 
.A(n_7675),
.Y(n_8993)
);

OR2x2_ASAP7_75t_L g8994 ( 
.A(n_7581),
.B(n_6938),
.Y(n_8994)
);

INVx2_ASAP7_75t_L g8995 ( 
.A(n_7460),
.Y(n_8995)
);

BUFx6f_ASAP7_75t_L g8996 ( 
.A(n_7682),
.Y(n_8996)
);

HB1xp67_ASAP7_75t_L g8997 ( 
.A(n_8004),
.Y(n_8997)
);

INVx1_ASAP7_75t_L g8998 ( 
.A(n_7812),
.Y(n_8998)
);

INVx2_ASAP7_75t_L g8999 ( 
.A(n_7460),
.Y(n_8999)
);

INVx1_ASAP7_75t_L g9000 ( 
.A(n_7675),
.Y(n_9000)
);

INVx2_ASAP7_75t_L g9001 ( 
.A(n_7461),
.Y(n_9001)
);

OR2x6_ASAP7_75t_L g9002 ( 
.A(n_8333),
.B(n_7291),
.Y(n_9002)
);

HB1xp67_ASAP7_75t_L g9003 ( 
.A(n_8010),
.Y(n_9003)
);

INVx1_ASAP7_75t_L g9004 ( 
.A(n_7763),
.Y(n_9004)
);

INVx2_ASAP7_75t_L g9005 ( 
.A(n_7461),
.Y(n_9005)
);

INVx3_ASAP7_75t_L g9006 ( 
.A(n_7584),
.Y(n_9006)
);

OAI21x1_ASAP7_75t_L g9007 ( 
.A1(n_7623),
.A2(n_6700),
.B(n_6792),
.Y(n_9007)
);

INVx3_ASAP7_75t_L g9008 ( 
.A(n_7623),
.Y(n_9008)
);

OAI21x1_ASAP7_75t_L g9009 ( 
.A1(n_7623),
.A2(n_6700),
.B(n_6792),
.Y(n_9009)
);

CKINVDCx6p67_ASAP7_75t_R g9010 ( 
.A(n_7682),
.Y(n_9010)
);

INVx3_ASAP7_75t_L g9011 ( 
.A(n_7623),
.Y(n_9011)
);

AO21x2_ASAP7_75t_L g9012 ( 
.A1(n_7480),
.A2(n_6559),
.B(n_6822),
.Y(n_9012)
);

AND2x2_ASAP7_75t_L g9013 ( 
.A(n_8049),
.B(n_6546),
.Y(n_9013)
);

INVx1_ASAP7_75t_L g9014 ( 
.A(n_7859),
.Y(n_9014)
);

AND2x2_ASAP7_75t_L g9015 ( 
.A(n_8311),
.B(n_7491),
.Y(n_9015)
);

AO31x2_ASAP7_75t_L g9016 ( 
.A1(n_7481),
.A2(n_7291),
.A3(n_6703),
.B(n_6471),
.Y(n_9016)
);

INVx1_ASAP7_75t_L g9017 ( 
.A(n_7971),
.Y(n_9017)
);

INVx2_ASAP7_75t_SL g9018 ( 
.A(n_8143),
.Y(n_9018)
);

INVx2_ASAP7_75t_L g9019 ( 
.A(n_7476),
.Y(n_9019)
);

OAI21xp5_ASAP7_75t_SL g9020 ( 
.A1(n_7886),
.A2(n_6607),
.B(n_6882),
.Y(n_9020)
);

AOI21x1_ASAP7_75t_L g9021 ( 
.A1(n_7466),
.A2(n_6981),
.B(n_6875),
.Y(n_9021)
);

AOI21x1_ASAP7_75t_L g9022 ( 
.A1(n_7466),
.A2(n_7336),
.B(n_7016),
.Y(n_9022)
);

AND2x2_ASAP7_75t_L g9023 ( 
.A(n_8311),
.B(n_6546),
.Y(n_9023)
);

INVx2_ASAP7_75t_L g9024 ( 
.A(n_7476),
.Y(n_9024)
);

AND2x2_ASAP7_75t_L g9025 ( 
.A(n_7491),
.B(n_6546),
.Y(n_9025)
);

INVx2_ASAP7_75t_L g9026 ( 
.A(n_8174),
.Y(n_9026)
);

AND2x2_ASAP7_75t_L g9027 ( 
.A(n_7851),
.B(n_6569),
.Y(n_9027)
);

AOI21xp5_ASAP7_75t_L g9028 ( 
.A1(n_7827),
.A2(n_7125),
.B(n_7082),
.Y(n_9028)
);

AO31x2_ASAP7_75t_L g9029 ( 
.A1(n_7481),
.A2(n_6703),
.A3(n_6471),
.B(n_6479),
.Y(n_9029)
);

INVx1_ASAP7_75t_L g9030 ( 
.A(n_7889),
.Y(n_9030)
);

INVx1_ASAP7_75t_L g9031 ( 
.A(n_7911),
.Y(n_9031)
);

INVx1_ASAP7_75t_L g9032 ( 
.A(n_7911),
.Y(n_9032)
);

INVx1_ASAP7_75t_L g9033 ( 
.A(n_7923),
.Y(n_9033)
);

INVx2_ASAP7_75t_L g9034 ( 
.A(n_8174),
.Y(n_9034)
);

HB1xp67_ASAP7_75t_L g9035 ( 
.A(n_8030),
.Y(n_9035)
);

INVx1_ASAP7_75t_L g9036 ( 
.A(n_7923),
.Y(n_9036)
);

OAI21xp5_ASAP7_75t_L g9037 ( 
.A1(n_8078),
.A2(n_6676),
.B(n_7082),
.Y(n_9037)
);

OAI21x1_ASAP7_75t_L g9038 ( 
.A1(n_7844),
.A2(n_6501),
.B(n_6607),
.Y(n_9038)
);

NAND2x1_ASAP7_75t_L g9039 ( 
.A(n_7485),
.B(n_6573),
.Y(n_9039)
);

OR2x2_ASAP7_75t_L g9040 ( 
.A(n_7752),
.B(n_6938),
.Y(n_9040)
);

INVx2_ASAP7_75t_L g9041 ( 
.A(n_8174),
.Y(n_9041)
);

AND2x2_ASAP7_75t_L g9042 ( 
.A(n_7851),
.B(n_6569),
.Y(n_9042)
);

NAND2xp5_ASAP7_75t_L g9043 ( 
.A(n_7726),
.B(n_7326),
.Y(n_9043)
);

INVx2_ASAP7_75t_L g9044 ( 
.A(n_7977),
.Y(n_9044)
);

INVx1_ASAP7_75t_L g9045 ( 
.A(n_7837),
.Y(n_9045)
);

NAND2x1_ASAP7_75t_L g9046 ( 
.A(n_7736),
.B(n_6684),
.Y(n_9046)
);

INVx1_ASAP7_75t_L g9047 ( 
.A(n_7837),
.Y(n_9047)
);

AOI22xp33_ASAP7_75t_L g9048 ( 
.A1(n_7778),
.A2(n_6443),
.B1(n_6653),
.B2(n_6644),
.Y(n_9048)
);

BUFx2_ASAP7_75t_L g9049 ( 
.A(n_8054),
.Y(n_9049)
);

AND2x4_ASAP7_75t_L g9050 ( 
.A(n_8266),
.B(n_7195),
.Y(n_9050)
);

AOI21xp5_ASAP7_75t_L g9051 ( 
.A1(n_8110),
.A2(n_7810),
.B(n_8162),
.Y(n_9051)
);

INVx3_ASAP7_75t_L g9052 ( 
.A(n_8116),
.Y(n_9052)
);

INVx1_ASAP7_75t_L g9053 ( 
.A(n_7862),
.Y(n_9053)
);

HB1xp67_ASAP7_75t_L g9054 ( 
.A(n_8076),
.Y(n_9054)
);

AO21x2_ASAP7_75t_L g9055 ( 
.A1(n_7481),
.A2(n_6822),
.B(n_6537),
.Y(n_9055)
);

INVx1_ASAP7_75t_L g9056 ( 
.A(n_7763),
.Y(n_9056)
);

INVx2_ASAP7_75t_L g9057 ( 
.A(n_7977),
.Y(n_9057)
);

INVx1_ASAP7_75t_L g9058 ( 
.A(n_7971),
.Y(n_9058)
);

OR2x6_ASAP7_75t_L g9059 ( 
.A(n_8333),
.B(n_6418),
.Y(n_9059)
);

INVx2_ASAP7_75t_SL g9060 ( 
.A(n_8143),
.Y(n_9060)
);

NOR2xp33_ASAP7_75t_L g9061 ( 
.A(n_7771),
.B(n_6274),
.Y(n_9061)
);

INVx1_ASAP7_75t_L g9062 ( 
.A(n_7951),
.Y(n_9062)
);

INVx1_ASAP7_75t_L g9063 ( 
.A(n_7951),
.Y(n_9063)
);

INVx2_ASAP7_75t_L g9064 ( 
.A(n_7983),
.Y(n_9064)
);

AND2x4_ASAP7_75t_L g9065 ( 
.A(n_8266),
.B(n_7195),
.Y(n_9065)
);

INVx1_ASAP7_75t_L g9066 ( 
.A(n_8036),
.Y(n_9066)
);

INVx1_ASAP7_75t_L g9067 ( 
.A(n_8036),
.Y(n_9067)
);

HB1xp67_ASAP7_75t_L g9068 ( 
.A(n_8107),
.Y(n_9068)
);

INVx1_ASAP7_75t_L g9069 ( 
.A(n_8048),
.Y(n_9069)
);

INVx1_ASAP7_75t_L g9070 ( 
.A(n_8048),
.Y(n_9070)
);

INVx3_ASAP7_75t_L g9071 ( 
.A(n_8116),
.Y(n_9071)
);

AND2x2_ASAP7_75t_L g9072 ( 
.A(n_7984),
.B(n_6569),
.Y(n_9072)
);

INVx1_ASAP7_75t_L g9073 ( 
.A(n_8082),
.Y(n_9073)
);

INVx1_ASAP7_75t_L g9074 ( 
.A(n_8082),
.Y(n_9074)
);

INVx1_ASAP7_75t_L g9075 ( 
.A(n_8103),
.Y(n_9075)
);

INVx1_ASAP7_75t_L g9076 ( 
.A(n_8103),
.Y(n_9076)
);

AO21x2_ASAP7_75t_L g9077 ( 
.A1(n_7483),
.A2(n_6822),
.B(n_6537),
.Y(n_9077)
);

INVx2_ASAP7_75t_L g9078 ( 
.A(n_7983),
.Y(n_9078)
);

HB1xp67_ASAP7_75t_L g9079 ( 
.A(n_8117),
.Y(n_9079)
);

AND2x4_ASAP7_75t_L g9080 ( 
.A(n_8266),
.B(n_7016),
.Y(n_9080)
);

INVx1_ASAP7_75t_L g9081 ( 
.A(n_7999),
.Y(n_9081)
);

INVx1_ASAP7_75t_L g9082 ( 
.A(n_7999),
.Y(n_9082)
);

INVx1_ASAP7_75t_L g9083 ( 
.A(n_8157),
.Y(n_9083)
);

INVx1_ASAP7_75t_L g9084 ( 
.A(n_8157),
.Y(n_9084)
);

OAI21x1_ASAP7_75t_L g9085 ( 
.A1(n_7844),
.A2(n_6659),
.B(n_7404),
.Y(n_9085)
);

NOR2xp33_ASAP7_75t_L g9086 ( 
.A(n_8075),
.B(n_6274),
.Y(n_9086)
);

INVx2_ASAP7_75t_L g9087 ( 
.A(n_7994),
.Y(n_9087)
);

INVx1_ASAP7_75t_L g9088 ( 
.A(n_7926),
.Y(n_9088)
);

INVx1_ASAP7_75t_L g9089 ( 
.A(n_7926),
.Y(n_9089)
);

INVx1_ASAP7_75t_L g9090 ( 
.A(n_7980),
.Y(n_9090)
);

OAI22xp5_ASAP7_75t_L g9091 ( 
.A1(n_7439),
.A2(n_6758),
.B1(n_7288),
.B2(n_7272),
.Y(n_9091)
);

INVx1_ASAP7_75t_L g9092 ( 
.A(n_7915),
.Y(n_9092)
);

HB1xp67_ASAP7_75t_L g9093 ( 
.A(n_8128),
.Y(n_9093)
);

INVx2_ASAP7_75t_L g9094 ( 
.A(n_7994),
.Y(n_9094)
);

INVx1_ASAP7_75t_L g9095 ( 
.A(n_7915),
.Y(n_9095)
);

AND2x2_ASAP7_75t_L g9096 ( 
.A(n_8059),
.B(n_6600),
.Y(n_9096)
);

BUFx3_ASAP7_75t_L g9097 ( 
.A(n_7682),
.Y(n_9097)
);

INVx2_ASAP7_75t_L g9098 ( 
.A(n_7996),
.Y(n_9098)
);

INVx1_ASAP7_75t_L g9099 ( 
.A(n_7919),
.Y(n_9099)
);

HB1xp67_ASAP7_75t_L g9100 ( 
.A(n_8153),
.Y(n_9100)
);

INVx3_ASAP7_75t_L g9101 ( 
.A(n_8116),
.Y(n_9101)
);

OAI21x1_ASAP7_75t_L g9102 ( 
.A1(n_7866),
.A2(n_6659),
.B(n_7404),
.Y(n_9102)
);

CKINVDCx5p33_ASAP7_75t_R g9103 ( 
.A(n_8005),
.Y(n_9103)
);

INVx1_ASAP7_75t_L g9104 ( 
.A(n_7919),
.Y(n_9104)
);

OA21x2_ASAP7_75t_L g9105 ( 
.A1(n_7719),
.A2(n_6786),
.B(n_6785),
.Y(n_9105)
);

OAI21x1_ASAP7_75t_L g9106 ( 
.A1(n_7866),
.A2(n_6659),
.B(n_6770),
.Y(n_9106)
);

AND2x2_ASAP7_75t_L g9107 ( 
.A(n_7984),
.B(n_6600),
.Y(n_9107)
);

INVx1_ASAP7_75t_L g9108 ( 
.A(n_7909),
.Y(n_9108)
);

INVx2_ASAP7_75t_L g9109 ( 
.A(n_7996),
.Y(n_9109)
);

OA21x2_ASAP7_75t_L g9110 ( 
.A1(n_7729),
.A2(n_6786),
.B(n_6785),
.Y(n_9110)
);

AO31x2_ASAP7_75t_L g9111 ( 
.A1(n_7483),
.A2(n_6471),
.A3(n_6479),
.B(n_6455),
.Y(n_9111)
);

INVx1_ASAP7_75t_L g9112 ( 
.A(n_7909),
.Y(n_9112)
);

INVx2_ASAP7_75t_L g9113 ( 
.A(n_8003),
.Y(n_9113)
);

INVx1_ASAP7_75t_L g9114 ( 
.A(n_7910),
.Y(n_9114)
);

INVxp67_ASAP7_75t_L g9115 ( 
.A(n_7545),
.Y(n_9115)
);

CKINVDCx5p33_ASAP7_75t_R g9116 ( 
.A(n_7721),
.Y(n_9116)
);

INVx2_ASAP7_75t_L g9117 ( 
.A(n_8003),
.Y(n_9117)
);

INVx1_ASAP7_75t_L g9118 ( 
.A(n_7826),
.Y(n_9118)
);

INVx1_ASAP7_75t_L g9119 ( 
.A(n_7854),
.Y(n_9119)
);

INVxp67_ASAP7_75t_SL g9120 ( 
.A(n_7575),
.Y(n_9120)
);

NOR2xp33_ASAP7_75t_L g9121 ( 
.A(n_7792),
.B(n_6275),
.Y(n_9121)
);

HB1xp67_ASAP7_75t_L g9122 ( 
.A(n_8193),
.Y(n_9122)
);

INVx1_ASAP7_75t_L g9123 ( 
.A(n_7933),
.Y(n_9123)
);

OAI22xp33_ASAP7_75t_L g9124 ( 
.A1(n_7680),
.A2(n_6843),
.B1(n_7029),
.B2(n_6882),
.Y(n_9124)
);

BUFx2_ASAP7_75t_L g9125 ( 
.A(n_8054),
.Y(n_9125)
);

INVx1_ASAP7_75t_L g9126 ( 
.A(n_7933),
.Y(n_9126)
);

BUFx3_ASAP7_75t_L g9127 ( 
.A(n_7748),
.Y(n_9127)
);

INVx1_ASAP7_75t_L g9128 ( 
.A(n_7935),
.Y(n_9128)
);

AND2x2_ASAP7_75t_L g9129 ( 
.A(n_8024),
.B(n_6600),
.Y(n_9129)
);

INVx1_ASAP7_75t_L g9130 ( 
.A(n_7935),
.Y(n_9130)
);

INVx2_ASAP7_75t_L g9131 ( 
.A(n_8061),
.Y(n_9131)
);

INVx2_ASAP7_75t_L g9132 ( 
.A(n_8061),
.Y(n_9132)
);

AND2x2_ASAP7_75t_L g9133 ( 
.A(n_8024),
.B(n_6947),
.Y(n_9133)
);

AO21x1_ASAP7_75t_L g9134 ( 
.A1(n_8283),
.A2(n_6947),
.B(n_6870),
.Y(n_9134)
);

NAND2xp5_ASAP7_75t_L g9135 ( 
.A(n_7939),
.B(n_7312),
.Y(n_9135)
);

INVx1_ASAP7_75t_L g9136 ( 
.A(n_8170),
.Y(n_9136)
);

AND2x2_ASAP7_75t_L g9137 ( 
.A(n_8126),
.B(n_8059),
.Y(n_9137)
);

INVx2_ASAP7_75t_L g9138 ( 
.A(n_8062),
.Y(n_9138)
);

INVx1_ASAP7_75t_L g9139 ( 
.A(n_8060),
.Y(n_9139)
);

INVx2_ASAP7_75t_L g9140 ( 
.A(n_8062),
.Y(n_9140)
);

INVx1_ASAP7_75t_SL g9141 ( 
.A(n_7504),
.Y(n_9141)
);

AND2x2_ASAP7_75t_L g9142 ( 
.A(n_8086),
.B(n_6646),
.Y(n_9142)
);

INVx2_ASAP7_75t_SL g9143 ( 
.A(n_8165),
.Y(n_9143)
);

INVxp67_ASAP7_75t_SL g9144 ( 
.A(n_7577),
.Y(n_9144)
);

OAI21x1_ASAP7_75t_L g9145 ( 
.A1(n_7925),
.A2(n_6770),
.B(n_7003),
.Y(n_9145)
);

AND2x4_ASAP7_75t_L g9146 ( 
.A(n_8291),
.B(n_6462),
.Y(n_9146)
);

INVx1_ASAP7_75t_L g9147 ( 
.A(n_7922),
.Y(n_9147)
);

AND2x2_ASAP7_75t_L g9148 ( 
.A(n_8086),
.B(n_8126),
.Y(n_9148)
);

INVx2_ASAP7_75t_L g9149 ( 
.A(n_8065),
.Y(n_9149)
);

INVx2_ASAP7_75t_L g9150 ( 
.A(n_8065),
.Y(n_9150)
);

AND2x2_ASAP7_75t_L g9151 ( 
.A(n_8175),
.B(n_6646),
.Y(n_9151)
);

OAI21x1_ASAP7_75t_L g9152 ( 
.A1(n_7925),
.A2(n_6770),
.B(n_7003),
.Y(n_9152)
);

INVx2_ASAP7_75t_L g9153 ( 
.A(n_8066),
.Y(n_9153)
);

INVx1_ASAP7_75t_L g9154 ( 
.A(n_7922),
.Y(n_9154)
);

CKINVDCx8_ASAP7_75t_R g9155 ( 
.A(n_7545),
.Y(n_9155)
);

OAI22xp5_ASAP7_75t_SL g9156 ( 
.A1(n_8338),
.A2(n_6705),
.B1(n_6280),
.B2(n_6284),
.Y(n_9156)
);

AND2x2_ASAP7_75t_L g9157 ( 
.A(n_8175),
.B(n_6646),
.Y(n_9157)
);

INVx1_ASAP7_75t_L g9158 ( 
.A(n_7970),
.Y(n_9158)
);

AND2x2_ASAP7_75t_L g9159 ( 
.A(n_8219),
.B(n_6646),
.Y(n_9159)
);

AND2x2_ASAP7_75t_L g9160 ( 
.A(n_8219),
.B(n_6646),
.Y(n_9160)
);

INVx1_ASAP7_75t_L g9161 ( 
.A(n_7970),
.Y(n_9161)
);

OAI21x1_ASAP7_75t_L g9162 ( 
.A1(n_8026),
.A2(n_6770),
.B(n_7003),
.Y(n_9162)
);

NAND2xp5_ASAP7_75t_L g9163 ( 
.A(n_9120),
.B(n_8102),
.Y(n_9163)
);

INVx2_ASAP7_75t_L g9164 ( 
.A(n_8491),
.Y(n_9164)
);

AO31x2_ASAP7_75t_L g9165 ( 
.A1(n_8457),
.A2(n_7492),
.A3(n_7483),
.B(n_8323),
.Y(n_9165)
);

BUFx6f_ASAP7_75t_SL g9166 ( 
.A(n_8378),
.Y(n_9166)
);

NAND2xp5_ASAP7_75t_L g9167 ( 
.A(n_9144),
.B(n_8457),
.Y(n_9167)
);

INVx2_ASAP7_75t_L g9168 ( 
.A(n_8491),
.Y(n_9168)
);

AOI22xp33_ASAP7_75t_L g9169 ( 
.A1(n_8681),
.A2(n_7700),
.B1(n_7693),
.B2(n_7422),
.Y(n_9169)
);

AND2x2_ASAP7_75t_L g9170 ( 
.A(n_8683),
.B(n_8145),
.Y(n_9170)
);

INVx1_ASAP7_75t_L g9171 ( 
.A(n_8357),
.Y(n_9171)
);

BUFx3_ASAP7_75t_L g9172 ( 
.A(n_8482),
.Y(n_9172)
);

OAI22xp5_ASAP7_75t_L g9173 ( 
.A1(n_9028),
.A2(n_7482),
.B1(n_7473),
.B2(n_7836),
.Y(n_9173)
);

AOI22xp33_ASAP7_75t_L g9174 ( 
.A1(n_8369),
.A2(n_7700),
.B1(n_7693),
.B2(n_7422),
.Y(n_9174)
);

AOI222xp33_ASAP7_75t_L g9175 ( 
.A1(n_8478),
.A2(n_8184),
.B1(n_8189),
.B2(n_8341),
.C1(n_8234),
.C2(n_8282),
.Y(n_9175)
);

OAI221xp5_ASAP7_75t_L g9176 ( 
.A1(n_8586),
.A2(n_8319),
.B1(n_8144),
.B2(n_8121),
.C(n_8341),
.Y(n_9176)
);

INVx2_ASAP7_75t_L g9177 ( 
.A(n_8815),
.Y(n_9177)
);

INVx1_ASAP7_75t_L g9178 ( 
.A(n_8376),
.Y(n_9178)
);

AOI22xp33_ASAP7_75t_SL g9179 ( 
.A1(n_8644),
.A2(n_6443),
.B1(n_7566),
.B2(n_8234),
.Y(n_9179)
);

INVx2_ASAP7_75t_L g9180 ( 
.A(n_8815),
.Y(n_9180)
);

OA21x2_ASAP7_75t_L g9181 ( 
.A1(n_8747),
.A2(n_7739),
.B(n_7729),
.Y(n_9181)
);

INVx1_ASAP7_75t_L g9182 ( 
.A(n_8472),
.Y(n_9182)
);

OR2x2_ASAP7_75t_L g9183 ( 
.A(n_8414),
.B(n_7752),
.Y(n_9183)
);

INVx1_ASAP7_75t_L g9184 ( 
.A(n_8472),
.Y(n_9184)
);

OR2x2_ASAP7_75t_L g9185 ( 
.A(n_8414),
.B(n_8432),
.Y(n_9185)
);

INVx1_ASAP7_75t_L g9186 ( 
.A(n_8474),
.Y(n_9186)
);

AO31x2_ASAP7_75t_L g9187 ( 
.A1(n_8586),
.A2(n_7492),
.A3(n_7739),
.B(n_7729),
.Y(n_9187)
);

OAI22xp5_ASAP7_75t_L g9188 ( 
.A1(n_8910),
.A2(n_7503),
.B1(n_7629),
.B2(n_7486),
.Y(n_9188)
);

OAI22xp33_ASAP7_75t_L g9189 ( 
.A1(n_8605),
.A2(n_7680),
.B1(n_7704),
.B2(n_7488),
.Y(n_9189)
);

AOI22xp5_ASAP7_75t_L g9190 ( 
.A1(n_8426),
.A2(n_8908),
.B1(n_8741),
.B2(n_8846),
.Y(n_9190)
);

OR2x2_ASAP7_75t_L g9191 ( 
.A(n_8432),
.B(n_7508),
.Y(n_9191)
);

INVx1_ASAP7_75t_L g9192 ( 
.A(n_8473),
.Y(n_9192)
);

OR2x2_ASAP7_75t_L g9193 ( 
.A(n_8513),
.B(n_7508),
.Y(n_9193)
);

AOI221xp5_ASAP7_75t_L g9194 ( 
.A1(n_8441),
.A2(n_7986),
.B1(n_8189),
.B2(n_8184),
.C(n_7426),
.Y(n_9194)
);

AOI22xp33_ASAP7_75t_L g9195 ( 
.A1(n_8417),
.A2(n_7700),
.B1(n_7693),
.B2(n_7422),
.Y(n_9195)
);

OAI211xp5_ASAP7_75t_SL g9196 ( 
.A1(n_9020),
.A2(n_8116),
.B(n_8237),
.C(n_8188),
.Y(n_9196)
);

AOI22xp33_ASAP7_75t_SL g9197 ( 
.A1(n_8753),
.A2(n_7566),
.B1(n_8282),
.B2(n_8245),
.Y(n_9197)
);

AOI21xp33_ASAP7_75t_L g9198 ( 
.A1(n_8735),
.A2(n_8427),
.B(n_8389),
.Y(n_9198)
);

AOI222xp33_ASAP7_75t_L g9199 ( 
.A1(n_8368),
.A2(n_8245),
.B1(n_8299),
.B2(n_7492),
.C1(n_7727),
.C2(n_7739),
.Y(n_9199)
);

OAI221xp5_ASAP7_75t_L g9200 ( 
.A1(n_8665),
.A2(n_8289),
.B1(n_8217),
.B2(n_7965),
.C(n_7998),
.Y(n_9200)
);

INVx2_ASAP7_75t_L g9201 ( 
.A(n_8683),
.Y(n_9201)
);

NOR2x1_ASAP7_75t_R g9202 ( 
.A(n_8482),
.B(n_7748),
.Y(n_9202)
);

AOI221xp5_ASAP7_75t_L g9203 ( 
.A1(n_8402),
.A2(n_8250),
.B1(n_8237),
.B2(n_8188),
.C(n_8066),
.Y(n_9203)
);

AND2x2_ASAP7_75t_L g9204 ( 
.A(n_8865),
.B(n_8145),
.Y(n_9204)
);

HB1xp67_ASAP7_75t_L g9205 ( 
.A(n_8452),
.Y(n_9205)
);

INVx1_ASAP7_75t_L g9206 ( 
.A(n_8474),
.Y(n_9206)
);

AND2x2_ASAP7_75t_L g9207 ( 
.A(n_8865),
.B(n_8145),
.Y(n_9207)
);

AO21x2_ASAP7_75t_L g9208 ( 
.A1(n_8692),
.A2(n_7495),
.B(n_7961),
.Y(n_9208)
);

AO21x2_ASAP7_75t_L g9209 ( 
.A1(n_9037),
.A2(n_7495),
.B(n_7961),
.Y(n_9209)
);

AOI22xp33_ASAP7_75t_SL g9210 ( 
.A1(n_8355),
.A2(n_7566),
.B1(n_8299),
.B2(n_8237),
.Y(n_9210)
);

INVx1_ASAP7_75t_L g9211 ( 
.A(n_8611),
.Y(n_9211)
);

INVx2_ASAP7_75t_L g9212 ( 
.A(n_8461),
.Y(n_9212)
);

AOI222xp33_ASAP7_75t_L g9213 ( 
.A1(n_8908),
.A2(n_8495),
.B1(n_8361),
.B2(n_8366),
.C1(n_8371),
.C2(n_8355),
.Y(n_9213)
);

OAI221xp5_ASAP7_75t_L g9214 ( 
.A1(n_8547),
.A2(n_7661),
.B1(n_7650),
.B2(n_7686),
.C(n_7566),
.Y(n_9214)
);

OR2x2_ASAP7_75t_L g9215 ( 
.A(n_8592),
.B(n_8262),
.Y(n_9215)
);

AND2x4_ASAP7_75t_L g9216 ( 
.A(n_8871),
.B(n_7829),
.Y(n_9216)
);

INVx1_ASAP7_75t_L g9217 ( 
.A(n_8473),
.Y(n_9217)
);

OAI22xp33_ASAP7_75t_L g9218 ( 
.A1(n_8733),
.A2(n_7704),
.B1(n_7488),
.B2(n_7422),
.Y(n_9218)
);

OAI211xp5_ASAP7_75t_L g9219 ( 
.A1(n_8562),
.A2(n_7840),
.B(n_7819),
.C(n_8295),
.Y(n_9219)
);

NAND2xp5_ASAP7_75t_L g9220 ( 
.A(n_8767),
.B(n_7946),
.Y(n_9220)
);

OAI21xp33_ASAP7_75t_SL g9221 ( 
.A1(n_8931),
.A2(n_8237),
.B(n_8188),
.Y(n_9221)
);

AO31x2_ASAP7_75t_L g9222 ( 
.A1(n_8702),
.A2(n_7501),
.A3(n_7507),
.B(n_7496),
.Y(n_9222)
);

AOI22xp33_ASAP7_75t_L g9223 ( 
.A1(n_8367),
.A2(n_7700),
.B1(n_7693),
.B2(n_7422),
.Y(n_9223)
);

AOI222xp33_ASAP7_75t_L g9224 ( 
.A1(n_8361),
.A2(n_8371),
.B1(n_8366),
.B2(n_8465),
.C1(n_8448),
.C2(n_8493),
.Y(n_9224)
);

INVx1_ASAP7_75t_L g9225 ( 
.A(n_8612),
.Y(n_9225)
);

INVx2_ASAP7_75t_L g9226 ( 
.A(n_8461),
.Y(n_9226)
);

AOI22xp33_ASAP7_75t_L g9227 ( 
.A1(n_8367),
.A2(n_7700),
.B1(n_7693),
.B2(n_7495),
.Y(n_9227)
);

INVx2_ASAP7_75t_L g9228 ( 
.A(n_8507),
.Y(n_9228)
);

INVx1_ASAP7_75t_L g9229 ( 
.A(n_8611),
.Y(n_9229)
);

INVx3_ASAP7_75t_L g9230 ( 
.A(n_8453),
.Y(n_9230)
);

INVx2_ASAP7_75t_L g9231 ( 
.A(n_8507),
.Y(n_9231)
);

OAI22xp5_ASAP7_75t_L g9232 ( 
.A1(n_8792),
.A2(n_7503),
.B1(n_7494),
.B2(n_7497),
.Y(n_9232)
);

AOI22xp33_ASAP7_75t_L g9233 ( 
.A1(n_8367),
.A2(n_7819),
.B1(n_6644),
.B2(n_8051),
.Y(n_9233)
);

INVx2_ASAP7_75t_L g9234 ( 
.A(n_8581),
.Y(n_9234)
);

AOI22xp5_ASAP7_75t_L g9235 ( 
.A1(n_9134),
.A2(n_8769),
.B1(n_8416),
.B2(n_8556),
.Y(n_9235)
);

OAI22xp5_ASAP7_75t_L g9236 ( 
.A1(n_9051),
.A2(n_8168),
.B1(n_8104),
.B2(n_7879),
.Y(n_9236)
);

AOI22xp33_ASAP7_75t_L g9237 ( 
.A1(n_9134),
.A2(n_7819),
.B1(n_6644),
.B2(n_8051),
.Y(n_9237)
);

INVx1_ASAP7_75t_L g9238 ( 
.A(n_8612),
.Y(n_9238)
);

AOI22xp33_ASAP7_75t_L g9239 ( 
.A1(n_8931),
.A2(n_7819),
.B1(n_6644),
.B2(n_8051),
.Y(n_9239)
);

OAI221xp5_ASAP7_75t_L g9240 ( 
.A1(n_8928),
.A2(n_8100),
.B1(n_8034),
.B2(n_7941),
.C(n_7917),
.Y(n_9240)
);

NAND2xp5_ASAP7_75t_L g9241 ( 
.A(n_8610),
.B(n_7962),
.Y(n_9241)
);

OR2x2_ASAP7_75t_L g9242 ( 
.A(n_8598),
.B(n_8538),
.Y(n_9242)
);

AO21x1_ASAP7_75t_SL g9243 ( 
.A1(n_8386),
.A2(n_8081),
.B(n_7354),
.Y(n_9243)
);

AOI22xp33_ASAP7_75t_L g9244 ( 
.A1(n_8442),
.A2(n_6644),
.B1(n_7493),
.B2(n_7517),
.Y(n_9244)
);

NAND2xp5_ASAP7_75t_L g9245 ( 
.A(n_8435),
.B(n_8002),
.Y(n_9245)
);

INVx1_ASAP7_75t_L g9246 ( 
.A(n_8613),
.Y(n_9246)
);

NAND3xp33_ASAP7_75t_L g9247 ( 
.A(n_8972),
.B(n_8541),
.C(n_8476),
.Y(n_9247)
);

INVx1_ASAP7_75t_L g9248 ( 
.A(n_8613),
.Y(n_9248)
);

OAI221xp5_ASAP7_75t_L g9249 ( 
.A1(n_9048),
.A2(n_7750),
.B1(n_8235),
.B2(n_8263),
.C(n_8238),
.Y(n_9249)
);

INVx1_ASAP7_75t_L g9250 ( 
.A(n_8614),
.Y(n_9250)
);

OAI21xp33_ASAP7_75t_L g9251 ( 
.A1(n_9135),
.A2(n_8135),
.B(n_8125),
.Y(n_9251)
);

NAND2xp5_ASAP7_75t_L g9252 ( 
.A(n_8450),
.B(n_8038),
.Y(n_9252)
);

INVx1_ASAP7_75t_L g9253 ( 
.A(n_8614),
.Y(n_9253)
);

OAI22xp33_ASAP7_75t_L g9254 ( 
.A1(n_8887),
.A2(n_8032),
.B1(n_8058),
.B2(n_7628),
.Y(n_9254)
);

AND2x4_ASAP7_75t_L g9255 ( 
.A(n_8871),
.B(n_7829),
.Y(n_9255)
);

BUFx8_ASAP7_75t_L g9256 ( 
.A(n_8881),
.Y(n_9256)
);

AOI22xp33_ASAP7_75t_L g9257 ( 
.A1(n_8541),
.A2(n_7519),
.B1(n_7715),
.B2(n_7717),
.Y(n_9257)
);

AO31x2_ASAP7_75t_L g9258 ( 
.A1(n_8698),
.A2(n_7501),
.A3(n_7507),
.B(n_7496),
.Y(n_9258)
);

INVx5_ASAP7_75t_SL g9259 ( 
.A(n_8470),
.Y(n_9259)
);

OAI21x1_ASAP7_75t_L g9260 ( 
.A1(n_8688),
.A2(n_7736),
.B(n_8026),
.Y(n_9260)
);

AOI221xp5_ASAP7_75t_L g9261 ( 
.A1(n_8544),
.A2(n_8250),
.B1(n_8188),
.B2(n_8087),
.C(n_8092),
.Y(n_9261)
);

AND2x2_ASAP7_75t_L g9262 ( 
.A(n_8903),
.B(n_8232),
.Y(n_9262)
);

AND2x2_ASAP7_75t_L g9263 ( 
.A(n_8903),
.B(n_8232),
.Y(n_9263)
);

AOI22xp33_ASAP7_75t_L g9264 ( 
.A1(n_8541),
.A2(n_7467),
.B1(n_7536),
.B2(n_7524),
.Y(n_9264)
);

AOI22xp33_ASAP7_75t_L g9265 ( 
.A1(n_8430),
.A2(n_7599),
.B1(n_7576),
.B2(n_7768),
.Y(n_9265)
);

AOI21xp33_ASAP7_75t_L g9266 ( 
.A1(n_8477),
.A2(n_7840),
.B(n_7699),
.Y(n_9266)
);

AOI21xp5_ASAP7_75t_L g9267 ( 
.A1(n_9124),
.A2(n_8147),
.B(n_7608),
.Y(n_9267)
);

AOI22xp33_ASAP7_75t_L g9268 ( 
.A1(n_8985),
.A2(n_7850),
.B1(n_6616),
.B2(n_7840),
.Y(n_9268)
);

OAI22xp5_ASAP7_75t_L g9269 ( 
.A1(n_8986),
.A2(n_7876),
.B1(n_7621),
.B2(n_7430),
.Y(n_9269)
);

INVx1_ASAP7_75t_L g9270 ( 
.A(n_8984),
.Y(n_9270)
);

BUFx6f_ASAP7_75t_L g9271 ( 
.A(n_8540),
.Y(n_9271)
);

AOI222xp33_ASAP7_75t_L g9272 ( 
.A1(n_9043),
.A2(n_7316),
.B1(n_8250),
.B2(n_7961),
.C1(n_7973),
.C2(n_7967),
.Y(n_9272)
);

INVx3_ASAP7_75t_L g9273 ( 
.A(n_8453),
.Y(n_9273)
);

OAI22xp5_ASAP7_75t_L g9274 ( 
.A1(n_8976),
.A2(n_8339),
.B1(n_8307),
.B2(n_7648),
.Y(n_9274)
);

OAI22xp5_ASAP7_75t_L g9275 ( 
.A1(n_9091),
.A2(n_7459),
.B1(n_7751),
.B2(n_7502),
.Y(n_9275)
);

OAI22xp5_ASAP7_75t_L g9276 ( 
.A1(n_8860),
.A2(n_7751),
.B1(n_7646),
.B2(n_7927),
.Y(n_9276)
);

NAND2xp5_ASAP7_75t_L g9277 ( 
.A(n_8454),
.B(n_8198),
.Y(n_9277)
);

AOI22xp33_ASAP7_75t_L g9278 ( 
.A1(n_8769),
.A2(n_6616),
.B1(n_7840),
.B2(n_7208),
.Y(n_9278)
);

AOI22xp33_ASAP7_75t_L g9279 ( 
.A1(n_8769),
.A2(n_6616),
.B1(n_7208),
.B2(n_7852),
.Y(n_9279)
);

INVx1_ASAP7_75t_L g9280 ( 
.A(n_8616),
.Y(n_9280)
);

AND2x2_ASAP7_75t_L g9281 ( 
.A(n_8757),
.B(n_8232),
.Y(n_9281)
);

OAI22xp5_ASAP7_75t_L g9282 ( 
.A1(n_8648),
.A2(n_7642),
.B1(n_7681),
.B2(n_7873),
.Y(n_9282)
);

INVx2_ASAP7_75t_L g9283 ( 
.A(n_8581),
.Y(n_9283)
);

OA21x2_ASAP7_75t_L g9284 ( 
.A1(n_8747),
.A2(n_8419),
.B(n_8392),
.Y(n_9284)
);

OR2x6_ASAP7_75t_L g9285 ( 
.A(n_8830),
.B(n_7863),
.Y(n_9285)
);

OAI221xp5_ASAP7_75t_L g9286 ( 
.A1(n_8562),
.A2(n_8250),
.B1(n_8091),
.B2(n_8092),
.C(n_8087),
.Y(n_9286)
);

INVx1_ASAP7_75t_L g9287 ( 
.A(n_8616),
.Y(n_9287)
);

AND2x2_ASAP7_75t_L g9288 ( 
.A(n_8757),
.B(n_8256),
.Y(n_9288)
);

NAND3xp33_ASAP7_75t_L g9289 ( 
.A(n_8477),
.B(n_8351),
.C(n_7049),
.Y(n_9289)
);

OR2x2_ASAP7_75t_L g9290 ( 
.A(n_8720),
.B(n_8262),
.Y(n_9290)
);

AO31x2_ASAP7_75t_L g9291 ( 
.A1(n_8702),
.A2(n_7501),
.A3(n_7507),
.B(n_7496),
.Y(n_9291)
);

AOI221xp5_ASAP7_75t_L g9292 ( 
.A1(n_8955),
.A2(n_8139),
.B1(n_8150),
.B2(n_8091),
.C(n_8069),
.Y(n_9292)
);

INVxp67_ASAP7_75t_L g9293 ( 
.A(n_8774),
.Y(n_9293)
);

OAI221xp5_ASAP7_75t_L g9294 ( 
.A1(n_8648),
.A2(n_8150),
.B1(n_8152),
.B2(n_8139),
.C(n_8069),
.Y(n_9294)
);

INVx2_ASAP7_75t_SL g9295 ( 
.A(n_8540),
.Y(n_9295)
);

INVx2_ASAP7_75t_L g9296 ( 
.A(n_9025),
.Y(n_9296)
);

AOI22xp33_ASAP7_75t_L g9297 ( 
.A1(n_8477),
.A2(n_6616),
.B1(n_7208),
.B2(n_7853),
.Y(n_9297)
);

INVx2_ASAP7_75t_L g9298 ( 
.A(n_9025),
.Y(n_9298)
);

OAI22xp5_ASAP7_75t_L g9299 ( 
.A1(n_8729),
.A2(n_7857),
.B1(n_8292),
.B2(n_8290),
.Y(n_9299)
);

AND2x2_ASAP7_75t_L g9300 ( 
.A(n_8757),
.B(n_8256),
.Y(n_9300)
);

AND2x2_ASAP7_75t_L g9301 ( 
.A(n_8757),
.B(n_8256),
.Y(n_9301)
);

AND2x2_ASAP7_75t_L g9302 ( 
.A(n_8936),
.B(n_7829),
.Y(n_9302)
);

NAND2xp5_ASAP7_75t_L g9303 ( 
.A(n_8709),
.B(n_7924),
.Y(n_9303)
);

OAI22xp5_ASAP7_75t_L g9304 ( 
.A1(n_8729),
.A2(n_8195),
.B1(n_8196),
.B2(n_8191),
.Y(n_9304)
);

OAI22xp5_ASAP7_75t_L g9305 ( 
.A1(n_8783),
.A2(n_8233),
.B1(n_7124),
.B2(n_7582),
.Y(n_9305)
);

AOI22xp33_ASAP7_75t_SL g9306 ( 
.A1(n_8696),
.A2(n_7152),
.B1(n_6603),
.B2(n_6616),
.Y(n_9306)
);

AOI221xp5_ASAP7_75t_L g9307 ( 
.A1(n_8945),
.A2(n_8760),
.B1(n_8778),
.B2(n_8732),
.C(n_8696),
.Y(n_9307)
);

OAI22xp5_ASAP7_75t_L g9308 ( 
.A1(n_8783),
.A2(n_7124),
.B1(n_7877),
.B2(n_7389),
.Y(n_9308)
);

INVx2_ASAP7_75t_L g9309 ( 
.A(n_9015),
.Y(n_9309)
);

BUFx8_ASAP7_75t_SL g9310 ( 
.A(n_8649),
.Y(n_9310)
);

OAI211xp5_ASAP7_75t_L g9311 ( 
.A1(n_9155),
.A2(n_8295),
.B(n_8351),
.C(n_8112),
.Y(n_9311)
);

AND2x2_ASAP7_75t_L g9312 ( 
.A(n_8936),
.B(n_7914),
.Y(n_9312)
);

AO21x2_ASAP7_75t_L g9313 ( 
.A1(n_8698),
.A2(n_7973),
.B(n_7967),
.Y(n_9313)
);

AOI22xp33_ASAP7_75t_L g9314 ( 
.A1(n_8535),
.A2(n_7208),
.B1(n_7637),
.B2(n_7723),
.Y(n_9314)
);

AOI21xp33_ASAP7_75t_L g9315 ( 
.A1(n_8535),
.A2(n_7699),
.B(n_7676),
.Y(n_9315)
);

INVx5_ASAP7_75t_SL g9316 ( 
.A(n_8571),
.Y(n_9316)
);

OAI21xp5_ASAP7_75t_SL g9317 ( 
.A1(n_8808),
.A2(n_7893),
.B(n_7336),
.Y(n_9317)
);

INVx2_ASAP7_75t_L g9318 ( 
.A(n_9015),
.Y(n_9318)
);

AOI221xp5_ASAP7_75t_L g9319 ( 
.A1(n_8696),
.A2(n_8222),
.B1(n_8223),
.B2(n_8163),
.C(n_8152),
.Y(n_9319)
);

INVx4_ASAP7_75t_L g9320 ( 
.A(n_8378),
.Y(n_9320)
);

AND2x2_ASAP7_75t_L g9321 ( 
.A(n_9049),
.B(n_7914),
.Y(n_9321)
);

OAI22xp5_ASAP7_75t_L g9322 ( 
.A1(n_8712),
.A2(n_7389),
.B1(n_8015),
.B2(n_7029),
.Y(n_9322)
);

OAI21xp5_ASAP7_75t_L g9323 ( 
.A1(n_8585),
.A2(n_8286),
.B(n_6696),
.Y(n_9323)
);

AOI22xp5_ASAP7_75t_L g9324 ( 
.A1(n_8536),
.A2(n_6840),
.B1(n_7316),
.B2(n_7944),
.Y(n_9324)
);

AOI22xp33_ASAP7_75t_L g9325 ( 
.A1(n_8535),
.A2(n_8348),
.B1(n_8318),
.B2(n_6653),
.Y(n_9325)
);

OAI211xp5_ASAP7_75t_L g9326 ( 
.A1(n_9155),
.A2(n_8136),
.B(n_8209),
.C(n_8112),
.Y(n_9326)
);

INVx1_ASAP7_75t_L g9327 ( 
.A(n_8991),
.Y(n_9327)
);

AOI22xp33_ASAP7_75t_L g9328 ( 
.A1(n_8536),
.A2(n_8348),
.B1(n_8318),
.B2(n_6653),
.Y(n_9328)
);

AND2x2_ASAP7_75t_L g9329 ( 
.A(n_9049),
.B(n_9125),
.Y(n_9329)
);

AND2x2_ASAP7_75t_L g9330 ( 
.A(n_9125),
.B(n_7914),
.Y(n_9330)
);

AOI22xp33_ASAP7_75t_L g9331 ( 
.A1(n_8536),
.A2(n_6653),
.B1(n_8222),
.B2(n_8163),
.Y(n_9331)
);

OAI22xp5_ASAP7_75t_L g9332 ( 
.A1(n_8859),
.A2(n_7688),
.B1(n_8261),
.B2(n_8214),
.Y(n_9332)
);

AOI21xp5_ASAP7_75t_L g9333 ( 
.A1(n_8489),
.A2(n_8147),
.B(n_7505),
.Y(n_9333)
);

AND2x2_ASAP7_75t_L g9334 ( 
.A(n_8520),
.B(n_8291),
.Y(n_9334)
);

INVx1_ASAP7_75t_L g9335 ( 
.A(n_8984),
.Y(n_9335)
);

INVx1_ASAP7_75t_L g9336 ( 
.A(n_8991),
.Y(n_9336)
);

AND2x2_ASAP7_75t_L g9337 ( 
.A(n_8520),
.B(n_8291),
.Y(n_9337)
);

OAI221xp5_ASAP7_75t_L g9338 ( 
.A1(n_8732),
.A2(n_8227),
.B1(n_8244),
.B2(n_8236),
.C(n_8223),
.Y(n_9338)
);

AOI22xp33_ASAP7_75t_L g9339 ( 
.A1(n_9146),
.A2(n_6653),
.B1(n_8236),
.B2(n_8227),
.Y(n_9339)
);

AO21x2_ASAP7_75t_L g9340 ( 
.A1(n_8392),
.A2(n_7973),
.B(n_7967),
.Y(n_9340)
);

AND2x2_ASAP7_75t_L g9341 ( 
.A(n_8452),
.B(n_7885),
.Y(n_9341)
);

AOI22xp33_ASAP7_75t_L g9342 ( 
.A1(n_9146),
.A2(n_6653),
.B1(n_8264),
.B2(n_8244),
.Y(n_9342)
);

OAI221xp5_ASAP7_75t_L g9343 ( 
.A1(n_8732),
.A2(n_8301),
.B1(n_8316),
.B2(n_8305),
.C(n_8264),
.Y(n_9343)
);

OAI22xp33_ASAP7_75t_L g9344 ( 
.A1(n_8760),
.A2(n_6740),
.B1(n_6870),
.B2(n_8225),
.Y(n_9344)
);

AOI22xp33_ASAP7_75t_L g9345 ( 
.A1(n_9146),
.A2(n_6653),
.B1(n_8305),
.B2(n_8301),
.Y(n_9345)
);

OAI211xp5_ASAP7_75t_SL g9346 ( 
.A1(n_8377),
.A2(n_8220),
.B(n_8007),
.C(n_7976),
.Y(n_9346)
);

OAI22xp33_ASAP7_75t_L g9347 ( 
.A1(n_8760),
.A2(n_8798),
.B1(n_8812),
.B2(n_8778),
.Y(n_9347)
);

OR2x2_ASAP7_75t_L g9348 ( 
.A(n_8720),
.B(n_7956),
.Y(n_9348)
);

OAI33xp33_ASAP7_75t_L g9349 ( 
.A1(n_8863),
.A2(n_9115),
.A3(n_8739),
.B1(n_8521),
.B2(n_9040),
.B3(n_8994),
.Y(n_9349)
);

AND2x2_ASAP7_75t_L g9350 ( 
.A(n_8632),
.B(n_7885),
.Y(n_9350)
);

BUFx6f_ASAP7_75t_L g9351 ( 
.A(n_8668),
.Y(n_9351)
);

AOI22xp33_ASAP7_75t_L g9352 ( 
.A1(n_8980),
.A2(n_6653),
.B1(n_8316),
.B2(n_6728),
.Y(n_9352)
);

INVx1_ASAP7_75t_L g9353 ( 
.A(n_8993),
.Y(n_9353)
);

OAI22xp5_ASAP7_75t_L g9354 ( 
.A1(n_8632),
.A2(n_8214),
.B1(n_8261),
.B2(n_7890),
.Y(n_9354)
);

OAI22xp5_ASAP7_75t_L g9355 ( 
.A1(n_8660),
.A2(n_7156),
.B1(n_6726),
.B2(n_7891),
.Y(n_9355)
);

AOI22xp33_ASAP7_75t_L g9356 ( 
.A1(n_8980),
.A2(n_6653),
.B1(n_6728),
.B2(n_6719),
.Y(n_9356)
);

AOI22xp33_ASAP7_75t_L g9357 ( 
.A1(n_8704),
.A2(n_6728),
.B1(n_6719),
.B2(n_7747),
.Y(n_9357)
);

AOI21xp33_ASAP7_75t_L g9358 ( 
.A1(n_8399),
.A2(n_7699),
.B(n_7676),
.Y(n_9358)
);

AO31x2_ASAP7_75t_L g9359 ( 
.A1(n_9026),
.A2(n_7587),
.A3(n_7512),
.B(n_7793),
.Y(n_9359)
);

NAND2xp5_ASAP7_75t_L g9360 ( 
.A(n_8654),
.B(n_7952),
.Y(n_9360)
);

AO31x2_ASAP7_75t_L g9361 ( 
.A1(n_9026),
.A2(n_7587),
.A3(n_7512),
.B(n_7793),
.Y(n_9361)
);

AND2x2_ASAP7_75t_L g9362 ( 
.A(n_8660),
.B(n_7885),
.Y(n_9362)
);

HB1xp67_ASAP7_75t_L g9363 ( 
.A(n_8537),
.Y(n_9363)
);

INVx2_ASAP7_75t_L g9364 ( 
.A(n_8669),
.Y(n_9364)
);

BUFx2_ASAP7_75t_SL g9365 ( 
.A(n_8649),
.Y(n_9365)
);

INVx1_ASAP7_75t_L g9366 ( 
.A(n_8993),
.Y(n_9366)
);

AND2x2_ASAP7_75t_L g9367 ( 
.A(n_8669),
.B(n_7885),
.Y(n_9367)
);

INVx1_ASAP7_75t_L g9368 ( 
.A(n_9000),
.Y(n_9368)
);

AOI21xp33_ASAP7_75t_L g9369 ( 
.A1(n_8399),
.A2(n_7699),
.B(n_7676),
.Y(n_9369)
);

BUFx2_ASAP7_75t_L g9370 ( 
.A(n_8881),
.Y(n_9370)
);

AOI221xp5_ASAP7_75t_L g9371 ( 
.A1(n_8778),
.A2(n_7432),
.B1(n_7429),
.B2(n_7428),
.C(n_7447),
.Y(n_9371)
);

AOI22xp5_ASAP7_75t_L g9372 ( 
.A1(n_8381),
.A2(n_6863),
.B1(n_7312),
.B2(n_6696),
.Y(n_9372)
);

AND2x2_ASAP7_75t_L g9373 ( 
.A(n_8679),
.B(n_8013),
.Y(n_9373)
);

AOI21xp5_ASAP7_75t_L g9374 ( 
.A1(n_8721),
.A2(n_7947),
.B(n_8328),
.Y(n_9374)
);

BUFx4f_ASAP7_75t_SL g9375 ( 
.A(n_8381),
.Y(n_9375)
);

OAI21xp33_ASAP7_75t_L g9376 ( 
.A1(n_8517),
.A2(n_7183),
.B(n_7170),
.Y(n_9376)
);

AOI21xp5_ASAP7_75t_L g9377 ( 
.A1(n_8486),
.A2(n_7156),
.B(n_8190),
.Y(n_9377)
);

OAI22xp5_ASAP7_75t_L g9378 ( 
.A1(n_8679),
.A2(n_6726),
.B1(n_7901),
.B2(n_8044),
.Y(n_9378)
);

INVx1_ASAP7_75t_L g9379 ( 
.A(n_9000),
.Y(n_9379)
);

INVx2_ASAP7_75t_L g9380 ( 
.A(n_9141),
.Y(n_9380)
);

BUFx6f_ASAP7_75t_L g9381 ( 
.A(n_8668),
.Y(n_9381)
);

NAND2x1_ASAP7_75t_L g9382 ( 
.A(n_8656),
.B(n_8190),
.Y(n_9382)
);

AOI22xp33_ASAP7_75t_L g9383 ( 
.A1(n_8704),
.A2(n_6728),
.B1(n_6719),
.B2(n_7747),
.Y(n_9383)
);

OA21x2_ASAP7_75t_L g9384 ( 
.A1(n_8419),
.A2(n_7587),
.B(n_7512),
.Y(n_9384)
);

AND2x2_ASAP7_75t_L g9385 ( 
.A(n_8923),
.B(n_8935),
.Y(n_9385)
);

OAI22xp5_ASAP7_75t_L g9386 ( 
.A1(n_8637),
.A2(n_7183),
.B1(n_7170),
.B2(n_8165),
.Y(n_9386)
);

OAI22xp5_ASAP7_75t_L g9387 ( 
.A1(n_8637),
.A2(n_8165),
.B1(n_7554),
.B2(n_7551),
.Y(n_9387)
);

AND2x2_ASAP7_75t_L g9388 ( 
.A(n_8923),
.B(n_8013),
.Y(n_9388)
);

AOI22xp33_ASAP7_75t_L g9389 ( 
.A1(n_8704),
.A2(n_6728),
.B1(n_6719),
.B2(n_7747),
.Y(n_9389)
);

CKINVDCx14_ASAP7_75t_R g9390 ( 
.A(n_8387),
.Y(n_9390)
);

NAND2xp5_ASAP7_75t_L g9391 ( 
.A(n_8654),
.B(n_7553),
.Y(n_9391)
);

AOI22xp33_ASAP7_75t_L g9392 ( 
.A1(n_8798),
.A2(n_6719),
.B1(n_7756),
.B2(n_7754),
.Y(n_9392)
);

INVx2_ASAP7_75t_L g9393 ( 
.A(n_8595),
.Y(n_9393)
);

AOI221xp5_ASAP7_75t_L g9394 ( 
.A1(n_8798),
.A2(n_7428),
.B1(n_7432),
.B2(n_7429),
.C(n_7447),
.Y(n_9394)
);

INVx1_ASAP7_75t_L g9395 ( 
.A(n_9004),
.Y(n_9395)
);

AOI22xp33_ASAP7_75t_L g9396 ( 
.A1(n_8812),
.A2(n_7756),
.B1(n_7773),
.B2(n_7754),
.Y(n_9396)
);

AOI22xp33_ASAP7_75t_SL g9397 ( 
.A1(n_8812),
.A2(n_6603),
.B1(n_7049),
.B2(n_6813),
.Y(n_9397)
);

AND2x2_ASAP7_75t_L g9398 ( 
.A(n_8935),
.B(n_8013),
.Y(n_9398)
);

AOI21xp5_ASAP7_75t_L g9399 ( 
.A1(n_8603),
.A2(n_7053),
.B(n_7162),
.Y(n_9399)
);

AOI21xp33_ASAP7_75t_L g9400 ( 
.A1(n_8399),
.A2(n_7676),
.B(n_7904),
.Y(n_9400)
);

AOI221xp5_ASAP7_75t_L g9401 ( 
.A1(n_8834),
.A2(n_7428),
.B1(n_7432),
.B2(n_7429),
.C(n_7904),
.Y(n_9401)
);

AOI22xp33_ASAP7_75t_L g9402 ( 
.A1(n_8834),
.A2(n_7756),
.B1(n_7773),
.B2(n_7754),
.Y(n_9402)
);

INVx1_ASAP7_75t_L g9403 ( 
.A(n_9004),
.Y(n_9403)
);

INVx1_ASAP7_75t_L g9404 ( 
.A(n_8358),
.Y(n_9404)
);

AOI221xp5_ASAP7_75t_L g9405 ( 
.A1(n_8834),
.A2(n_7904),
.B1(n_8240),
.B2(n_7957),
.C(n_8337),
.Y(n_9405)
);

OAI22xp33_ASAP7_75t_L g9406 ( 
.A1(n_8835),
.A2(n_6740),
.B1(n_6815),
.B2(n_7398),
.Y(n_9406)
);

AOI22xp33_ASAP7_75t_L g9407 ( 
.A1(n_8835),
.A2(n_7777),
.B1(n_7773),
.B2(n_7793),
.Y(n_9407)
);

OAI22xp5_ASAP7_75t_L g9408 ( 
.A1(n_8637),
.A2(n_8165),
.B1(n_8021),
.B2(n_8020),
.Y(n_9408)
);

INVx1_ASAP7_75t_L g9409 ( 
.A(n_8360),
.Y(n_9409)
);

AOI22xp33_ASAP7_75t_L g9410 ( 
.A1(n_8835),
.A2(n_7777),
.B1(n_7806),
.B2(n_7797),
.Y(n_9410)
);

OR2x6_ASAP7_75t_L g9411 ( 
.A(n_8830),
.B(n_8734),
.Y(n_9411)
);

OAI211xp5_ASAP7_75t_L g9412 ( 
.A1(n_8602),
.A2(n_8112),
.B(n_8209),
.C(n_8136),
.Y(n_9412)
);

AOI22xp5_ASAP7_75t_L g9413 ( 
.A1(n_8601),
.A2(n_6863),
.B1(n_7049),
.B2(n_6858),
.Y(n_9413)
);

AOI21xp33_ASAP7_75t_L g9414 ( 
.A1(n_8643),
.A2(n_8136),
.B(n_8112),
.Y(n_9414)
);

AOI22xp33_ASAP7_75t_L g9415 ( 
.A1(n_8603),
.A2(n_8680),
.B1(n_8740),
.B2(n_8451),
.Y(n_9415)
);

AOI22xp33_ASAP7_75t_L g9416 ( 
.A1(n_8603),
.A2(n_7777),
.B1(n_7806),
.B2(n_7797),
.Y(n_9416)
);

BUFx3_ASAP7_75t_L g9417 ( 
.A(n_8514),
.Y(n_9417)
);

AOI22xp5_ASAP7_75t_L g9418 ( 
.A1(n_8618),
.A2(n_7049),
.B1(n_6858),
.B2(n_7559),
.Y(n_9418)
);

AND2x2_ASAP7_75t_L g9419 ( 
.A(n_8451),
.B(n_8013),
.Y(n_9419)
);

AOI22xp33_ASAP7_75t_L g9420 ( 
.A1(n_8680),
.A2(n_7806),
.B1(n_7817),
.B2(n_7797),
.Y(n_9420)
);

OR2x2_ASAP7_75t_L g9421 ( 
.A(n_8517),
.B(n_7956),
.Y(n_9421)
);

OAI22xp5_ASAP7_75t_L g9422 ( 
.A1(n_8643),
.A2(n_7753),
.B1(n_7860),
.B2(n_7588),
.Y(n_9422)
);

AOI221xp5_ASAP7_75t_L g9423 ( 
.A1(n_8643),
.A2(n_7957),
.B1(n_8337),
.B2(n_7817),
.C(n_7842),
.Y(n_9423)
);

BUFx2_ASAP7_75t_L g9424 ( 
.A(n_8455),
.Y(n_9424)
);

INVx1_ASAP7_75t_L g9425 ( 
.A(n_8362),
.Y(n_9425)
);

AOI221xp5_ASAP7_75t_L g9426 ( 
.A1(n_8690),
.A2(n_8337),
.B1(n_7817),
.B2(n_7842),
.C(n_7834),
.Y(n_9426)
);

AOI22xp33_ASAP7_75t_L g9427 ( 
.A1(n_8680),
.A2(n_7834),
.B1(n_7842),
.B2(n_7818),
.Y(n_9427)
);

BUFx6f_ASAP7_75t_L g9428 ( 
.A(n_8383),
.Y(n_9428)
);

OAI22xp5_ASAP7_75t_L g9429 ( 
.A1(n_8635),
.A2(n_7753),
.B1(n_7860),
.B2(n_7588),
.Y(n_9429)
);

BUFx3_ASAP7_75t_L g9430 ( 
.A(n_8387),
.Y(n_9430)
);

OR2x6_ASAP7_75t_L g9431 ( 
.A(n_8830),
.B(n_7863),
.Y(n_9431)
);

OAI211xp5_ASAP7_75t_SL g9432 ( 
.A1(n_8521),
.A2(n_8304),
.B(n_8101),
.C(n_7541),
.Y(n_9432)
);

OAI21xp5_ASAP7_75t_L g9433 ( 
.A1(n_8585),
.A2(n_8286),
.B(n_6791),
.Y(n_9433)
);

INVx2_ASAP7_75t_L g9434 ( 
.A(n_8595),
.Y(n_9434)
);

INVx1_ASAP7_75t_L g9435 ( 
.A(n_8363),
.Y(n_9435)
);

AND2x2_ASAP7_75t_SL g9436 ( 
.A(n_8740),
.B(n_8178),
.Y(n_9436)
);

OAI22xp5_ASAP7_75t_L g9437 ( 
.A1(n_8635),
.A2(n_7753),
.B1(n_7860),
.B2(n_7588),
.Y(n_9437)
);

AOI22xp33_ASAP7_75t_L g9438 ( 
.A1(n_8740),
.A2(n_7834),
.B1(n_7847),
.B2(n_7818),
.Y(n_9438)
);

INVx1_ASAP7_75t_L g9439 ( 
.A(n_8364),
.Y(n_9439)
);

AND2x2_ASAP7_75t_L g9440 ( 
.A(n_8856),
.B(n_8201),
.Y(n_9440)
);

INVx1_ASAP7_75t_L g9441 ( 
.A(n_8370),
.Y(n_9441)
);

AOI22xp33_ASAP7_75t_L g9442 ( 
.A1(n_9044),
.A2(n_9064),
.B1(n_9078),
.B2(n_9057),
.Y(n_9442)
);

AND2x2_ASAP7_75t_L g9443 ( 
.A(n_8856),
.B(n_8201),
.Y(n_9443)
);

OAI22xp5_ASAP7_75t_L g9444 ( 
.A1(n_9050),
.A2(n_7753),
.B1(n_7860),
.B2(n_7588),
.Y(n_9444)
);

AOI211xp5_ASAP7_75t_L g9445 ( 
.A1(n_8587),
.A2(n_8211),
.B(n_6623),
.C(n_8119),
.Y(n_9445)
);

INVx1_ASAP7_75t_L g9446 ( 
.A(n_8374),
.Y(n_9446)
);

NOR2xp33_ASAP7_75t_L g9447 ( 
.A(n_8802),
.B(n_7748),
.Y(n_9447)
);

BUFx4f_ASAP7_75t_SL g9448 ( 
.A(n_8455),
.Y(n_9448)
);

AOI22xp33_ASAP7_75t_L g9449 ( 
.A1(n_9044),
.A2(n_7847),
.B1(n_7848),
.B2(n_7818),
.Y(n_9449)
);

AND2x2_ASAP7_75t_L g9450 ( 
.A(n_8817),
.B(n_8201),
.Y(n_9450)
);

AND2x2_ASAP7_75t_L g9451 ( 
.A(n_8817),
.B(n_8201),
.Y(n_9451)
);

HB1xp67_ASAP7_75t_L g9452 ( 
.A(n_8560),
.Y(n_9452)
);

OR2x2_ASAP7_75t_L g9453 ( 
.A(n_8626),
.B(n_8115),
.Y(n_9453)
);

INVx1_ASAP7_75t_L g9454 ( 
.A(n_8380),
.Y(n_9454)
);

AOI22xp33_ASAP7_75t_L g9455 ( 
.A1(n_9057),
.A2(n_7848),
.B1(n_7856),
.B2(n_7847),
.Y(n_9455)
);

AOI22xp33_ASAP7_75t_L g9456 ( 
.A1(n_9064),
.A2(n_7856),
.B1(n_7848),
.B2(n_6813),
.Y(n_9456)
);

AOI22xp33_ASAP7_75t_L g9457 ( 
.A1(n_9078),
.A2(n_7856),
.B1(n_6813),
.B2(n_6794),
.Y(n_9457)
);

OAI22xp5_ASAP7_75t_L g9458 ( 
.A1(n_9050),
.A2(n_7908),
.B1(n_7988),
.B2(n_7931),
.Y(n_9458)
);

A2O1A1Ixp33_ASAP7_75t_L g9459 ( 
.A1(n_8587),
.A2(n_7053),
.B(n_6688),
.C(n_6791),
.Y(n_9459)
);

AOI21xp5_ASAP7_75t_L g9460 ( 
.A1(n_9156),
.A2(n_7162),
.B(n_8178),
.Y(n_9460)
);

OAI22xp5_ASAP7_75t_L g9461 ( 
.A1(n_9050),
.A2(n_7908),
.B1(n_7988),
.B2(n_7931),
.Y(n_9461)
);

OAI221xp5_ASAP7_75t_L g9462 ( 
.A1(n_8794),
.A2(n_7807),
.B1(n_7757),
.B2(n_6740),
.C(n_6813),
.Y(n_9462)
);

INVx1_ASAP7_75t_L g9463 ( 
.A(n_8382),
.Y(n_9463)
);

AOI22xp33_ASAP7_75t_L g9464 ( 
.A1(n_9087),
.A2(n_6813),
.B1(n_6794),
.B2(n_7475),
.Y(n_9464)
);

AOI22xp5_ASAP7_75t_L g9465 ( 
.A1(n_8916),
.A2(n_7049),
.B1(n_6978),
.B2(n_6794),
.Y(n_9465)
);

INVx1_ASAP7_75t_L g9466 ( 
.A(n_8388),
.Y(n_9466)
);

INVx2_ASAP7_75t_L g9467 ( 
.A(n_8619),
.Y(n_9467)
);

AOI22xp33_ASAP7_75t_L g9468 ( 
.A1(n_9087),
.A2(n_6794),
.B1(n_7578),
.B2(n_7475),
.Y(n_9468)
);

NAND2xp5_ASAP7_75t_L g9469 ( 
.A(n_8675),
.B(n_7585),
.Y(n_9469)
);

INVx3_ASAP7_75t_L g9470 ( 
.A(n_8836),
.Y(n_9470)
);

AOI22xp33_ASAP7_75t_SL g9471 ( 
.A1(n_8690),
.A2(n_6794),
.B1(n_6694),
.B2(n_6993),
.Y(n_9471)
);

NAND3xp33_ASAP7_75t_L g9472 ( 
.A(n_8675),
.B(n_7534),
.C(n_7529),
.Y(n_9472)
);

AOI22xp33_ASAP7_75t_L g9473 ( 
.A1(n_9094),
.A2(n_7578),
.B1(n_7596),
.B2(n_7475),
.Y(n_9473)
);

BUFx2_ASAP7_75t_L g9474 ( 
.A(n_8383),
.Y(n_9474)
);

AOI21xp5_ASAP7_75t_L g9475 ( 
.A1(n_8359),
.A2(n_8072),
.B(n_8070),
.Y(n_9475)
);

AOI22xp33_ASAP7_75t_SL g9476 ( 
.A1(n_8707),
.A2(n_6694),
.B1(n_6993),
.B2(n_8136),
.Y(n_9476)
);

AND2x4_ASAP7_75t_L g9477 ( 
.A(n_8699),
.B(n_8248),
.Y(n_9477)
);

AOI22xp33_ASAP7_75t_L g9478 ( 
.A1(n_9094),
.A2(n_7578),
.B1(n_7596),
.B2(n_7475),
.Y(n_9478)
);

OAI221xp5_ASAP7_75t_L g9479 ( 
.A1(n_8794),
.A2(n_6694),
.B1(n_8186),
.B2(n_7858),
.C(n_8109),
.Y(n_9479)
);

AOI22xp33_ASAP7_75t_L g9480 ( 
.A1(n_9098),
.A2(n_7596),
.B1(n_7606),
.B2(n_7578),
.Y(n_9480)
);

NAND2xp5_ASAP7_75t_L g9481 ( 
.A(n_8699),
.B(n_7585),
.Y(n_9481)
);

AOI21xp5_ASAP7_75t_L g9482 ( 
.A1(n_8359),
.A2(n_7075),
.B(n_7731),
.Y(n_9482)
);

INVx2_ASAP7_75t_L g9483 ( 
.A(n_8619),
.Y(n_9483)
);

INVx1_ASAP7_75t_L g9484 ( 
.A(n_8390),
.Y(n_9484)
);

AOI22xp33_ASAP7_75t_L g9485 ( 
.A1(n_9098),
.A2(n_7606),
.B1(n_7626),
.B2(n_7596),
.Y(n_9485)
);

AOI21xp5_ASAP7_75t_L g9486 ( 
.A1(n_8359),
.A2(n_7075),
.B(n_8343),
.Y(n_9486)
);

OAI211xp5_ASAP7_75t_L g9487 ( 
.A1(n_8602),
.A2(n_8209),
.B(n_8221),
.C(n_7838),
.Y(n_9487)
);

OAI21x1_ASAP7_75t_L g9488 ( 
.A1(n_8688),
.A2(n_8142),
.B(n_8129),
.Y(n_9488)
);

HB1xp67_ASAP7_75t_L g9489 ( 
.A(n_8572),
.Y(n_9489)
);

BUFx6f_ASAP7_75t_L g9490 ( 
.A(n_8397),
.Y(n_9490)
);

AOI22xp33_ASAP7_75t_L g9491 ( 
.A1(n_9109),
.A2(n_7626),
.B1(n_7627),
.B2(n_7606),
.Y(n_9491)
);

CKINVDCx20_ASAP7_75t_R g9492 ( 
.A(n_8848),
.Y(n_9492)
);

AOI21xp5_ASAP7_75t_SL g9493 ( 
.A1(n_8761),
.A2(n_7520),
.B(n_7235),
.Y(n_9493)
);

AOI21xp33_ASAP7_75t_L g9494 ( 
.A1(n_8625),
.A2(n_8209),
.B(n_7930),
.Y(n_9494)
);

OAI22xp5_ASAP7_75t_L g9495 ( 
.A1(n_9065),
.A2(n_7908),
.B1(n_7988),
.B2(n_7931),
.Y(n_9495)
);

OAI221xp5_ASAP7_75t_L g9496 ( 
.A1(n_8833),
.A2(n_6694),
.B1(n_8074),
.B2(n_7338),
.C(n_7036),
.Y(n_9496)
);

NAND2xp5_ASAP7_75t_L g9497 ( 
.A(n_8615),
.B(n_7616),
.Y(n_9497)
);

OAI21xp33_ASAP7_75t_L g9498 ( 
.A1(n_8833),
.A2(n_7036),
.B(n_7031),
.Y(n_9498)
);

AO21x2_ASAP7_75t_L g9499 ( 
.A1(n_9034),
.A2(n_7868),
.B(n_7867),
.Y(n_9499)
);

AOI22xp33_ASAP7_75t_L g9500 ( 
.A1(n_9109),
.A2(n_9117),
.B1(n_9113),
.B2(n_8832),
.Y(n_9500)
);

NAND2xp5_ASAP7_75t_L g9501 ( 
.A(n_8624),
.B(n_7789),
.Y(n_9501)
);

AOI22xp33_ASAP7_75t_L g9502 ( 
.A1(n_9113),
.A2(n_7626),
.B1(n_7627),
.B2(n_7606),
.Y(n_9502)
);

AOI22xp33_ASAP7_75t_SL g9503 ( 
.A1(n_8707),
.A2(n_6694),
.B1(n_6993),
.B2(n_6688),
.Y(n_9503)
);

OAI221xp5_ASAP7_75t_L g9504 ( 
.A1(n_8981),
.A2(n_7338),
.B1(n_7031),
.B2(n_8268),
.C(n_8246),
.Y(n_9504)
);

AOI22xp33_ASAP7_75t_L g9505 ( 
.A1(n_9117),
.A2(n_7627),
.B1(n_7633),
.B2(n_7626),
.Y(n_9505)
);

AOI221xp5_ASAP7_75t_L g9506 ( 
.A1(n_8401),
.A2(n_7125),
.B1(n_7869),
.B2(n_7868),
.C(n_7867),
.Y(n_9506)
);

BUFx3_ASAP7_75t_L g9507 ( 
.A(n_8848),
.Y(n_9507)
);

NAND2xp5_ASAP7_75t_L g9508 ( 
.A(n_8627),
.B(n_7789),
.Y(n_9508)
);

OAI22xp5_ASAP7_75t_L g9509 ( 
.A1(n_9065),
.A2(n_7908),
.B1(n_7988),
.B2(n_7931),
.Y(n_9509)
);

OR2x2_ASAP7_75t_L g9510 ( 
.A(n_8626),
.B(n_8115),
.Y(n_9510)
);

AOI22xp33_ASAP7_75t_L g9511 ( 
.A1(n_8829),
.A2(n_7633),
.B1(n_7709),
.B2(n_7627),
.Y(n_9511)
);

AOI221xp5_ASAP7_75t_L g9512 ( 
.A1(n_8401),
.A2(n_7869),
.B1(n_7912),
.B2(n_7897),
.C(n_7882),
.Y(n_9512)
);

AO31x2_ASAP7_75t_L g9513 ( 
.A1(n_9034),
.A2(n_7897),
.A3(n_7912),
.B(n_7882),
.Y(n_9513)
);

AOI22xp33_ASAP7_75t_L g9514 ( 
.A1(n_8829),
.A2(n_7709),
.B1(n_7761),
.B2(n_7633),
.Y(n_9514)
);

CKINVDCx11_ASAP7_75t_R g9515 ( 
.A(n_8970),
.Y(n_9515)
);

BUFx3_ASAP7_75t_L g9516 ( 
.A(n_8879),
.Y(n_9516)
);

AOI22xp33_ASAP7_75t_L g9517 ( 
.A1(n_8832),
.A2(n_7709),
.B1(n_7761),
.B2(n_7633),
.Y(n_9517)
);

BUFx2_ASAP7_75t_L g9518 ( 
.A(n_8796),
.Y(n_9518)
);

NOR2xp33_ASAP7_75t_L g9519 ( 
.A(n_8670),
.B(n_8347),
.Y(n_9519)
);

AND2x4_ASAP7_75t_L g9520 ( 
.A(n_8852),
.B(n_8248),
.Y(n_9520)
);

AND2x2_ASAP7_75t_L g9521 ( 
.A(n_8852),
.B(n_8673),
.Y(n_9521)
);

INVx1_ASAP7_75t_L g9522 ( 
.A(n_8394),
.Y(n_9522)
);

INVx4_ASAP7_75t_L g9523 ( 
.A(n_8397),
.Y(n_9523)
);

AOI221xp5_ASAP7_75t_L g9524 ( 
.A1(n_8408),
.A2(n_7097),
.B1(n_7964),
.B2(n_7005),
.C(n_7067),
.Y(n_9524)
);

INVx1_ASAP7_75t_L g9525 ( 
.A(n_8395),
.Y(n_9525)
);

OAI221xp5_ASAP7_75t_L g9526 ( 
.A1(n_8981),
.A2(n_9021),
.B1(n_9022),
.B2(n_8521),
.C(n_9059),
.Y(n_9526)
);

AOI222xp33_ASAP7_75t_L g9527 ( 
.A1(n_8521),
.A2(n_6580),
.B1(n_7067),
.B2(n_7076),
.C1(n_7005),
.C2(n_7097),
.Y(n_9527)
);

AOI22xp33_ASAP7_75t_L g9528 ( 
.A1(n_8839),
.A2(n_7761),
.B1(n_7770),
.B2(n_7709),
.Y(n_9528)
);

AND2x2_ASAP7_75t_L g9529 ( 
.A(n_8673),
.B(n_8248),
.Y(n_9529)
);

AOI22xp33_ASAP7_75t_L g9530 ( 
.A1(n_8839),
.A2(n_7770),
.B1(n_7784),
.B2(n_7761),
.Y(n_9530)
);

INVx1_ASAP7_75t_L g9531 ( 
.A(n_8396),
.Y(n_9531)
);

AOI22xp33_ASAP7_75t_L g9532 ( 
.A1(n_8853),
.A2(n_7784),
.B1(n_7835),
.B2(n_7770),
.Y(n_9532)
);

AOI21xp33_ASAP7_75t_L g9533 ( 
.A1(n_8625),
.A2(n_7930),
.B(n_7902),
.Y(n_9533)
);

OR2x2_ASAP7_75t_L g9534 ( 
.A(n_8677),
.B(n_8134),
.Y(n_9534)
);

INVx1_ASAP7_75t_L g9535 ( 
.A(n_8403),
.Y(n_9535)
);

AND2x2_ASAP7_75t_SL g9536 ( 
.A(n_8992),
.B(n_8248),
.Y(n_9536)
);

OAI22xp33_ASAP7_75t_L g9537 ( 
.A1(n_8521),
.A2(n_6815),
.B1(n_7398),
.B2(n_7189),
.Y(n_9537)
);

BUFx6f_ASAP7_75t_L g9538 ( 
.A(n_8407),
.Y(n_9538)
);

INVx4_ASAP7_75t_L g9539 ( 
.A(n_8407),
.Y(n_9539)
);

OAI21xp5_ASAP7_75t_L g9540 ( 
.A1(n_8480),
.A2(n_6634),
.B(n_8129),
.Y(n_9540)
);

AOI22xp33_ASAP7_75t_L g9541 ( 
.A1(n_8853),
.A2(n_8867),
.B1(n_8869),
.B2(n_8855),
.Y(n_9541)
);

AOI221xp5_ASAP7_75t_L g9542 ( 
.A1(n_8408),
.A2(n_7964),
.B1(n_6822),
.B2(n_7021),
.C(n_7079),
.Y(n_9542)
);

AND2x2_ASAP7_75t_L g9543 ( 
.A(n_8682),
.B(n_8255),
.Y(n_9543)
);

OAI22xp5_ASAP7_75t_L g9544 ( 
.A1(n_9065),
.A2(n_8068),
.B1(n_8031),
.B2(n_8221),
.Y(n_9544)
);

AOI22xp33_ASAP7_75t_L g9545 ( 
.A1(n_8855),
.A2(n_7784),
.B1(n_7835),
.B2(n_7770),
.Y(n_9545)
);

INVx2_ASAP7_75t_L g9546 ( 
.A(n_8629),
.Y(n_9546)
);

AOI22xp33_ASAP7_75t_L g9547 ( 
.A1(n_8867),
.A2(n_7835),
.B1(n_7839),
.B2(n_7784),
.Y(n_9547)
);

OAI221xp5_ASAP7_75t_L g9548 ( 
.A1(n_9021),
.A2(n_7338),
.B1(n_8268),
.B2(n_8246),
.C(n_7902),
.Y(n_9548)
);

NAND2x1_ASAP7_75t_L g9549 ( 
.A(n_8656),
.B(n_6684),
.Y(n_9549)
);

NAND2xp5_ASAP7_75t_SL g9550 ( 
.A(n_8836),
.B(n_7529),
.Y(n_9550)
);

INVx3_ASAP7_75t_SL g9551 ( 
.A(n_8730),
.Y(n_9551)
);

INVx4_ASAP7_75t_L g9552 ( 
.A(n_8734),
.Y(n_9552)
);

BUFx3_ASAP7_75t_L g9553 ( 
.A(n_8730),
.Y(n_9553)
);

AOI221xp5_ASAP7_75t_L g9554 ( 
.A1(n_8869),
.A2(n_7964),
.B1(n_6822),
.B2(n_7021),
.C(n_7079),
.Y(n_9554)
);

AND2x2_ASAP7_75t_L g9555 ( 
.A(n_8682),
.B(n_8255),
.Y(n_9555)
);

INVx1_ASAP7_75t_L g9556 ( 
.A(n_8404),
.Y(n_9556)
);

NAND2xp5_ASAP7_75t_L g9557 ( 
.A(n_8678),
.B(n_7845),
.Y(n_9557)
);

AND2x4_ASAP7_75t_L g9558 ( 
.A(n_8629),
.B(n_8255),
.Y(n_9558)
);

AND2x2_ASAP7_75t_L g9559 ( 
.A(n_9137),
.B(n_8255),
.Y(n_9559)
);

NAND3xp33_ASAP7_75t_L g9560 ( 
.A(n_8685),
.B(n_7534),
.C(n_7529),
.Y(n_9560)
);

AOI22xp33_ASAP7_75t_SL g9561 ( 
.A1(n_8431),
.A2(n_6993),
.B1(n_6688),
.B2(n_7062),
.Y(n_9561)
);

OAI22xp5_ASAP7_75t_L g9562 ( 
.A1(n_8431),
.A2(n_8068),
.B1(n_8031),
.B2(n_7289),
.Y(n_9562)
);

BUFx2_ASAP7_75t_L g9563 ( 
.A(n_8487),
.Y(n_9563)
);

OAI221xp5_ASAP7_75t_L g9564 ( 
.A1(n_9022),
.A2(n_7338),
.B1(n_8268),
.B2(n_8246),
.C(n_7902),
.Y(n_9564)
);

AOI22xp33_ASAP7_75t_SL g9565 ( 
.A1(n_8446),
.A2(n_6993),
.B1(n_7062),
.B2(n_8246),
.Y(n_9565)
);

OAI22xp5_ASAP7_75t_L g9566 ( 
.A1(n_8446),
.A2(n_8068),
.B1(n_8031),
.B2(n_7289),
.Y(n_9566)
);

OAI221xp5_ASAP7_75t_L g9567 ( 
.A1(n_9059),
.A2(n_7338),
.B1(n_8268),
.B2(n_7902),
.C(n_7989),
.Y(n_9567)
);

AOI22xp33_ASAP7_75t_L g9568 ( 
.A1(n_8873),
.A2(n_7839),
.B1(n_7861),
.B2(n_7835),
.Y(n_9568)
);

OAI22xp5_ASAP7_75t_L g9569 ( 
.A1(n_8460),
.A2(n_8031),
.B1(n_8068),
.B2(n_7076),
.Y(n_9569)
);

INVx1_ASAP7_75t_L g9570 ( 
.A(n_8405),
.Y(n_9570)
);

AO31x2_ASAP7_75t_L g9571 ( 
.A1(n_9041),
.A2(n_8029),
.A3(n_7974),
.B(n_8041),
.Y(n_9571)
);

INVx2_ASAP7_75t_L g9572 ( 
.A(n_8429),
.Y(n_9572)
);

NAND3xp33_ASAP7_75t_SL g9573 ( 
.A(n_8808),
.B(n_7884),
.C(n_7838),
.Y(n_9573)
);

OAI22xp5_ASAP7_75t_L g9574 ( 
.A1(n_8460),
.A2(n_7991),
.B1(n_7354),
.B2(n_6708),
.Y(n_9574)
);

OAI211xp5_ASAP7_75t_SL g9575 ( 
.A1(n_8372),
.A2(n_7662),
.B(n_7903),
.C(n_7845),
.Y(n_9575)
);

AOI21xp5_ASAP7_75t_L g9576 ( 
.A1(n_8480),
.A2(n_7010),
.B(n_7158),
.Y(n_9576)
);

AOI21xp5_ASAP7_75t_L g9577 ( 
.A1(n_8481),
.A2(n_7010),
.B(n_7158),
.Y(n_9577)
);

AOI22xp5_ASAP7_75t_L g9578 ( 
.A1(n_8723),
.A2(n_6978),
.B1(n_6993),
.B2(n_6623),
.Y(n_9578)
);

AOI22xp33_ASAP7_75t_L g9579 ( 
.A1(n_8873),
.A2(n_7861),
.B1(n_7865),
.B2(n_7839),
.Y(n_9579)
);

AOI22xp33_ASAP7_75t_L g9580 ( 
.A1(n_8876),
.A2(n_7861),
.B1(n_7865),
.B2(n_7839),
.Y(n_9580)
);

BUFx2_ASAP7_75t_L g9581 ( 
.A(n_8845),
.Y(n_9581)
);

AO31x2_ASAP7_75t_L g9582 ( 
.A1(n_9041),
.A2(n_8029),
.A3(n_7974),
.B(n_8019),
.Y(n_9582)
);

AOI22xp33_ASAP7_75t_L g9583 ( 
.A1(n_8876),
.A2(n_7865),
.B1(n_7905),
.B2(n_7861),
.Y(n_9583)
);

HB1xp67_ASAP7_75t_L g9584 ( 
.A(n_8701),
.Y(n_9584)
);

OAI221xp5_ASAP7_75t_L g9585 ( 
.A1(n_9059),
.A2(n_7989),
.B1(n_8000),
.B2(n_7930),
.C(n_7759),
.Y(n_9585)
);

AND2x2_ASAP7_75t_L g9586 ( 
.A(n_9137),
.B(n_7529),
.Y(n_9586)
);

AOI221xp5_ASAP7_75t_L g9587 ( 
.A1(n_8878),
.A2(n_7987),
.B1(n_8029),
.B2(n_7974),
.C(n_8039),
.Y(n_9587)
);

INVx3_ASAP7_75t_L g9588 ( 
.A(n_8836),
.Y(n_9588)
);

INVx1_ASAP7_75t_L g9589 ( 
.A(n_8406),
.Y(n_9589)
);

OAI21xp33_ASAP7_75t_L g9590 ( 
.A1(n_8772),
.A2(n_8156),
.B(n_8142),
.Y(n_9590)
);

AOI221xp5_ASAP7_75t_L g9591 ( 
.A1(n_8878),
.A2(n_8039),
.B1(n_8043),
.B2(n_8042),
.C(n_8040),
.Y(n_9591)
);

AOI22xp33_ASAP7_75t_L g9592 ( 
.A1(n_8880),
.A2(n_7905),
.B1(n_7955),
.B2(n_7865),
.Y(n_9592)
);

OAI21xp5_ASAP7_75t_L g9593 ( 
.A1(n_8481),
.A2(n_8479),
.B(n_8439),
.Y(n_9593)
);

OAI221xp5_ASAP7_75t_L g9594 ( 
.A1(n_9059),
.A2(n_8858),
.B1(n_8889),
.B2(n_8411),
.C(n_8656),
.Y(n_9594)
);

NAND2xp5_ASAP7_75t_L g9595 ( 
.A(n_8708),
.B(n_7903),
.Y(n_9595)
);

INVx2_ASAP7_75t_SL g9596 ( 
.A(n_8670),
.Y(n_9596)
);

AOI222xp33_ASAP7_75t_L g9597 ( 
.A1(n_8638),
.A2(n_6580),
.B1(n_8042),
.B2(n_8043),
.C1(n_8040),
.C2(n_8039),
.Y(n_9597)
);

INVxp33_ASAP7_75t_L g9598 ( 
.A(n_8764),
.Y(n_9598)
);

AOI22xp33_ASAP7_75t_L g9599 ( 
.A1(n_8880),
.A2(n_7955),
.B1(n_7905),
.B2(n_7534),
.Y(n_9599)
);

OAI22xp33_ASAP7_75t_L g9600 ( 
.A1(n_8411),
.A2(n_7166),
.B1(n_7189),
.B2(n_7759),
.Y(n_9600)
);

OAI22xp5_ASAP7_75t_L g9601 ( 
.A1(n_8638),
.A2(n_6708),
.B1(n_6917),
.B2(n_7310),
.Y(n_9601)
);

INVx5_ASAP7_75t_L g9602 ( 
.A(n_8734),
.Y(n_9602)
);

AOI22xp33_ASAP7_75t_SL g9603 ( 
.A1(n_8663),
.A2(n_9038),
.B1(n_8777),
.B2(n_8800),
.Y(n_9603)
);

OAI21xp33_ASAP7_75t_L g9604 ( 
.A1(n_8663),
.A2(n_7351),
.B(n_7920),
.Y(n_9604)
);

INVx3_ASAP7_75t_L g9605 ( 
.A(n_8895),
.Y(n_9605)
);

OR2x6_ASAP7_75t_L g9606 ( 
.A(n_8830),
.B(n_7899),
.Y(n_9606)
);

NAND2x1_ASAP7_75t_L g9607 ( 
.A(n_8656),
.B(n_8247),
.Y(n_9607)
);

OR2x6_ASAP7_75t_L g9608 ( 
.A(n_8734),
.B(n_7899),
.Y(n_9608)
);

AOI22xp33_ASAP7_75t_L g9609 ( 
.A1(n_8885),
.A2(n_7955),
.B1(n_7905),
.B2(n_7534),
.Y(n_9609)
);

INVx1_ASAP7_75t_L g9610 ( 
.A(n_8409),
.Y(n_9610)
);

AOI221xp5_ASAP7_75t_SL g9611 ( 
.A1(n_8429),
.A2(n_7221),
.B1(n_7884),
.B2(n_8140),
.C(n_8094),
.Y(n_9611)
);

AOI21xp33_ASAP7_75t_SL g9612 ( 
.A1(n_8553),
.A2(n_7878),
.B(n_7795),
.Y(n_9612)
);

OAI221xp5_ASAP7_75t_L g9613 ( 
.A1(n_8858),
.A2(n_7989),
.B1(n_8000),
.B2(n_7930),
.C(n_7759),
.Y(n_9613)
);

AOI22xp33_ASAP7_75t_SL g9614 ( 
.A1(n_9038),
.A2(n_8777),
.B1(n_8800),
.B2(n_8746),
.Y(n_9614)
);

INVx1_ASAP7_75t_L g9615 ( 
.A(n_8412),
.Y(n_9615)
);

INVx2_ASAP7_75t_SL g9616 ( 
.A(n_8676),
.Y(n_9616)
);

A2O1A1Ixp33_ASAP7_75t_L g9617 ( 
.A1(n_8439),
.A2(n_7039),
.B(n_7030),
.C(n_7955),
.Y(n_9617)
);

OR2x2_ASAP7_75t_L g9618 ( 
.A(n_8677),
.B(n_8134),
.Y(n_9618)
);

AOI22xp33_ASAP7_75t_L g9619 ( 
.A1(n_8885),
.A2(n_7534),
.B1(n_7685),
.B2(n_7529),
.Y(n_9619)
);

AO21x2_ASAP7_75t_L g9620 ( 
.A1(n_8365),
.A2(n_8019),
.B(n_8009),
.Y(n_9620)
);

AND2x2_ASAP7_75t_L g9621 ( 
.A(n_9148),
.B(n_7529),
.Y(n_9621)
);

HB1xp67_ASAP7_75t_L g9622 ( 
.A(n_8714),
.Y(n_9622)
);

AOI211xp5_ASAP7_75t_L g9623 ( 
.A1(n_8479),
.A2(n_6647),
.B(n_6652),
.C(n_6577),
.Y(n_9623)
);

NAND2xp5_ASAP7_75t_L g9624 ( 
.A(n_8724),
.B(n_7920),
.Y(n_9624)
);

AOI22xp33_ASAP7_75t_L g9625 ( 
.A1(n_8886),
.A2(n_7685),
.B1(n_7762),
.B2(n_7534),
.Y(n_9625)
);

INVx2_ASAP7_75t_L g9626 ( 
.A(n_8429),
.Y(n_9626)
);

CKINVDCx5p33_ASAP7_75t_R g9627 ( 
.A(n_9103),
.Y(n_9627)
);

AND2x2_ASAP7_75t_L g9628 ( 
.A(n_9148),
.B(n_7685),
.Y(n_9628)
);

INVx2_ASAP7_75t_L g9629 ( 
.A(n_8429),
.Y(n_9629)
);

AOI22xp33_ASAP7_75t_L g9630 ( 
.A1(n_8886),
.A2(n_7762),
.B1(n_7785),
.B2(n_7685),
.Y(n_9630)
);

OR2x2_ASAP7_75t_L g9631 ( 
.A(n_8684),
.B(n_7072),
.Y(n_9631)
);

OAI221xp5_ASAP7_75t_L g9632 ( 
.A1(n_8889),
.A2(n_8000),
.B1(n_7989),
.B2(n_8096),
.C(n_7039),
.Y(n_9632)
);

CKINVDCx5p33_ASAP7_75t_R g9633 ( 
.A(n_9103),
.Y(n_9633)
);

BUFx3_ASAP7_75t_L g9634 ( 
.A(n_8676),
.Y(n_9634)
);

OAI22xp5_ASAP7_75t_L g9635 ( 
.A1(n_8496),
.A2(n_6917),
.B1(n_7310),
.B2(n_6955),
.Y(n_9635)
);

OAI22xp33_ASAP7_75t_L g9636 ( 
.A1(n_8411),
.A2(n_7189),
.B1(n_7166),
.B2(n_7410),
.Y(n_9636)
);

AOI22xp33_ASAP7_75t_L g9637 ( 
.A1(n_8897),
.A2(n_7762),
.B1(n_7785),
.B2(n_7685),
.Y(n_9637)
);

HB1xp67_ASAP7_75t_L g9638 ( 
.A(n_8736),
.Y(n_9638)
);

OR2x2_ASAP7_75t_L g9639 ( 
.A(n_8684),
.B(n_7072),
.Y(n_9639)
);

OAI22xp33_ASAP7_75t_L g9640 ( 
.A1(n_8411),
.A2(n_7166),
.B1(n_7410),
.B2(n_7213),
.Y(n_9640)
);

AND2x2_ASAP7_75t_L g9641 ( 
.A(n_8969),
.B(n_7685),
.Y(n_9641)
);

INVx1_ASAP7_75t_L g9642 ( 
.A(n_8415),
.Y(n_9642)
);

INVx1_ASAP7_75t_L g9643 ( 
.A(n_8418),
.Y(n_9643)
);

OAI21xp33_ASAP7_75t_SL g9644 ( 
.A1(n_8356),
.A2(n_9152),
.B(n_9145),
.Y(n_9644)
);

AOI221xp5_ASAP7_75t_L g9645 ( 
.A1(n_8897),
.A2(n_8042),
.B1(n_8050),
.B2(n_8043),
.C(n_8040),
.Y(n_9645)
);

NAND2xp5_ASAP7_75t_L g9646 ( 
.A(n_8752),
.B(n_7993),
.Y(n_9646)
);

AOI222xp33_ASAP7_75t_SL g9647 ( 
.A1(n_8640),
.A2(n_8094),
.B1(n_8181),
.B2(n_8140),
.C1(n_8205),
.C2(n_8200),
.Y(n_9647)
);

AO21x2_ASAP7_75t_L g9648 ( 
.A1(n_8365),
.A2(n_8009),
.B(n_8050),
.Y(n_9648)
);

NOR2xp33_ASAP7_75t_L g9649 ( 
.A(n_8758),
.B(n_8199),
.Y(n_9649)
);

INVx1_ASAP7_75t_L g9650 ( 
.A(n_8424),
.Y(n_9650)
);

HB1xp67_ASAP7_75t_L g9651 ( 
.A(n_8785),
.Y(n_9651)
);

AOI22xp33_ASAP7_75t_L g9652 ( 
.A1(n_8898),
.A2(n_7785),
.B1(n_7762),
.B2(n_6993),
.Y(n_9652)
);

AND2x2_ASAP7_75t_L g9653 ( 
.A(n_8969),
.B(n_7762),
.Y(n_9653)
);

OAI22xp5_ASAP7_75t_SL g9654 ( 
.A1(n_8591),
.A2(n_6280),
.B1(n_6284),
.B2(n_6275),
.Y(n_9654)
);

AND2x2_ASAP7_75t_L g9655 ( 
.A(n_8989),
.B(n_7762),
.Y(n_9655)
);

INVx2_ASAP7_75t_L g9656 ( 
.A(n_8429),
.Y(n_9656)
);

AOI22xp33_ASAP7_75t_L g9657 ( 
.A1(n_8898),
.A2(n_7785),
.B1(n_6993),
.B2(n_6866),
.Y(n_9657)
);

BUFx12f_ASAP7_75t_L g9658 ( 
.A(n_9116),
.Y(n_9658)
);

AOI22xp33_ASAP7_75t_L g9659 ( 
.A1(n_8909),
.A2(n_7785),
.B1(n_6993),
.B2(n_6866),
.Y(n_9659)
);

AOI221xp5_ASAP7_75t_L g9660 ( 
.A1(n_8909),
.A2(n_8108),
.B1(n_8122),
.B2(n_8106),
.C(n_8050),
.Y(n_9660)
);

AOI221xp5_ASAP7_75t_L g9661 ( 
.A1(n_8913),
.A2(n_8122),
.B1(n_8127),
.B2(n_8108),
.C(n_8106),
.Y(n_9661)
);

AOI22xp5_ASAP7_75t_L g9662 ( 
.A1(n_9086),
.A2(n_6993),
.B1(n_7213),
.B2(n_7161),
.Y(n_9662)
);

AOI22xp33_ASAP7_75t_L g9663 ( 
.A1(n_8913),
.A2(n_7785),
.B1(n_6468),
.B2(n_6491),
.Y(n_9663)
);

NAND2xp5_ASAP7_75t_L g9664 ( 
.A(n_8791),
.B(n_7993),
.Y(n_9664)
);

AND2x2_ASAP7_75t_L g9665 ( 
.A(n_8989),
.B(n_8149),
.Y(n_9665)
);

OAI22xp5_ASAP7_75t_L g9666 ( 
.A1(n_8496),
.A2(n_7310),
.B1(n_6955),
.B2(n_6760),
.Y(n_9666)
);

AOI221xp5_ASAP7_75t_L g9667 ( 
.A1(n_8915),
.A2(n_8108),
.B1(n_8127),
.B2(n_8122),
.C(n_8106),
.Y(n_9667)
);

CKINVDCx5p33_ASAP7_75t_R g9668 ( 
.A(n_9116),
.Y(n_9668)
);

OAI211xp5_ASAP7_75t_L g9669 ( 
.A1(n_8772),
.A2(n_8181),
.B(n_8000),
.C(n_6652),
.Y(n_9669)
);

AOI221xp5_ASAP7_75t_L g9670 ( 
.A1(n_8915),
.A2(n_8131),
.B1(n_8137),
.B2(n_8132),
.C(n_8127),
.Y(n_9670)
);

AOI222xp33_ASAP7_75t_L g9671 ( 
.A1(n_8917),
.A2(n_8131),
.B1(n_8137),
.B2(n_8160),
.C1(n_8146),
.C2(n_8132),
.Y(n_9671)
);

INVx1_ASAP7_75t_L g9672 ( 
.A(n_8433),
.Y(n_9672)
);

AOI22xp33_ASAP7_75t_L g9673 ( 
.A1(n_8917),
.A2(n_6468),
.B1(n_6491),
.B2(n_6458),
.Y(n_9673)
);

OAI22xp5_ASAP7_75t_L g9674 ( 
.A1(n_8510),
.A2(n_8623),
.B1(n_8713),
.B2(n_8686),
.Y(n_9674)
);

AOI21xp5_ASAP7_75t_L g9675 ( 
.A1(n_8505),
.A2(n_8302),
.B(n_8001),
.Y(n_9675)
);

AOI22xp33_ASAP7_75t_L g9676 ( 
.A1(n_8920),
.A2(n_6468),
.B1(n_6491),
.B2(n_6458),
.Y(n_9676)
);

AOI221xp5_ASAP7_75t_L g9677 ( 
.A1(n_8920),
.A2(n_8132),
.B1(n_8146),
.B2(n_8137),
.C(n_8131),
.Y(n_9677)
);

AOI221xp5_ASAP7_75t_L g9678 ( 
.A1(n_8924),
.A2(n_8160),
.B1(n_8203),
.B2(n_8197),
.C(n_8146),
.Y(n_9678)
);

AOI22xp33_ASAP7_75t_L g9679 ( 
.A1(n_8924),
.A2(n_6468),
.B1(n_6491),
.B2(n_6458),
.Y(n_9679)
);

OR2x2_ASAP7_75t_L g9680 ( 
.A(n_8686),
.B(n_7072),
.Y(n_9680)
);

AOI21xp5_ASAP7_75t_L g9681 ( 
.A1(n_8505),
.A2(n_8302),
.B(n_8001),
.Y(n_9681)
);

OAI22xp5_ASAP7_75t_L g9682 ( 
.A1(n_8510),
.A2(n_6760),
.B1(n_8247),
.B2(n_8096),
.Y(n_9682)
);

AOI22xp33_ASAP7_75t_SL g9683 ( 
.A1(n_8746),
.A2(n_6820),
.B1(n_6458),
.B2(n_6491),
.Y(n_9683)
);

NAND2x1_ASAP7_75t_L g9684 ( 
.A(n_8447),
.B(n_8247),
.Y(n_9684)
);

O2A1O1Ixp33_ASAP7_75t_L g9685 ( 
.A1(n_8793),
.A2(n_8260),
.B(n_8280),
.C(n_8229),
.Y(n_9685)
);

INVx3_ASAP7_75t_L g9686 ( 
.A(n_8895),
.Y(n_9686)
);

A2O1A1Ixp33_ASAP7_75t_L g9687 ( 
.A1(n_9106),
.A2(n_7030),
.B(n_6807),
.C(n_6972),
.Y(n_9687)
);

HB1xp67_ASAP7_75t_L g9688 ( 
.A(n_8900),
.Y(n_9688)
);

AND2x4_ASAP7_75t_SL g9689 ( 
.A(n_8571),
.B(n_6352),
.Y(n_9689)
);

NAND2x1p5_ASAP7_75t_L g9690 ( 
.A(n_8895),
.B(n_7113),
.Y(n_9690)
);

AOI221xp5_ASAP7_75t_L g9691 ( 
.A1(n_8925),
.A2(n_8160),
.B1(n_8207),
.B2(n_8203),
.C(n_8197),
.Y(n_9691)
);

OAI22xp5_ASAP7_75t_L g9692 ( 
.A1(n_8623),
.A2(n_8247),
.B1(n_8096),
.B2(n_7161),
.Y(n_9692)
);

AOI22xp33_ASAP7_75t_L g9693 ( 
.A1(n_8925),
.A2(n_6468),
.B1(n_6491),
.B2(n_6458),
.Y(n_9693)
);

AOI21xp33_ASAP7_75t_L g9694 ( 
.A1(n_8393),
.A2(n_8462),
.B(n_8443),
.Y(n_9694)
);

AOI22xp33_ASAP7_75t_L g9695 ( 
.A1(n_8927),
.A2(n_6468),
.B1(n_6885),
.B2(n_6458),
.Y(n_9695)
);

AOI22xp5_ASAP7_75t_L g9696 ( 
.A1(n_8801),
.A2(n_7222),
.B1(n_8296),
.B2(n_8243),
.Y(n_9696)
);

INVx1_ASAP7_75t_L g9697 ( 
.A(n_8434),
.Y(n_9697)
);

AOI22xp33_ASAP7_75t_L g9698 ( 
.A1(n_8927),
.A2(n_6913),
.B1(n_6885),
.B2(n_7520),
.Y(n_9698)
);

OAI21xp33_ASAP7_75t_L g9699 ( 
.A1(n_8738),
.A2(n_7351),
.B(n_8340),
.Y(n_9699)
);

INVx2_ASAP7_75t_L g9700 ( 
.A(n_8492),
.Y(n_9700)
);

INVx2_ASAP7_75t_L g9701 ( 
.A(n_8492),
.Y(n_9701)
);

AOI22xp33_ASAP7_75t_L g9702 ( 
.A1(n_8929),
.A2(n_6913),
.B1(n_6885),
.B2(n_7520),
.Y(n_9702)
);

AOI22xp33_ASAP7_75t_L g9703 ( 
.A1(n_8929),
.A2(n_6913),
.B1(n_6885),
.B2(n_7520),
.Y(n_9703)
);

AOI221xp5_ASAP7_75t_L g9704 ( 
.A1(n_8934),
.A2(n_8197),
.B1(n_8208),
.B2(n_8207),
.C(n_8203),
.Y(n_9704)
);

OR2x2_ASAP7_75t_L g9705 ( 
.A(n_8713),
.B(n_7041),
.Y(n_9705)
);

OAI22xp5_ASAP7_75t_L g9706 ( 
.A1(n_8738),
.A2(n_8096),
.B1(n_8354),
.B2(n_7698),
.Y(n_9706)
);

OR2x6_ASAP7_75t_L g9707 ( 
.A(n_8734),
.B(n_8022),
.Y(n_9707)
);

INVx1_ASAP7_75t_L g9708 ( 
.A(n_8436),
.Y(n_9708)
);

INVx4_ASAP7_75t_L g9709 ( 
.A(n_8837),
.Y(n_9709)
);

AOI22xp33_ASAP7_75t_L g9710 ( 
.A1(n_8934),
.A2(n_6913),
.B1(n_6885),
.B2(n_6807),
.Y(n_9710)
);

AOI22xp33_ASAP7_75t_L g9711 ( 
.A1(n_8938),
.A2(n_8941),
.B1(n_8951),
.B2(n_8940),
.Y(n_9711)
);

AOI22xp33_ASAP7_75t_L g9712 ( 
.A1(n_8938),
.A2(n_6913),
.B1(n_6885),
.B2(n_6807),
.Y(n_9712)
);

AOI221xp5_ASAP7_75t_L g9713 ( 
.A1(n_8940),
.A2(n_8207),
.B1(n_8269),
.B2(n_8251),
.C(n_8208),
.Y(n_9713)
);

INVx1_ASAP7_75t_L g9714 ( 
.A(n_8437),
.Y(n_9714)
);

INVx2_ASAP7_75t_L g9715 ( 
.A(n_8492),
.Y(n_9715)
);

AOI22xp33_ASAP7_75t_SL g9716 ( 
.A1(n_8813),
.A2(n_6820),
.B1(n_6913),
.B2(n_7222),
.Y(n_9716)
);

INVx2_ASAP7_75t_L g9717 ( 
.A(n_8492),
.Y(n_9717)
);

NAND2xp5_ASAP7_75t_L g9718 ( 
.A(n_8919),
.B(n_8340),
.Y(n_9718)
);

AOI221xp5_ASAP7_75t_L g9719 ( 
.A1(n_8941),
.A2(n_8269),
.B1(n_8285),
.B2(n_8251),
.C(n_8208),
.Y(n_9719)
);

AOI22xp33_ASAP7_75t_L g9720 ( 
.A1(n_8951),
.A2(n_7950),
.B1(n_7963),
.B2(n_7894),
.Y(n_9720)
);

CKINVDCx5p33_ASAP7_75t_R g9721 ( 
.A(n_8758),
.Y(n_9721)
);

AOI22xp5_ASAP7_75t_L g9722 ( 
.A1(n_8801),
.A2(n_6280),
.B1(n_6284),
.B2(n_6275),
.Y(n_9722)
);

OR2x2_ASAP7_75t_L g9723 ( 
.A(n_8994),
.B(n_7041),
.Y(n_9723)
);

OAI22xp33_ASAP7_75t_L g9724 ( 
.A1(n_8744),
.A2(n_6960),
.B1(n_7407),
.B2(n_7041),
.Y(n_9724)
);

AOI222xp33_ASAP7_75t_L g9725 ( 
.A1(n_8953),
.A2(n_8718),
.B1(n_8706),
.B2(n_8719),
.C1(n_8716),
.C2(n_8705),
.Y(n_9725)
);

AOI22xp33_ASAP7_75t_L g9726 ( 
.A1(n_8953),
.A2(n_7950),
.B1(n_7963),
.B2(n_7894),
.Y(n_9726)
);

AOI33xp33_ASAP7_75t_L g9727 ( 
.A1(n_8771),
.A2(n_6964),
.A3(n_6953),
.B1(n_6976),
.B2(n_6957),
.B3(n_8342),
.Y(n_9727)
);

INVx1_ASAP7_75t_L g9728 ( 
.A(n_8438),
.Y(n_9728)
);

INVx2_ASAP7_75t_SL g9729 ( 
.A(n_8567),
.Y(n_9729)
);

INVx2_ASAP7_75t_L g9730 ( 
.A(n_8492),
.Y(n_9730)
);

OAI221xp5_ASAP7_75t_L g9731 ( 
.A1(n_8447),
.A2(n_8563),
.B1(n_8662),
.B2(n_8620),
.C(n_8862),
.Y(n_9731)
);

INVx1_ASAP7_75t_L g9732 ( 
.A(n_8440),
.Y(n_9732)
);

OAI222xp33_ASAP7_75t_L g9733 ( 
.A1(n_8744),
.A2(n_8171),
.B1(n_8176),
.B2(n_8156),
.C1(n_6797),
.C2(n_6625),
.Y(n_9733)
);

HB1xp67_ASAP7_75t_L g9734 ( 
.A(n_8948),
.Y(n_9734)
);

AND2x4_ASAP7_75t_L g9735 ( 
.A(n_8921),
.B(n_7113),
.Y(n_9735)
);

OA21x2_ASAP7_75t_L g9736 ( 
.A1(n_8379),
.A2(n_8918),
.B(n_8781),
.Y(n_9736)
);

OAI21xp5_ASAP7_75t_L g9737 ( 
.A1(n_8781),
.A2(n_6634),
.B(n_8171),
.Y(n_9737)
);

AOI21xp33_ASAP7_75t_L g9738 ( 
.A1(n_8393),
.A2(n_8462),
.B(n_8443),
.Y(n_9738)
);

AOI22xp33_ASAP7_75t_SL g9739 ( 
.A1(n_8813),
.A2(n_6577),
.B1(n_6562),
.B2(n_6936),
.Y(n_9739)
);

HB1xp67_ASAP7_75t_L g9740 ( 
.A(n_8979),
.Y(n_9740)
);

INVx11_ASAP7_75t_L g9741 ( 
.A(n_8845),
.Y(n_9741)
);

BUFx12f_ASAP7_75t_L g9742 ( 
.A(n_8566),
.Y(n_9742)
);

OAI211xp5_ASAP7_75t_L g9743 ( 
.A1(n_8640),
.A2(n_8176),
.B(n_7110),
.C(n_7221),
.Y(n_9743)
);

AOI221xp5_ASAP7_75t_L g9744 ( 
.A1(n_8373),
.A2(n_8251),
.B1(n_8325),
.B2(n_8285),
.C(n_8269),
.Y(n_9744)
);

AOI22xp5_ASAP7_75t_L g9745 ( 
.A1(n_8801),
.A2(n_6280),
.B1(n_6284),
.B2(n_6275),
.Y(n_9745)
);

OAI221xp5_ASAP7_75t_SL g9746 ( 
.A1(n_8862),
.A2(n_6972),
.B1(n_7407),
.B2(n_7240),
.C(n_6960),
.Y(n_9746)
);

OAI22xp33_ASAP7_75t_L g9747 ( 
.A1(n_8447),
.A2(n_7269),
.B1(n_7216),
.B2(n_7223),
.Y(n_9747)
);

AOI221xp5_ASAP7_75t_L g9748 ( 
.A1(n_8373),
.A2(n_8285),
.B1(n_8325),
.B2(n_7344),
.C(n_7409),
.Y(n_9748)
);

NAND3xp33_ASAP7_75t_L g9749 ( 
.A(n_8997),
.B(n_7950),
.C(n_7894),
.Y(n_9749)
);

AOI22xp33_ASAP7_75t_L g9750 ( 
.A1(n_8705),
.A2(n_7950),
.B1(n_7963),
.B2(n_7894),
.Y(n_9750)
);

INVx2_ASAP7_75t_L g9751 ( 
.A(n_8566),
.Y(n_9751)
);

INVx3_ASAP7_75t_L g9752 ( 
.A(n_8911),
.Y(n_9752)
);

AOI222xp33_ASAP7_75t_L g9753 ( 
.A1(n_8706),
.A2(n_8325),
.B1(n_7214),
.B2(n_6953),
.C1(n_6964),
.C2(n_6976),
.Y(n_9753)
);

NAND2xp33_ASAP7_75t_R g9754 ( 
.A(n_8447),
.B(n_6098),
.Y(n_9754)
);

OAI21xp5_ASAP7_75t_L g9755 ( 
.A1(n_8551),
.A2(n_6634),
.B(n_6577),
.Y(n_9755)
);

NAND2xp5_ASAP7_75t_L g9756 ( 
.A(n_9003),
.B(n_6806),
.Y(n_9756)
);

AOI21xp5_ASAP7_75t_L g9757 ( 
.A1(n_9039),
.A2(n_8130),
.B(n_6861),
.Y(n_9757)
);

NAND2xp5_ASAP7_75t_L g9758 ( 
.A(n_9035),
.B(n_6806),
.Y(n_9758)
);

AOI33xp33_ASAP7_75t_L g9759 ( 
.A1(n_8771),
.A2(n_6964),
.A3(n_6953),
.B1(n_6976),
.B2(n_6957),
.B3(n_8342),
.Y(n_9759)
);

OAI22xp5_ASAP7_75t_L g9760 ( 
.A1(n_8563),
.A2(n_8890),
.B1(n_8958),
.B2(n_8944),
.Y(n_9760)
);

AOI222xp33_ASAP7_75t_L g9761 ( 
.A1(n_8716),
.A2(n_7214),
.B1(n_6957),
.B2(n_6564),
.C1(n_6861),
.C2(n_7372),
.Y(n_9761)
);

OAI221xp5_ASAP7_75t_L g9762 ( 
.A1(n_8563),
.A2(n_7192),
.B1(n_7197),
.B2(n_6988),
.C(n_7020),
.Y(n_9762)
);

AND2x2_ASAP7_75t_L g9763 ( 
.A(n_8990),
.B(n_8149),
.Y(n_9763)
);

INVx2_ASAP7_75t_L g9764 ( 
.A(n_8566),
.Y(n_9764)
);

AOI22xp33_ASAP7_75t_L g9765 ( 
.A1(n_8718),
.A2(n_8728),
.B1(n_8745),
.B2(n_8719),
.Y(n_9765)
);

OAI22xp33_ASAP7_75t_L g9766 ( 
.A1(n_8563),
.A2(n_7269),
.B1(n_7216),
.B2(n_7223),
.Y(n_9766)
);

AOI22xp33_ASAP7_75t_L g9767 ( 
.A1(n_8728),
.A2(n_7950),
.B1(n_7963),
.B2(n_7894),
.Y(n_9767)
);

HB1xp67_ASAP7_75t_L g9768 ( 
.A(n_9054),
.Y(n_9768)
);

AOI22xp33_ASAP7_75t_L g9769 ( 
.A1(n_8745),
.A2(n_7950),
.B1(n_7963),
.B2(n_7894),
.Y(n_9769)
);

NAND3xp33_ASAP7_75t_SL g9770 ( 
.A(n_8930),
.B(n_8795),
.C(n_8558),
.Y(n_9770)
);

AO31x2_ASAP7_75t_L g9771 ( 
.A1(n_8375),
.A2(n_8346),
.A3(n_8350),
.B(n_8345),
.Y(n_9771)
);

AOI221xp5_ASAP7_75t_L g9772 ( 
.A1(n_8375),
.A2(n_7344),
.B1(n_7409),
.B2(n_8346),
.C(n_8345),
.Y(n_9772)
);

OR2x6_ASAP7_75t_L g9773 ( 
.A(n_8837),
.B(n_8022),
.Y(n_9773)
);

OAI22xp33_ASAP7_75t_L g9774 ( 
.A1(n_9002),
.A2(n_7223),
.B1(n_6617),
.B2(n_6773),
.Y(n_9774)
);

AOI22xp33_ASAP7_75t_L g9775 ( 
.A1(n_8748),
.A2(n_8012),
.B1(n_8089),
.B2(n_7963),
.Y(n_9775)
);

HB1xp67_ASAP7_75t_L g9776 ( 
.A(n_9068),
.Y(n_9776)
);

AOI22xp33_ASAP7_75t_L g9777 ( 
.A1(n_8748),
.A2(n_8750),
.B1(n_8751),
.B2(n_8749),
.Y(n_9777)
);

OAI221xp5_ASAP7_75t_L g9778 ( 
.A1(n_8620),
.A2(n_7192),
.B1(n_7197),
.B2(n_6988),
.C(n_7020),
.Y(n_9778)
);

OAI22xp5_ASAP7_75t_L g9779 ( 
.A1(n_8890),
.A2(n_8354),
.B1(n_7959),
.B2(n_7960),
.Y(n_9779)
);

OA21x2_ASAP7_75t_L g9780 ( 
.A1(n_8379),
.A2(n_8315),
.B(n_7427),
.Y(n_9780)
);

AND2x2_ASAP7_75t_L g9781 ( 
.A(n_8990),
.B(n_9013),
.Y(n_9781)
);

NAND2xp5_ASAP7_75t_L g9782 ( 
.A(n_9079),
.B(n_6806),
.Y(n_9782)
);

OAI22xp5_ASAP7_75t_L g9783 ( 
.A1(n_8944),
.A2(n_8354),
.B1(n_7959),
.B2(n_7960),
.Y(n_9783)
);

NAND2xp5_ASAP7_75t_L g9784 ( 
.A(n_9093),
.B(n_6806),
.Y(n_9784)
);

INVx2_ASAP7_75t_L g9785 ( 
.A(n_8566),
.Y(n_9785)
);

INVx2_ASAP7_75t_L g9786 ( 
.A(n_8566),
.Y(n_9786)
);

OAI22xp33_ASAP7_75t_L g9787 ( 
.A1(n_9002),
.A2(n_7223),
.B1(n_6617),
.B2(n_6773),
.Y(n_9787)
);

AOI22xp33_ASAP7_75t_L g9788 ( 
.A1(n_8749),
.A2(n_8012),
.B1(n_8105),
.B2(n_8089),
.Y(n_9788)
);

AOI221xp5_ASAP7_75t_L g9789 ( 
.A1(n_8384),
.A2(n_8353),
.B1(n_8352),
.B2(n_8350),
.C(n_7402),
.Y(n_9789)
);

OAI21xp33_ASAP7_75t_SL g9790 ( 
.A1(n_8356),
.A2(n_8315),
.B(n_6564),
.Y(n_9790)
);

INVx4_ASAP7_75t_L g9791 ( 
.A(n_8837),
.Y(n_9791)
);

AOI222xp33_ASAP7_75t_L g9792 ( 
.A1(n_8750),
.A2(n_7402),
.B1(n_6462),
.B2(n_7069),
.C1(n_6562),
.C2(n_8352),
.Y(n_9792)
);

INVx1_ASAP7_75t_L g9793 ( 
.A(n_8445),
.Y(n_9793)
);

AOI22xp33_ASAP7_75t_L g9794 ( 
.A1(n_8751),
.A2(n_8012),
.B1(n_8105),
.B2(n_8089),
.Y(n_9794)
);

OAI211xp5_ASAP7_75t_L g9795 ( 
.A1(n_8717),
.A2(n_7095),
.B(n_7253),
.C(n_8254),
.Y(n_9795)
);

AO21x2_ASAP7_75t_L g9796 ( 
.A1(n_8918),
.A2(n_8353),
.B(n_7862),
.Y(n_9796)
);

AOI22xp33_ASAP7_75t_SL g9797 ( 
.A1(n_8844),
.A2(n_6562),
.B1(n_6959),
.B2(n_6936),
.Y(n_9797)
);

OAI21x1_ASAP7_75t_L g9798 ( 
.A1(n_8722),
.A2(n_7427),
.B(n_7820),
.Y(n_9798)
);

OAI22xp5_ASAP7_75t_L g9799 ( 
.A1(n_8958),
.A2(n_8073),
.B1(n_7936),
.B2(n_7332),
.Y(n_9799)
);

AND2x2_ASAP7_75t_L g9800 ( 
.A(n_9013),
.B(n_8182),
.Y(n_9800)
);

AOI22xp33_ASAP7_75t_SL g9801 ( 
.A1(n_8844),
.A2(n_6959),
.B1(n_6988),
.B2(n_6936),
.Y(n_9801)
);

OR2x2_ASAP7_75t_L g9802 ( 
.A(n_9040),
.B(n_8300),
.Y(n_9802)
);

OAI22xp5_ASAP7_75t_L g9803 ( 
.A1(n_8973),
.A2(n_8073),
.B1(n_7936),
.B2(n_7332),
.Y(n_9803)
);

AOI22xp5_ASAP7_75t_L g9804 ( 
.A1(n_8851),
.A2(n_7024),
.B1(n_7132),
.B2(n_5833),
.Y(n_9804)
);

OAI22xp33_ASAP7_75t_L g9805 ( 
.A1(n_9002),
.A2(n_7223),
.B1(n_6617),
.B2(n_6773),
.Y(n_9805)
);

OR2x2_ASAP7_75t_L g9806 ( 
.A(n_8633),
.B(n_7069),
.Y(n_9806)
);

OAI22xp5_ASAP7_75t_L g9807 ( 
.A1(n_8973),
.A2(n_7298),
.B1(n_8071),
.B2(n_6581),
.Y(n_9807)
);

AOI22xp33_ASAP7_75t_L g9808 ( 
.A1(n_8754),
.A2(n_8012),
.B1(n_8105),
.B2(n_8089),
.Y(n_9808)
);

AND2x2_ASAP7_75t_L g9809 ( 
.A(n_9023),
.B(n_8182),
.Y(n_9809)
);

HB1xp67_ASAP7_75t_L g9810 ( 
.A(n_9100),
.Y(n_9810)
);

HB1xp67_ASAP7_75t_L g9811 ( 
.A(n_9122),
.Y(n_9811)
);

OAI22xp5_ASAP7_75t_L g9812 ( 
.A1(n_8975),
.A2(n_7298),
.B1(n_8071),
.B2(n_6581),
.Y(n_9812)
);

OR2x6_ASAP7_75t_L g9813 ( 
.A(n_8837),
.B(n_7647),
.Y(n_9813)
);

INVx3_ASAP7_75t_L g9814 ( 
.A(n_8911),
.Y(n_9814)
);

OAI22xp33_ASAP7_75t_L g9815 ( 
.A1(n_9002),
.A2(n_7223),
.B1(n_6617),
.B2(n_6773),
.Y(n_9815)
);

NAND2xp5_ASAP7_75t_L g9816 ( 
.A(n_8996),
.B(n_6806),
.Y(n_9816)
);

AOI22xp33_ASAP7_75t_SL g9817 ( 
.A1(n_8902),
.A2(n_6959),
.B1(n_6988),
.B2(n_6936),
.Y(n_9817)
);

AOI22xp33_ASAP7_75t_L g9818 ( 
.A1(n_8754),
.A2(n_8012),
.B1(n_8105),
.B2(n_8089),
.Y(n_9818)
);

OAI22xp5_ASAP7_75t_L g9819 ( 
.A1(n_8975),
.A2(n_9018),
.B1(n_9060),
.B2(n_8987),
.Y(n_9819)
);

AOI22xp33_ASAP7_75t_L g9820 ( 
.A1(n_8756),
.A2(n_8012),
.B1(n_8105),
.B2(n_8089),
.Y(n_9820)
);

INVx2_ASAP7_75t_L g9821 ( 
.A(n_8621),
.Y(n_9821)
);

OAI22xp33_ASAP7_75t_L g9822 ( 
.A1(n_8742),
.A2(n_6617),
.B1(n_6773),
.B2(n_6625),
.Y(n_9822)
);

INVx1_ASAP7_75t_L g9823 ( 
.A(n_8463),
.Y(n_9823)
);

INVx1_ASAP7_75t_L g9824 ( 
.A(n_8464),
.Y(n_9824)
);

AND2x2_ASAP7_75t_L g9825 ( 
.A(n_9023),
.B(n_8185),
.Y(n_9825)
);

AOI21xp33_ASAP7_75t_L g9826 ( 
.A1(n_8483),
.A2(n_8530),
.B(n_8987),
.Y(n_9826)
);

INVx4_ASAP7_75t_L g9827 ( 
.A(n_8837),
.Y(n_9827)
);

INVx1_ASAP7_75t_L g9828 ( 
.A(n_8466),
.Y(n_9828)
);

INVx1_ASAP7_75t_L g9829 ( 
.A(n_8469),
.Y(n_9829)
);

AND2x2_ASAP7_75t_L g9830 ( 
.A(n_8726),
.B(n_8185),
.Y(n_9830)
);

AOI22xp33_ASAP7_75t_L g9831 ( 
.A1(n_8756),
.A2(n_8105),
.B1(n_8151),
.B2(n_8113),
.Y(n_9831)
);

OA21x2_ASAP7_75t_L g9832 ( 
.A1(n_9145),
.A2(n_7833),
.B(n_7820),
.Y(n_9832)
);

NOR2xp67_ASAP7_75t_L g9833 ( 
.A(n_8717),
.B(n_8254),
.Y(n_9833)
);

AO21x2_ASAP7_75t_L g9834 ( 
.A1(n_8384),
.A2(n_7875),
.B(n_7854),
.Y(n_9834)
);

AOI21xp5_ASAP7_75t_L g9835 ( 
.A1(n_9039),
.A2(n_9046),
.B(n_8617),
.Y(n_9835)
);

AND2x2_ASAP7_75t_L g9836 ( 
.A(n_8726),
.B(n_8113),
.Y(n_9836)
);

NOR2xp33_ASAP7_75t_L g9837 ( 
.A(n_8717),
.B(n_7063),
.Y(n_9837)
);

OAI211xp5_ASAP7_75t_L g9838 ( 
.A1(n_9018),
.A2(n_7095),
.B(n_7253),
.C(n_8254),
.Y(n_9838)
);

INVx2_ASAP7_75t_SL g9839 ( 
.A(n_8621),
.Y(n_9839)
);

AND2x2_ASAP7_75t_L g9840 ( 
.A(n_8731),
.B(n_8113),
.Y(n_9840)
);

AOI22xp33_ASAP7_75t_L g9841 ( 
.A1(n_8759),
.A2(n_8113),
.B1(n_8206),
.B2(n_8151),
.Y(n_9841)
);

INVx1_ASAP7_75t_L g9842 ( 
.A(n_8485),
.Y(n_9842)
);

AND2x2_ASAP7_75t_L g9843 ( 
.A(n_8731),
.B(n_8113),
.Y(n_9843)
);

HB1xp67_ASAP7_75t_L g9844 ( 
.A(n_8600),
.Y(n_9844)
);

OR2x2_ASAP7_75t_L g9845 ( 
.A(n_8633),
.B(n_7325),
.Y(n_9845)
);

INVx1_ASAP7_75t_L g9846 ( 
.A(n_9185),
.Y(n_9846)
);

INVx2_ASAP7_75t_L g9847 ( 
.A(n_9424),
.Y(n_9847)
);

HB1xp67_ASAP7_75t_L g9848 ( 
.A(n_9167),
.Y(n_9848)
);

NAND2x1_ASAP7_75t_L g9849 ( 
.A(n_9470),
.B(n_9080),
.Y(n_9849)
);

INVx2_ASAP7_75t_L g9850 ( 
.A(n_9474),
.Y(n_9850)
);

OR2x2_ASAP7_75t_L g9851 ( 
.A(n_9290),
.B(n_8645),
.Y(n_9851)
);

NAND2xp5_ASAP7_75t_L g9852 ( 
.A(n_9213),
.B(n_8488),
.Y(n_9852)
);

INVx1_ASAP7_75t_L g9853 ( 
.A(n_9363),
.Y(n_9853)
);

INVx2_ASAP7_75t_L g9854 ( 
.A(n_9375),
.Y(n_9854)
);

OR2x2_ASAP7_75t_L g9855 ( 
.A(n_9193),
.B(n_8645),
.Y(n_9855)
);

NOR2xp33_ASAP7_75t_L g9856 ( 
.A(n_9351),
.B(n_8621),
.Y(n_9856)
);

AND2x2_ASAP7_75t_L g9857 ( 
.A(n_9259),
.B(n_9010),
.Y(n_9857)
);

INVx2_ASAP7_75t_L g9858 ( 
.A(n_9164),
.Y(n_9858)
);

INVx1_ASAP7_75t_L g9859 ( 
.A(n_9452),
.Y(n_9859)
);

INVx1_ASAP7_75t_L g9860 ( 
.A(n_9489),
.Y(n_9860)
);

AND2x2_ASAP7_75t_L g9861 ( 
.A(n_9259),
.B(n_9010),
.Y(n_9861)
);

AND2x2_ASAP7_75t_L g9862 ( 
.A(n_9563),
.B(n_8532),
.Y(n_9862)
);

AND2x4_ASAP7_75t_L g9863 ( 
.A(n_9168),
.B(n_8921),
.Y(n_9863)
);

AND2x2_ASAP7_75t_L g9864 ( 
.A(n_9365),
.B(n_8532),
.Y(n_9864)
);

INVx2_ASAP7_75t_L g9865 ( 
.A(n_9230),
.Y(n_9865)
);

INVx2_ASAP7_75t_L g9866 ( 
.A(n_9230),
.Y(n_9866)
);

HB1xp67_ASAP7_75t_L g9867 ( 
.A(n_9844),
.Y(n_9867)
);

INVx1_ASAP7_75t_L g9868 ( 
.A(n_9584),
.Y(n_9868)
);

AND2x2_ASAP7_75t_L g9869 ( 
.A(n_9177),
.B(n_8617),
.Y(n_9869)
);

INVx2_ASAP7_75t_L g9870 ( 
.A(n_9273),
.Y(n_9870)
);

INVx1_ASAP7_75t_L g9871 ( 
.A(n_9622),
.Y(n_9871)
);

INVx1_ASAP7_75t_SL g9872 ( 
.A(n_9310),
.Y(n_9872)
);

BUFx2_ASAP7_75t_L g9873 ( 
.A(n_9256),
.Y(n_9873)
);

INVx2_ASAP7_75t_L g9874 ( 
.A(n_9273),
.Y(n_9874)
);

INVx1_ASAP7_75t_L g9875 ( 
.A(n_9638),
.Y(n_9875)
);

INVx3_ASAP7_75t_L g9876 ( 
.A(n_9351),
.Y(n_9876)
);

AND2x2_ASAP7_75t_L g9877 ( 
.A(n_9180),
.B(n_8821),
.Y(n_9877)
);

INVx1_ASAP7_75t_L g9878 ( 
.A(n_9651),
.Y(n_9878)
);

AND2x4_ASAP7_75t_L g9879 ( 
.A(n_9216),
.B(n_8926),
.Y(n_9879)
);

INVx1_ASAP7_75t_L g9880 ( 
.A(n_9688),
.Y(n_9880)
);

INVx3_ASAP7_75t_L g9881 ( 
.A(n_9351),
.Y(n_9881)
);

INVx1_ASAP7_75t_L g9882 ( 
.A(n_9734),
.Y(n_9882)
);

HB1xp67_ASAP7_75t_L g9883 ( 
.A(n_9380),
.Y(n_9883)
);

INVx1_ASAP7_75t_L g9884 ( 
.A(n_9740),
.Y(n_9884)
);

BUFx3_ASAP7_75t_L g9885 ( 
.A(n_9256),
.Y(n_9885)
);

AND2x2_ASAP7_75t_L g9886 ( 
.A(n_9329),
.B(n_8821),
.Y(n_9886)
);

INVx1_ASAP7_75t_L g9887 ( 
.A(n_9768),
.Y(n_9887)
);

NAND2x1p5_ASAP7_75t_L g9888 ( 
.A(n_9602),
.B(n_8621),
.Y(n_9888)
);

INVx1_ASAP7_75t_L g9889 ( 
.A(n_9776),
.Y(n_9889)
);

OR2x2_ASAP7_75t_L g9890 ( 
.A(n_9348),
.B(n_8600),
.Y(n_9890)
);

INVx2_ASAP7_75t_L g9891 ( 
.A(n_9295),
.Y(n_9891)
);

AND2x4_ASAP7_75t_SL g9892 ( 
.A(n_9381),
.B(n_8621),
.Y(n_9892)
);

INVx2_ASAP7_75t_L g9893 ( 
.A(n_9729),
.Y(n_9893)
);

NAND2xp5_ASAP7_75t_L g9894 ( 
.A(n_9324),
.B(n_8497),
.Y(n_9894)
);

INVx1_ASAP7_75t_L g9895 ( 
.A(n_9810),
.Y(n_9895)
);

HB1xp67_ASAP7_75t_L g9896 ( 
.A(n_9205),
.Y(n_9896)
);

AND2x2_ASAP7_75t_L g9897 ( 
.A(n_9302),
.B(n_8840),
.Y(n_9897)
);

HB1xp67_ASAP7_75t_L g9898 ( 
.A(n_9811),
.Y(n_9898)
);

INVx1_ASAP7_75t_L g9899 ( 
.A(n_9182),
.Y(n_9899)
);

BUFx2_ASAP7_75t_L g9900 ( 
.A(n_9381),
.Y(n_9900)
);

INVx1_ASAP7_75t_L g9901 ( 
.A(n_9184),
.Y(n_9901)
);

INVx2_ASAP7_75t_L g9902 ( 
.A(n_9165),
.Y(n_9902)
);

AND2x2_ASAP7_75t_L g9903 ( 
.A(n_9312),
.B(n_8840),
.Y(n_9903)
);

INVx2_ASAP7_75t_L g9904 ( 
.A(n_9586),
.Y(n_9904)
);

INVx3_ASAP7_75t_L g9905 ( 
.A(n_9381),
.Y(n_9905)
);

BUFx4f_ASAP7_75t_SL g9906 ( 
.A(n_9492),
.Y(n_9906)
);

INVx4_ASAP7_75t_L g9907 ( 
.A(n_9448),
.Y(n_9907)
);

AND2x2_ASAP7_75t_L g9908 ( 
.A(n_9321),
.B(n_8926),
.Y(n_9908)
);

INVx1_ASAP7_75t_L g9909 ( 
.A(n_9186),
.Y(n_9909)
);

NAND2xp5_ASAP7_75t_L g9910 ( 
.A(n_9324),
.B(n_8498),
.Y(n_9910)
);

AND2x2_ASAP7_75t_L g9911 ( 
.A(n_9330),
.B(n_8988),
.Y(n_9911)
);

INVx1_ASAP7_75t_L g9912 ( 
.A(n_9192),
.Y(n_9912)
);

INVx1_ASAP7_75t_L g9913 ( 
.A(n_9206),
.Y(n_9913)
);

AND2x2_ASAP7_75t_L g9914 ( 
.A(n_9170),
.B(n_8988),
.Y(n_9914)
);

AND2x2_ASAP7_75t_L g9915 ( 
.A(n_9581),
.B(n_9781),
.Y(n_9915)
);

INVx1_ASAP7_75t_L g9916 ( 
.A(n_9211),
.Y(n_9916)
);

BUFx2_ASAP7_75t_L g9917 ( 
.A(n_9202),
.Y(n_9917)
);

AND2x2_ASAP7_75t_L g9918 ( 
.A(n_9436),
.B(n_9097),
.Y(n_9918)
);

INVx1_ASAP7_75t_L g9919 ( 
.A(n_9217),
.Y(n_9919)
);

OR2x2_ASAP7_75t_L g9920 ( 
.A(n_9191),
.B(n_8600),
.Y(n_9920)
);

HB1xp67_ASAP7_75t_L g9921 ( 
.A(n_9165),
.Y(n_9921)
);

INVx3_ASAP7_75t_L g9922 ( 
.A(n_9516),
.Y(n_9922)
);

INVx1_ASAP7_75t_L g9923 ( 
.A(n_9225),
.Y(n_9923)
);

INVx2_ASAP7_75t_L g9924 ( 
.A(n_9621),
.Y(n_9924)
);

AND2x2_ASAP7_75t_L g9925 ( 
.A(n_9559),
.B(n_9097),
.Y(n_9925)
);

NAND2xp5_ASAP7_75t_L g9926 ( 
.A(n_9190),
.B(n_8500),
.Y(n_9926)
);

INVx2_ASAP7_75t_L g9927 ( 
.A(n_9628),
.Y(n_9927)
);

OR2x2_ASAP7_75t_L g9928 ( 
.A(n_9242),
.B(n_8600),
.Y(n_9928)
);

INVx3_ASAP7_75t_L g9929 ( 
.A(n_9271),
.Y(n_9929)
);

AND2x2_ASAP7_75t_L g9930 ( 
.A(n_9521),
.B(n_9127),
.Y(n_9930)
);

INVx2_ASAP7_75t_SL g9931 ( 
.A(n_9417),
.Y(n_9931)
);

INVx2_ASAP7_75t_L g9932 ( 
.A(n_9836),
.Y(n_9932)
);

INVx1_ASAP7_75t_L g9933 ( 
.A(n_9229),
.Y(n_9933)
);

INVx1_ASAP7_75t_L g9934 ( 
.A(n_9238),
.Y(n_9934)
);

OAI21xp33_ASAP7_75t_L g9935 ( 
.A1(n_9432),
.A2(n_9127),
.B(n_8542),
.Y(n_9935)
);

INVx1_ASAP7_75t_L g9936 ( 
.A(n_9246),
.Y(n_9936)
);

INVx2_ASAP7_75t_L g9937 ( 
.A(n_9840),
.Y(n_9937)
);

BUFx3_ASAP7_75t_L g9938 ( 
.A(n_9172),
.Y(n_9938)
);

INVx2_ASAP7_75t_L g9939 ( 
.A(n_9843),
.Y(n_9939)
);

INVx2_ASAP7_75t_L g9940 ( 
.A(n_9165),
.Y(n_9940)
);

INVx2_ASAP7_75t_L g9941 ( 
.A(n_9385),
.Y(n_9941)
);

INVx1_ASAP7_75t_L g9942 ( 
.A(n_9248),
.Y(n_9942)
);

INVx2_ASAP7_75t_L g9943 ( 
.A(n_9641),
.Y(n_9943)
);

INVx2_ASAP7_75t_L g9944 ( 
.A(n_9653),
.Y(n_9944)
);

HB1xp67_ASAP7_75t_L g9945 ( 
.A(n_9247),
.Y(n_9945)
);

INVx1_ASAP7_75t_L g9946 ( 
.A(n_9250),
.Y(n_9946)
);

INVx1_ASAP7_75t_L g9947 ( 
.A(n_9253),
.Y(n_9947)
);

OR2x2_ASAP7_75t_L g9948 ( 
.A(n_9183),
.B(n_8600),
.Y(n_9948)
);

OR2x2_ASAP7_75t_L g9949 ( 
.A(n_9421),
.B(n_9453),
.Y(n_9949)
);

INVx1_ASAP7_75t_L g9950 ( 
.A(n_9270),
.Y(n_9950)
);

BUFx6f_ASAP7_75t_L g9951 ( 
.A(n_9271),
.Y(n_9951)
);

HB1xp67_ASAP7_75t_L g9952 ( 
.A(n_9212),
.Y(n_9952)
);

INVx2_ASAP7_75t_L g9953 ( 
.A(n_9655),
.Y(n_9953)
);

INVx2_ASAP7_75t_L g9954 ( 
.A(n_9271),
.Y(n_9954)
);

BUFx2_ASAP7_75t_L g9955 ( 
.A(n_9202),
.Y(n_9955)
);

AND2x2_ASAP7_75t_L g9956 ( 
.A(n_9334),
.B(n_8483),
.Y(n_9956)
);

AND2x2_ASAP7_75t_L g9957 ( 
.A(n_9337),
.B(n_8530),
.Y(n_9957)
);

HB1xp67_ASAP7_75t_L g9958 ( 
.A(n_9226),
.Y(n_9958)
);

INVx1_ASAP7_75t_L g9959 ( 
.A(n_9280),
.Y(n_9959)
);

INVx2_ASAP7_75t_L g9960 ( 
.A(n_9204),
.Y(n_9960)
);

NAND2xp5_ASAP7_75t_L g9961 ( 
.A(n_9190),
.B(n_8506),
.Y(n_9961)
);

AND2x2_ASAP7_75t_L g9962 ( 
.A(n_9519),
.B(n_8996),
.Y(n_9962)
);

INVx1_ASAP7_75t_L g9963 ( 
.A(n_9287),
.Y(n_9963)
);

HB1xp67_ASAP7_75t_L g9964 ( 
.A(n_9228),
.Y(n_9964)
);

BUFx3_ASAP7_75t_L g9965 ( 
.A(n_9507),
.Y(n_9965)
);

AND2x2_ASAP7_75t_L g9966 ( 
.A(n_9419),
.B(n_8996),
.Y(n_9966)
);

OR2x2_ASAP7_75t_L g9967 ( 
.A(n_9510),
.B(n_8471),
.Y(n_9967)
);

INVx1_ASAP7_75t_L g9968 ( 
.A(n_9327),
.Y(n_9968)
);

AND2x2_ASAP7_75t_L g9969 ( 
.A(n_9529),
.B(n_8996),
.Y(n_9969)
);

OR2x2_ASAP7_75t_L g9970 ( 
.A(n_9220),
.B(n_9802),
.Y(n_9970)
);

AND2x4_ASAP7_75t_L g9971 ( 
.A(n_9216),
.B(n_8642),
.Y(n_9971)
);

AND2x2_ASAP7_75t_L g9972 ( 
.A(n_9543),
.B(n_8996),
.Y(n_9972)
);

INVx2_ASAP7_75t_L g9973 ( 
.A(n_9207),
.Y(n_9973)
);

INVx1_ASAP7_75t_L g9974 ( 
.A(n_9335),
.Y(n_9974)
);

AND2x2_ASAP7_75t_L g9975 ( 
.A(n_9555),
.B(n_8642),
.Y(n_9975)
);

INVx1_ASAP7_75t_L g9976 ( 
.A(n_9336),
.Y(n_9976)
);

OR2x2_ASAP7_75t_L g9977 ( 
.A(n_9534),
.B(n_8471),
.Y(n_9977)
);

INVx3_ASAP7_75t_L g9978 ( 
.A(n_9430),
.Y(n_9978)
);

NAND2xp5_ASAP7_75t_L g9979 ( 
.A(n_9235),
.B(n_8511),
.Y(n_9979)
);

AND2x2_ASAP7_75t_L g9980 ( 
.A(n_9388),
.B(n_8642),
.Y(n_9980)
);

INVx2_ASAP7_75t_L g9981 ( 
.A(n_9262),
.Y(n_9981)
);

INVx1_ASAP7_75t_L g9982 ( 
.A(n_9353),
.Y(n_9982)
);

INVx2_ASAP7_75t_L g9983 ( 
.A(n_9796),
.Y(n_9983)
);

AND2x2_ASAP7_75t_L g9984 ( 
.A(n_9398),
.B(n_8642),
.Y(n_9984)
);

AND2x2_ASAP7_75t_L g9985 ( 
.A(n_9447),
.B(n_8642),
.Y(n_9985)
);

AND2x2_ASAP7_75t_L g9986 ( 
.A(n_9281),
.B(n_8647),
.Y(n_9986)
);

INVx1_ASAP7_75t_L g9987 ( 
.A(n_9366),
.Y(n_9987)
);

INVx2_ASAP7_75t_L g9988 ( 
.A(n_9263),
.Y(n_9988)
);

AND2x2_ASAP7_75t_L g9989 ( 
.A(n_9288),
.B(n_8647),
.Y(n_9989)
);

INVx2_ASAP7_75t_L g9990 ( 
.A(n_9796),
.Y(n_9990)
);

NAND2x1p5_ASAP7_75t_L g9991 ( 
.A(n_9602),
.B(n_8647),
.Y(n_9991)
);

AND2x2_ASAP7_75t_L g9992 ( 
.A(n_9300),
.B(n_8647),
.Y(n_9992)
);

NOR2xp67_ASAP7_75t_SL g9993 ( 
.A(n_9658),
.B(n_8647),
.Y(n_9993)
);

INVx1_ASAP7_75t_L g9994 ( 
.A(n_9368),
.Y(n_9994)
);

OR2x2_ASAP7_75t_L g9995 ( 
.A(n_9618),
.B(n_8512),
.Y(n_9995)
);

OR2x2_ASAP7_75t_L g9996 ( 
.A(n_9241),
.B(n_8515),
.Y(n_9996)
);

BUFx2_ASAP7_75t_L g9997 ( 
.A(n_9370),
.Y(n_9997)
);

HB1xp67_ASAP7_75t_L g9998 ( 
.A(n_9231),
.Y(n_9998)
);

OR2x2_ASAP7_75t_L g9999 ( 
.A(n_9171),
.B(n_8518),
.Y(n_9999)
);

AND2x2_ASAP7_75t_L g10000 ( 
.A(n_9301),
.B(n_9060),
.Y(n_10000)
);

INVx3_ASAP7_75t_L g10001 ( 
.A(n_9634),
.Y(n_10001)
);

INVx2_ASAP7_75t_L g10002 ( 
.A(n_9515),
.Y(n_10002)
);

AND2x2_ASAP7_75t_L g10003 ( 
.A(n_9689),
.B(n_9143),
.Y(n_10003)
);

BUFx3_ASAP7_75t_L g10004 ( 
.A(n_9553),
.Y(n_10004)
);

INVx1_ASAP7_75t_L g10005 ( 
.A(n_9379),
.Y(n_10005)
);

OR2x2_ASAP7_75t_L g10006 ( 
.A(n_9178),
.B(n_8522),
.Y(n_10006)
);

HB1xp67_ASAP7_75t_L g10007 ( 
.A(n_9234),
.Y(n_10007)
);

INVxp67_ASAP7_75t_L g10008 ( 
.A(n_9428),
.Y(n_10008)
);

AO31x2_ASAP7_75t_L g10009 ( 
.A1(n_9163),
.A2(n_9121),
.A3(n_8391),
.B(n_8398),
.Y(n_10009)
);

HB1xp67_ASAP7_75t_L g10010 ( 
.A(n_9283),
.Y(n_10010)
);

INVx3_ASAP7_75t_L g10011 ( 
.A(n_9741),
.Y(n_10011)
);

AND2x2_ASAP7_75t_L g10012 ( 
.A(n_9411),
.B(n_9143),
.Y(n_10012)
);

NAND2xp5_ASAP7_75t_L g10013 ( 
.A(n_9235),
.B(n_8526),
.Y(n_10013)
);

INVx2_ASAP7_75t_L g10014 ( 
.A(n_9834),
.Y(n_10014)
);

AND2x4_ASAP7_75t_L g10015 ( 
.A(n_9255),
.B(n_8911),
.Y(n_10015)
);

OR2x2_ASAP7_75t_L g10016 ( 
.A(n_9705),
.B(n_8527),
.Y(n_10016)
);

OR2x2_ASAP7_75t_L g10017 ( 
.A(n_9674),
.B(n_8528),
.Y(n_10017)
);

BUFx2_ASAP7_75t_L g10018 ( 
.A(n_9293),
.Y(n_10018)
);

INVx1_ASAP7_75t_L g10019 ( 
.A(n_9395),
.Y(n_10019)
);

INVx1_ASAP7_75t_L g10020 ( 
.A(n_9403),
.Y(n_10020)
);

AND2x2_ASAP7_75t_L g10021 ( 
.A(n_9411),
.B(n_8930),
.Y(n_10021)
);

INVx2_ASAP7_75t_L g10022 ( 
.A(n_9834),
.Y(n_10022)
);

INVx2_ASAP7_75t_L g10023 ( 
.A(n_9572),
.Y(n_10023)
);

AND2x2_ASAP7_75t_L g10024 ( 
.A(n_9411),
.B(n_8930),
.Y(n_10024)
);

OR2x2_ASAP7_75t_L g10025 ( 
.A(n_9303),
.B(n_8529),
.Y(n_10025)
);

OR2x2_ASAP7_75t_L g10026 ( 
.A(n_9201),
.B(n_8534),
.Y(n_10026)
);

INVx1_ASAP7_75t_L g10027 ( 
.A(n_9404),
.Y(n_10027)
);

AND2x2_ASAP7_75t_L g10028 ( 
.A(n_9813),
.B(n_8113),
.Y(n_10028)
);

NOR2x1_ASAP7_75t_L g10029 ( 
.A(n_9608),
.B(n_9061),
.Y(n_10029)
);

AND2x2_ASAP7_75t_L g10030 ( 
.A(n_9813),
.B(n_8151),
.Y(n_10030)
);

INVx1_ASAP7_75t_L g10031 ( 
.A(n_9409),
.Y(n_10031)
);

INVxp67_ASAP7_75t_SL g10032 ( 
.A(n_9537),
.Y(n_10032)
);

INVx2_ASAP7_75t_L g10033 ( 
.A(n_9626),
.Y(n_10033)
);

INVxp67_ASAP7_75t_SL g10034 ( 
.A(n_9289),
.Y(n_10034)
);

NAND2xp5_ASAP7_75t_L g10035 ( 
.A(n_9198),
.B(n_8546),
.Y(n_10035)
);

OR2x2_ASAP7_75t_L g10036 ( 
.A(n_9215),
.B(n_8549),
.Y(n_10036)
);

NAND2xp5_ASAP7_75t_L g10037 ( 
.A(n_9224),
.B(n_9527),
.Y(n_10037)
);

NOR2xp33_ASAP7_75t_L g10038 ( 
.A(n_9390),
.B(n_9349),
.Y(n_10038)
);

HB1xp67_ASAP7_75t_L g10039 ( 
.A(n_9284),
.Y(n_10039)
);

AND2x2_ASAP7_75t_L g10040 ( 
.A(n_9813),
.B(n_8151),
.Y(n_10040)
);

INVx2_ASAP7_75t_L g10041 ( 
.A(n_9629),
.Y(n_10041)
);

INVx2_ASAP7_75t_L g10042 ( 
.A(n_9656),
.Y(n_10042)
);

OR2x2_ASAP7_75t_L g10043 ( 
.A(n_9631),
.B(n_8550),
.Y(n_10043)
);

NAND2xp5_ASAP7_75t_L g10044 ( 
.A(n_9197),
.B(n_8552),
.Y(n_10044)
);

INVx1_ASAP7_75t_L g10045 ( 
.A(n_9425),
.Y(n_10045)
);

AND2x2_ASAP7_75t_L g10046 ( 
.A(n_9830),
.B(n_8151),
.Y(n_10046)
);

OR2x2_ASAP7_75t_L g10047 ( 
.A(n_9639),
.B(n_9680),
.Y(n_10047)
);

BUFx2_ASAP7_75t_L g10048 ( 
.A(n_9742),
.Y(n_10048)
);

INVx1_ASAP7_75t_L g10049 ( 
.A(n_9435),
.Y(n_10049)
);

OR2x2_ASAP7_75t_L g10050 ( 
.A(n_9360),
.B(n_8555),
.Y(n_10050)
);

INVx2_ASAP7_75t_L g10051 ( 
.A(n_9700),
.Y(n_10051)
);

AND2x2_ASAP7_75t_L g10052 ( 
.A(n_9440),
.B(n_8151),
.Y(n_10052)
);

NAND2xp5_ASAP7_75t_L g10053 ( 
.A(n_9189),
.B(n_8559),
.Y(n_10053)
);

HB1xp67_ASAP7_75t_L g10054 ( 
.A(n_9284),
.Y(n_10054)
);

AND2x2_ASAP7_75t_L g10055 ( 
.A(n_9443),
.B(n_8206),
.Y(n_10055)
);

NAND2xp5_ASAP7_75t_L g10056 ( 
.A(n_9498),
.B(n_8569),
.Y(n_10056)
);

AND2x4_ASAP7_75t_L g10057 ( 
.A(n_9255),
.B(n_8742),
.Y(n_10057)
);

INVx1_ASAP7_75t_L g10058 ( 
.A(n_9439),
.Y(n_10058)
);

INVx1_ASAP7_75t_L g10059 ( 
.A(n_9441),
.Y(n_10059)
);

BUFx6f_ASAP7_75t_L g10060 ( 
.A(n_9428),
.Y(n_10060)
);

INVx2_ASAP7_75t_SL g10061 ( 
.A(n_9428),
.Y(n_10061)
);

AND2x2_ASAP7_75t_L g10062 ( 
.A(n_9665),
.B(n_8206),
.Y(n_10062)
);

INVx2_ASAP7_75t_L g10063 ( 
.A(n_9701),
.Y(n_10063)
);

INVx1_ASAP7_75t_L g10064 ( 
.A(n_9446),
.Y(n_10064)
);

INVx5_ASAP7_75t_L g10065 ( 
.A(n_9490),
.Y(n_10065)
);

INVx1_ASAP7_75t_L g10066 ( 
.A(n_9454),
.Y(n_10066)
);

OR2x2_ASAP7_75t_L g10067 ( 
.A(n_9309),
.B(n_8573),
.Y(n_10067)
);

INVx1_ASAP7_75t_L g10068 ( 
.A(n_9463),
.Y(n_10068)
);

INVx1_ASAP7_75t_L g10069 ( 
.A(n_9466),
.Y(n_10069)
);

INVx2_ASAP7_75t_L g10070 ( 
.A(n_9715),
.Y(n_10070)
);

AND2x2_ASAP7_75t_L g10071 ( 
.A(n_9763),
.B(n_8206),
.Y(n_10071)
);

NAND2x1p5_ASAP7_75t_L g10072 ( 
.A(n_9602),
.B(n_9552),
.Y(n_10072)
);

INVx1_ASAP7_75t_L g10073 ( 
.A(n_9484),
.Y(n_10073)
);

AND2x2_ASAP7_75t_L g10074 ( 
.A(n_9800),
.B(n_8206),
.Y(n_10074)
);

AND2x2_ASAP7_75t_L g10075 ( 
.A(n_9809),
.B(n_8206),
.Y(n_10075)
);

INVx2_ASAP7_75t_L g10076 ( 
.A(n_9717),
.Y(n_10076)
);

INVx1_ASAP7_75t_L g10077 ( 
.A(n_9522),
.Y(n_10077)
);

INVx2_ASAP7_75t_L g10078 ( 
.A(n_9730),
.Y(n_10078)
);

INVx1_ASAP7_75t_L g10079 ( 
.A(n_9525),
.Y(n_10079)
);

AND2x2_ASAP7_75t_L g10080 ( 
.A(n_9825),
.B(n_8210),
.Y(n_10080)
);

NOR2xp33_ASAP7_75t_L g10081 ( 
.A(n_9551),
.B(n_5810),
.Y(n_10081)
);

AOI22xp33_ASAP7_75t_L g10082 ( 
.A1(n_9194),
.A2(n_8765),
.B1(n_8773),
.B2(n_8759),
.Y(n_10082)
);

AND2x2_ASAP7_75t_L g10083 ( 
.A(n_9690),
.B(n_8210),
.Y(n_10083)
);

INVx1_ASAP7_75t_L g10084 ( 
.A(n_9531),
.Y(n_10084)
);

HB1xp67_ASAP7_75t_L g10085 ( 
.A(n_9364),
.Y(n_10085)
);

OR2x2_ASAP7_75t_L g10086 ( 
.A(n_9318),
.B(n_8575),
.Y(n_10086)
);

AND2x2_ASAP7_75t_L g10087 ( 
.A(n_9243),
.B(n_8210),
.Y(n_10087)
);

INVx2_ASAP7_75t_L g10088 ( 
.A(n_9751),
.Y(n_10088)
);

BUFx3_ASAP7_75t_L g10089 ( 
.A(n_9721),
.Y(n_10089)
);

AND2x2_ASAP7_75t_L g10090 ( 
.A(n_9450),
.B(n_8210),
.Y(n_10090)
);

AO31x2_ASAP7_75t_L g10091 ( 
.A1(n_9386),
.A2(n_8391),
.A3(n_8398),
.B(n_8385),
.Y(n_10091)
);

AND2x2_ASAP7_75t_L g10092 ( 
.A(n_9451),
.B(n_8210),
.Y(n_10092)
);

INVx1_ASAP7_75t_L g10093 ( 
.A(n_9535),
.Y(n_10093)
);

INVx2_ASAP7_75t_L g10094 ( 
.A(n_9764),
.Y(n_10094)
);

OR2x2_ASAP7_75t_L g10095 ( 
.A(n_9723),
.B(n_8582),
.Y(n_10095)
);

AND2x4_ASAP7_75t_L g10096 ( 
.A(n_9596),
.B(n_8742),
.Y(n_10096)
);

AND2x2_ASAP7_75t_SL g10097 ( 
.A(n_9233),
.B(n_8210),
.Y(n_10097)
);

AND2x2_ASAP7_75t_L g10098 ( 
.A(n_9316),
.B(n_8215),
.Y(n_10098)
);

INVx1_ASAP7_75t_L g10099 ( 
.A(n_9556),
.Y(n_10099)
);

AND2x2_ASAP7_75t_L g10100 ( 
.A(n_9316),
.B(n_8215),
.Y(n_10100)
);

INVx1_ASAP7_75t_L g10101 ( 
.A(n_9570),
.Y(n_10101)
);

INVx1_ASAP7_75t_L g10102 ( 
.A(n_9589),
.Y(n_10102)
);

NAND2xp5_ASAP7_75t_L g10103 ( 
.A(n_9498),
.B(n_8583),
.Y(n_10103)
);

INVxp67_ASAP7_75t_SL g10104 ( 
.A(n_9347),
.Y(n_10104)
);

AND2x2_ASAP7_75t_L g10105 ( 
.A(n_9285),
.B(n_9431),
.Y(n_10105)
);

INVx1_ASAP7_75t_L g10106 ( 
.A(n_9610),
.Y(n_10106)
);

HB1xp67_ASAP7_75t_L g10107 ( 
.A(n_9209),
.Y(n_10107)
);

INVx2_ASAP7_75t_L g10108 ( 
.A(n_9785),
.Y(n_10108)
);

INVx1_ASAP7_75t_L g10109 ( 
.A(n_9615),
.Y(n_10109)
);

INVx1_ASAP7_75t_L g10110 ( 
.A(n_9642),
.Y(n_10110)
);

AND2x2_ASAP7_75t_L g10111 ( 
.A(n_9285),
.B(n_8215),
.Y(n_10111)
);

INVx2_ASAP7_75t_SL g10112 ( 
.A(n_9490),
.Y(n_10112)
);

AND2x2_ASAP7_75t_L g10113 ( 
.A(n_9285),
.B(n_9431),
.Y(n_10113)
);

HB1xp67_ASAP7_75t_L g10114 ( 
.A(n_9209),
.Y(n_10114)
);

INVx2_ASAP7_75t_L g10115 ( 
.A(n_9786),
.Y(n_10115)
);

INVx2_ASAP7_75t_L g10116 ( 
.A(n_9821),
.Y(n_10116)
);

HB1xp67_ASAP7_75t_L g10117 ( 
.A(n_9393),
.Y(n_10117)
);

INVx1_ASAP7_75t_L g10118 ( 
.A(n_9643),
.Y(n_10118)
);

INVx1_ASAP7_75t_L g10119 ( 
.A(n_9650),
.Y(n_10119)
);

OR2x2_ASAP7_75t_L g10120 ( 
.A(n_9845),
.B(n_8584),
.Y(n_10120)
);

INVx1_ASAP7_75t_L g10121 ( 
.A(n_9672),
.Y(n_10121)
);

INVx1_ASAP7_75t_L g10122 ( 
.A(n_9697),
.Y(n_10122)
);

AND2x2_ASAP7_75t_L g10123 ( 
.A(n_9431),
.B(n_9606),
.Y(n_10123)
);

INVx2_ASAP7_75t_L g10124 ( 
.A(n_9208),
.Y(n_10124)
);

INVx2_ASAP7_75t_SL g10125 ( 
.A(n_9490),
.Y(n_10125)
);

INVx3_ASAP7_75t_L g10126 ( 
.A(n_9320),
.Y(n_10126)
);

INVxp67_ASAP7_75t_SL g10127 ( 
.A(n_9175),
.Y(n_10127)
);

OR2x2_ASAP7_75t_L g10128 ( 
.A(n_9277),
.B(n_8593),
.Y(n_10128)
);

INVx1_ASAP7_75t_L g10129 ( 
.A(n_9708),
.Y(n_10129)
);

BUFx2_ASAP7_75t_L g10130 ( 
.A(n_9518),
.Y(n_10130)
);

AND2x2_ASAP7_75t_L g10131 ( 
.A(n_9606),
.B(n_8215),
.Y(n_10131)
);

CKINVDCx16_ASAP7_75t_R g10132 ( 
.A(n_9166),
.Y(n_10132)
);

INVx2_ASAP7_75t_L g10133 ( 
.A(n_9839),
.Y(n_10133)
);

INVx3_ASAP7_75t_L g10134 ( 
.A(n_9320),
.Y(n_10134)
);

NAND2xp5_ASAP7_75t_L g10135 ( 
.A(n_9179),
.B(n_8596),
.Y(n_10135)
);

INVxp67_ASAP7_75t_L g10136 ( 
.A(n_9616),
.Y(n_10136)
);

NAND2xp5_ASAP7_75t_L g10137 ( 
.A(n_9376),
.B(n_8597),
.Y(n_10137)
);

OR2x2_ASAP7_75t_L g10138 ( 
.A(n_9245),
.B(n_8599),
.Y(n_10138)
);

INVx1_ASAP7_75t_L g10139 ( 
.A(n_9714),
.Y(n_10139)
);

INVx1_ASAP7_75t_L g10140 ( 
.A(n_9728),
.Y(n_10140)
);

INVx2_ASAP7_75t_L g10141 ( 
.A(n_9736),
.Y(n_10141)
);

INVx3_ASAP7_75t_L g10142 ( 
.A(n_9538),
.Y(n_10142)
);

HB1xp67_ASAP7_75t_L g10143 ( 
.A(n_9434),
.Y(n_10143)
);

AND2x2_ASAP7_75t_L g10144 ( 
.A(n_9606),
.B(n_8215),
.Y(n_10144)
);

INVx1_ASAP7_75t_L g10145 ( 
.A(n_9732),
.Y(n_10145)
);

INVx1_ASAP7_75t_L g10146 ( 
.A(n_9793),
.Y(n_10146)
);

BUFx6f_ASAP7_75t_L g10147 ( 
.A(n_9538),
.Y(n_10147)
);

INVx2_ASAP7_75t_L g10148 ( 
.A(n_9736),
.Y(n_10148)
);

NAND2xp5_ASAP7_75t_L g10149 ( 
.A(n_9272),
.B(n_8604),
.Y(n_10149)
);

AND2x2_ASAP7_75t_L g10150 ( 
.A(n_9350),
.B(n_8215),
.Y(n_10150)
);

NAND2xp5_ASAP7_75t_L g10151 ( 
.A(n_9372),
.B(n_8606),
.Y(n_10151)
);

AND2x2_ASAP7_75t_L g10152 ( 
.A(n_9362),
.B(n_8224),
.Y(n_10152)
);

INVx1_ASAP7_75t_L g10153 ( 
.A(n_9823),
.Y(n_10153)
);

INVx1_ASAP7_75t_L g10154 ( 
.A(n_9824),
.Y(n_10154)
);

NAND2xp5_ASAP7_75t_L g10155 ( 
.A(n_9372),
.B(n_8628),
.Y(n_10155)
);

AND2x2_ASAP7_75t_L g10156 ( 
.A(n_9367),
.B(n_8224),
.Y(n_10156)
);

AND2x2_ASAP7_75t_L g10157 ( 
.A(n_9373),
.B(n_8224),
.Y(n_10157)
);

INVx1_ASAP7_75t_L g10158 ( 
.A(n_9828),
.Y(n_10158)
);

INVx2_ASAP7_75t_L g10159 ( 
.A(n_9467),
.Y(n_10159)
);

INVx3_ASAP7_75t_L g10160 ( 
.A(n_9538),
.Y(n_10160)
);

INVx4_ASAP7_75t_L g10161 ( 
.A(n_9166),
.Y(n_10161)
);

AND2x2_ASAP7_75t_L g10162 ( 
.A(n_9536),
.B(n_8224),
.Y(n_10162)
);

AND2x4_ASAP7_75t_L g10163 ( 
.A(n_9735),
.B(n_8742),
.Y(n_10163)
);

INVx2_ASAP7_75t_L g10164 ( 
.A(n_9483),
.Y(n_10164)
);

INVxp67_ASAP7_75t_L g10165 ( 
.A(n_9546),
.Y(n_10165)
);

INVx1_ASAP7_75t_L g10166 ( 
.A(n_9829),
.Y(n_10166)
);

AOI22xp5_ASAP7_75t_L g10167 ( 
.A1(n_9506),
.A2(n_8899),
.B1(n_8851),
.B2(n_9055),
.Y(n_10167)
);

INVx1_ASAP7_75t_L g10168 ( 
.A(n_9842),
.Y(n_10168)
);

INVx2_ASAP7_75t_L g10169 ( 
.A(n_9341),
.Y(n_10169)
);

INVx2_ASAP7_75t_L g10170 ( 
.A(n_9771),
.Y(n_10170)
);

INVx1_ASAP7_75t_L g10171 ( 
.A(n_9771),
.Y(n_10171)
);

AND2x4_ASAP7_75t_SL g10172 ( 
.A(n_9558),
.B(n_8224),
.Y(n_10172)
);

INVx2_ASAP7_75t_L g10173 ( 
.A(n_9771),
.Y(n_10173)
);

AND2x2_ASAP7_75t_L g10174 ( 
.A(n_9558),
.B(n_8224),
.Y(n_10174)
);

INVx1_ASAP7_75t_L g10175 ( 
.A(n_9497),
.Y(n_10175)
);

NOR2xp33_ASAP7_75t_L g10176 ( 
.A(n_9598),
.B(n_5810),
.Y(n_10176)
);

AND2x2_ASAP7_75t_L g10177 ( 
.A(n_9296),
.B(n_8287),
.Y(n_10177)
);

BUFx2_ASAP7_75t_L g10178 ( 
.A(n_9523),
.Y(n_10178)
);

INVx2_ASAP7_75t_L g10179 ( 
.A(n_9298),
.Y(n_10179)
);

NAND2x1_ASAP7_75t_L g10180 ( 
.A(n_9470),
.B(n_9080),
.Y(n_10180)
);

AND2x2_ASAP7_75t_L g10181 ( 
.A(n_9477),
.B(n_9735),
.Y(n_10181)
);

INVx1_ASAP7_75t_L g10182 ( 
.A(n_9501),
.Y(n_10182)
);

NOR2xp33_ASAP7_75t_L g10183 ( 
.A(n_9668),
.B(n_5833),
.Y(n_10183)
);

OR2x2_ASAP7_75t_L g10184 ( 
.A(n_9252),
.B(n_8630),
.Y(n_10184)
);

INVx1_ASAP7_75t_L g10185 ( 
.A(n_9508),
.Y(n_10185)
);

INVx2_ASAP7_75t_SL g10186 ( 
.A(n_9627),
.Y(n_10186)
);

INVx1_ASAP7_75t_L g10187 ( 
.A(n_9557),
.Y(n_10187)
);

INVx3_ASAP7_75t_L g10188 ( 
.A(n_9523),
.Y(n_10188)
);

AND2x2_ASAP7_75t_L g10189 ( 
.A(n_9477),
.B(n_8287),
.Y(n_10189)
);

AND2x2_ASAP7_75t_L g10190 ( 
.A(n_9520),
.B(n_8287),
.Y(n_10190)
);

INVx2_ASAP7_75t_L g10191 ( 
.A(n_9588),
.Y(n_10191)
);

NAND2xp5_ASAP7_75t_L g10192 ( 
.A(n_9554),
.B(n_8631),
.Y(n_10192)
);

INVx1_ASAP7_75t_L g10193 ( 
.A(n_9595),
.Y(n_10193)
);

INVx1_ASAP7_75t_L g10194 ( 
.A(n_9624),
.Y(n_10194)
);

INVx1_ASAP7_75t_L g10195 ( 
.A(n_9646),
.Y(n_10195)
);

INVx2_ASAP7_75t_L g10196 ( 
.A(n_9588),
.Y(n_10196)
);

OR2x2_ASAP7_75t_L g10197 ( 
.A(n_9806),
.B(n_8646),
.Y(n_10197)
);

INVx1_ASAP7_75t_L g10198 ( 
.A(n_9664),
.Y(n_10198)
);

NAND2xp5_ASAP7_75t_L g10199 ( 
.A(n_9210),
.B(n_8650),
.Y(n_10199)
);

INVx1_ASAP7_75t_L g10200 ( 
.A(n_9718),
.Y(n_10200)
);

OR2x2_ASAP7_75t_L g10201 ( 
.A(n_9391),
.B(n_8651),
.Y(n_10201)
);

AND2x2_ASAP7_75t_L g10202 ( 
.A(n_9520),
.B(n_9605),
.Y(n_10202)
);

BUFx3_ASAP7_75t_L g10203 ( 
.A(n_9633),
.Y(n_10203)
);

INVx2_ASAP7_75t_SL g10204 ( 
.A(n_9539),
.Y(n_10204)
);

OR2x2_ASAP7_75t_L g10205 ( 
.A(n_9469),
.B(n_8655),
.Y(n_10205)
);

INVx3_ASAP7_75t_L g10206 ( 
.A(n_9539),
.Y(n_10206)
);

NOR2x1p5_ASAP7_75t_L g10207 ( 
.A(n_9607),
.B(n_8218),
.Y(n_10207)
);

AND2x2_ASAP7_75t_L g10208 ( 
.A(n_9605),
.B(n_8287),
.Y(n_10208)
);

OR2x2_ASAP7_75t_L g10209 ( 
.A(n_9481),
.B(n_8664),
.Y(n_10209)
);

CKINVDCx5p33_ASAP7_75t_R g10210 ( 
.A(n_9649),
.Y(n_10210)
);

INVx2_ASAP7_75t_L g10211 ( 
.A(n_9686),
.Y(n_10211)
);

INVx2_ASAP7_75t_L g10212 ( 
.A(n_9686),
.Y(n_10212)
);

AND2x2_ASAP7_75t_L g10213 ( 
.A(n_9752),
.B(n_8287),
.Y(n_10213)
);

INVx1_ASAP7_75t_L g10214 ( 
.A(n_9685),
.Y(n_10214)
);

BUFx2_ASAP7_75t_L g10215 ( 
.A(n_9608),
.Y(n_10215)
);

INVx1_ASAP7_75t_L g10216 ( 
.A(n_9725),
.Y(n_10216)
);

AND2x2_ASAP7_75t_L g10217 ( 
.A(n_9752),
.B(n_8287),
.Y(n_10217)
);

BUFx2_ASAP7_75t_L g10218 ( 
.A(n_9608),
.Y(n_10218)
);

INVx1_ASAP7_75t_L g10219 ( 
.A(n_9571),
.Y(n_10219)
);

INVx2_ASAP7_75t_L g10220 ( 
.A(n_9814),
.Y(n_10220)
);

AND2x2_ASAP7_75t_L g10221 ( 
.A(n_9814),
.B(n_9027),
.Y(n_10221)
);

INVx1_ASAP7_75t_L g10222 ( 
.A(n_9571),
.Y(n_10222)
);

INVx2_ASAP7_75t_L g10223 ( 
.A(n_9552),
.Y(n_10223)
);

INVx1_ASAP7_75t_L g10224 ( 
.A(n_9571),
.Y(n_10224)
);

AOI22xp33_ASAP7_75t_SL g10225 ( 
.A1(n_9176),
.A2(n_8449),
.B1(n_8456),
.B2(n_8372),
.Y(n_10225)
);

INVx2_ASAP7_75t_L g10226 ( 
.A(n_9709),
.Y(n_10226)
);

NAND2xp5_ASAP7_75t_L g10227 ( 
.A(n_9237),
.B(n_9524),
.Y(n_10227)
);

INVxp67_ASAP7_75t_SL g10228 ( 
.A(n_9315),
.Y(n_10228)
);

AND2x2_ASAP7_75t_L g10229 ( 
.A(n_9415),
.B(n_9027),
.Y(n_10229)
);

NAND2xp5_ASAP7_75t_L g10230 ( 
.A(n_9542),
.B(n_8666),
.Y(n_10230)
);

HB1xp67_ASAP7_75t_L g10231 ( 
.A(n_9340),
.Y(n_10231)
);

INVx3_ASAP7_75t_L g10232 ( 
.A(n_9382),
.Y(n_10232)
);

INVx1_ASAP7_75t_L g10233 ( 
.A(n_9582),
.Y(n_10233)
);

INVx1_ASAP7_75t_L g10234 ( 
.A(n_9582),
.Y(n_10234)
);

INVx2_ASAP7_75t_L g10235 ( 
.A(n_9709),
.Y(n_10235)
);

INVx1_ASAP7_75t_L g10236 ( 
.A(n_9582),
.Y(n_10236)
);

OR2x2_ASAP7_75t_L g10237 ( 
.A(n_9819),
.B(n_8667),
.Y(n_10237)
);

HB1xp67_ASAP7_75t_L g10238 ( 
.A(n_9340),
.Y(n_10238)
);

NAND2xp5_ASAP7_75t_L g10239 ( 
.A(n_9772),
.B(n_8671),
.Y(n_10239)
);

INVx2_ASAP7_75t_L g10240 ( 
.A(n_9791),
.Y(n_10240)
);

INVx2_ASAP7_75t_L g10241 ( 
.A(n_9791),
.Y(n_10241)
);

INVx1_ASAP7_75t_L g10242 ( 
.A(n_9313),
.Y(n_10242)
);

AND2x2_ASAP7_75t_L g10243 ( 
.A(n_9707),
.B(n_9042),
.Y(n_10243)
);

INVx2_ASAP7_75t_L g10244 ( 
.A(n_9827),
.Y(n_10244)
);

INVx2_ASAP7_75t_L g10245 ( 
.A(n_9827),
.Y(n_10245)
);

INVx1_ASAP7_75t_L g10246 ( 
.A(n_9313),
.Y(n_10246)
);

AND2x4_ASAP7_75t_L g10247 ( 
.A(n_9707),
.B(n_8428),
.Y(n_10247)
);

AOI22xp5_ASAP7_75t_L g10248 ( 
.A1(n_9218),
.A2(n_9188),
.B1(n_9199),
.B2(n_9413),
.Y(n_10248)
);

HB1xp67_ASAP7_75t_L g10249 ( 
.A(n_9181),
.Y(n_10249)
);

INVx2_ASAP7_75t_L g10250 ( 
.A(n_9208),
.Y(n_10250)
);

HB1xp67_ASAP7_75t_L g10251 ( 
.A(n_9181),
.Y(n_10251)
);

AND2x4_ASAP7_75t_SL g10252 ( 
.A(n_9707),
.B(n_9773),
.Y(n_10252)
);

INVx1_ASAP7_75t_L g10253 ( 
.A(n_9513),
.Y(n_10253)
);

OR2x2_ASAP7_75t_L g10254 ( 
.A(n_9282),
.B(n_8674),
.Y(n_10254)
);

INVx1_ASAP7_75t_L g10255 ( 
.A(n_9513),
.Y(n_10255)
);

INVx1_ASAP7_75t_L g10256 ( 
.A(n_9513),
.Y(n_10256)
);

INVx2_ASAP7_75t_L g10257 ( 
.A(n_9780),
.Y(n_10257)
);

INVx2_ASAP7_75t_L g10258 ( 
.A(n_9780),
.Y(n_10258)
);

INVx2_ASAP7_75t_L g10259 ( 
.A(n_9187),
.Y(n_10259)
);

HB1xp67_ASAP7_75t_L g10260 ( 
.A(n_9401),
.Y(n_10260)
);

INVx1_ASAP7_75t_L g10261 ( 
.A(n_9359),
.Y(n_10261)
);

INVx2_ASAP7_75t_L g10262 ( 
.A(n_9187),
.Y(n_10262)
);

OR2x2_ASAP7_75t_L g10263 ( 
.A(n_9699),
.B(n_8687),
.Y(n_10263)
);

INVxp67_ASAP7_75t_SL g10264 ( 
.A(n_9266),
.Y(n_10264)
);

AND2x2_ASAP7_75t_L g10265 ( 
.A(n_9773),
.B(n_9042),
.Y(n_10265)
);

AND2x2_ASAP7_75t_L g10266 ( 
.A(n_9773),
.B(n_9072),
.Y(n_10266)
);

AND2x2_ASAP7_75t_L g10267 ( 
.A(n_9837),
.B(n_9072),
.Y(n_10267)
);

AND2x2_ASAP7_75t_L g10268 ( 
.A(n_9612),
.B(n_9096),
.Y(n_10268)
);

CKINVDCx5p33_ASAP7_75t_R g10269 ( 
.A(n_9654),
.Y(n_10269)
);

INVx1_ASAP7_75t_L g10270 ( 
.A(n_9359),
.Y(n_10270)
);

INVx2_ASAP7_75t_L g10271 ( 
.A(n_9187),
.Y(n_10271)
);

INVx1_ASAP7_75t_L g10272 ( 
.A(n_9359),
.Y(n_10272)
);

INVx1_ASAP7_75t_L g10273 ( 
.A(n_9361),
.Y(n_10273)
);

BUFx3_ASAP7_75t_L g10274 ( 
.A(n_9684),
.Y(n_10274)
);

INVx1_ASAP7_75t_L g10275 ( 
.A(n_9361),
.Y(n_10275)
);

HB1xp67_ASAP7_75t_L g10276 ( 
.A(n_9560),
.Y(n_10276)
);

BUFx2_ASAP7_75t_L g10277 ( 
.A(n_9221),
.Y(n_10277)
);

AND2x2_ASAP7_75t_L g10278 ( 
.A(n_9612),
.B(n_9096),
.Y(n_10278)
);

HB1xp67_ASAP7_75t_L g10279 ( 
.A(n_9749),
.Y(n_10279)
);

AND2x2_ASAP7_75t_L g10280 ( 
.A(n_9475),
.B(n_9107),
.Y(n_10280)
);

INVx1_ASAP7_75t_L g10281 ( 
.A(n_9361),
.Y(n_10281)
);

AND2x2_ASAP7_75t_L g10282 ( 
.A(n_9333),
.B(n_9107),
.Y(n_10282)
);

AND2x2_ASAP7_75t_L g10283 ( 
.A(n_9493),
.B(n_9129),
.Y(n_10283)
);

AND2x2_ASAP7_75t_L g10284 ( 
.A(n_9444),
.B(n_9129),
.Y(n_10284)
);

INVx2_ASAP7_75t_L g10285 ( 
.A(n_9832),
.Y(n_10285)
);

INVx3_ASAP7_75t_L g10286 ( 
.A(n_9549),
.Y(n_10286)
);

OR2x2_ASAP7_75t_L g10287 ( 
.A(n_9573),
.B(n_8689),
.Y(n_10287)
);

AND2x2_ASAP7_75t_L g10288 ( 
.A(n_9458),
.B(n_9133),
.Y(n_10288)
);

NOR2xp33_ASAP7_75t_L g10289 ( 
.A(n_9346),
.B(n_5968),
.Y(n_10289)
);

AND2x2_ASAP7_75t_L g10290 ( 
.A(n_9461),
.B(n_9133),
.Y(n_10290)
);

NAND2xp5_ASAP7_75t_L g10291 ( 
.A(n_9239),
.B(n_8691),
.Y(n_10291)
);

INVx1_ASAP7_75t_L g10292 ( 
.A(n_9499),
.Y(n_10292)
);

BUFx2_ASAP7_75t_L g10293 ( 
.A(n_9221),
.Y(n_10293)
);

INVx1_ASAP7_75t_L g10294 ( 
.A(n_9499),
.Y(n_10294)
);

INVxp67_ASAP7_75t_SL g10295 ( 
.A(n_9465),
.Y(n_10295)
);

NAND2xp5_ASAP7_75t_L g10296 ( 
.A(n_9789),
.B(n_8694),
.Y(n_10296)
);

INVx2_ASAP7_75t_L g10297 ( 
.A(n_9832),
.Y(n_10297)
);

AOI22xp33_ASAP7_75t_SL g10298 ( 
.A1(n_9526),
.A2(n_8449),
.B1(n_8456),
.B2(n_8372),
.Y(n_10298)
);

INVx2_ASAP7_75t_L g10299 ( 
.A(n_9260),
.Y(n_10299)
);

INVxp67_ASAP7_75t_SL g10300 ( 
.A(n_9465),
.Y(n_10300)
);

AND2x4_ASAP7_75t_L g10301 ( 
.A(n_9472),
.B(n_8428),
.Y(n_10301)
);

INVx1_ASAP7_75t_L g10302 ( 
.A(n_9222),
.Y(n_10302)
);

AOI22xp33_ASAP7_75t_L g10303 ( 
.A1(n_9251),
.A2(n_8773),
.B1(n_8779),
.B2(n_8765),
.Y(n_10303)
);

AND2x2_ASAP7_75t_L g10304 ( 
.A(n_9495),
.B(n_9142),
.Y(n_10304)
);

INVx1_ASAP7_75t_L g10305 ( 
.A(n_9222),
.Y(n_10305)
);

INVx1_ASAP7_75t_L g10306 ( 
.A(n_9222),
.Y(n_10306)
);

INVx1_ASAP7_75t_L g10307 ( 
.A(n_9258),
.Y(n_10307)
);

INVx2_ASAP7_75t_L g10308 ( 
.A(n_9798),
.Y(n_10308)
);

NAND2xp5_ASAP7_75t_L g10309 ( 
.A(n_9278),
.B(n_8695),
.Y(n_10309)
);

AND2x4_ASAP7_75t_L g10310 ( 
.A(n_9833),
.B(n_8428),
.Y(n_10310)
);

INVx2_ASAP7_75t_L g10311 ( 
.A(n_9620),
.Y(n_10311)
);

INVx1_ASAP7_75t_L g10312 ( 
.A(n_9258),
.Y(n_10312)
);

NAND2xp5_ASAP7_75t_L g10313 ( 
.A(n_9254),
.B(n_8697),
.Y(n_10313)
);

BUFx2_ASAP7_75t_SL g10314 ( 
.A(n_9833),
.Y(n_10314)
);

HB1xp67_ASAP7_75t_L g10315 ( 
.A(n_9400),
.Y(n_10315)
);

AOI222xp33_ASAP7_75t_L g10316 ( 
.A1(n_9405),
.A2(n_8545),
.B1(n_8542),
.B2(n_8548),
.C1(n_8543),
.C2(n_8539),
.Y(n_10316)
);

AND2x2_ASAP7_75t_L g10317 ( 
.A(n_9509),
.B(n_9142),
.Y(n_10317)
);

INVx1_ASAP7_75t_L g10318 ( 
.A(n_9258),
.Y(n_10318)
);

INVx2_ASAP7_75t_L g10319 ( 
.A(n_9620),
.Y(n_10319)
);

BUFx2_ASAP7_75t_L g10320 ( 
.A(n_9429),
.Y(n_10320)
);

AND2x2_ASAP7_75t_L g10321 ( 
.A(n_9437),
.B(n_9151),
.Y(n_10321)
);

INVx4_ASAP7_75t_L g10322 ( 
.A(n_9754),
.Y(n_10322)
);

INVx2_ASAP7_75t_L g10323 ( 
.A(n_9648),
.Y(n_10323)
);

AND2x2_ASAP7_75t_L g10324 ( 
.A(n_9544),
.B(n_9151),
.Y(n_10324)
);

INVx2_ASAP7_75t_L g10325 ( 
.A(n_9648),
.Y(n_10325)
);

INVx1_ASAP7_75t_L g10326 ( 
.A(n_9291),
.Y(n_10326)
);

INVxp67_ASAP7_75t_SL g10327 ( 
.A(n_9358),
.Y(n_10327)
);

AND2x2_ASAP7_75t_L g10328 ( 
.A(n_9422),
.B(n_9157),
.Y(n_10328)
);

INVx2_ASAP7_75t_L g10329 ( 
.A(n_9488),
.Y(n_10329)
);

BUFx3_ASAP7_75t_L g10330 ( 
.A(n_9722),
.Y(n_10330)
);

AND2x2_ASAP7_75t_L g10331 ( 
.A(n_9377),
.B(n_9157),
.Y(n_10331)
);

INVx2_ASAP7_75t_L g10332 ( 
.A(n_9384),
.Y(n_10332)
);

INVx2_ASAP7_75t_L g10333 ( 
.A(n_9384),
.Y(n_10333)
);

INVx1_ASAP7_75t_L g10334 ( 
.A(n_9291),
.Y(n_10334)
);

INVx1_ASAP7_75t_L g10335 ( 
.A(n_9291),
.Y(n_10335)
);

INVx3_ASAP7_75t_L g10336 ( 
.A(n_9816),
.Y(n_10336)
);

INVx1_ASAP7_75t_L g10337 ( 
.A(n_9338),
.Y(n_10337)
);

NAND2xp5_ASAP7_75t_L g10338 ( 
.A(n_9727),
.B(n_8700),
.Y(n_10338)
);

INVx4_ASAP7_75t_L g10339 ( 
.A(n_9770),
.Y(n_10339)
);

AND2x2_ASAP7_75t_L g10340 ( 
.A(n_9374),
.B(n_9159),
.Y(n_10340)
);

AND2x2_ASAP7_75t_L g10341 ( 
.A(n_9550),
.B(n_9159),
.Y(n_10341)
);

INVx1_ASAP7_75t_L g10342 ( 
.A(n_9343),
.Y(n_10342)
);

NAND2xp5_ASAP7_75t_L g10343 ( 
.A(n_9759),
.B(n_8703),
.Y(n_10343)
);

OR2x2_ASAP7_75t_L g10344 ( 
.A(n_9354),
.B(n_8710),
.Y(n_10344)
);

INVx3_ASAP7_75t_L g10345 ( 
.A(n_9756),
.Y(n_10345)
);

AO31x2_ASAP7_75t_L g10346 ( 
.A1(n_9276),
.A2(n_8400),
.A3(n_8410),
.B(n_8385),
.Y(n_10346)
);

NAND2xp5_ASAP7_75t_L g10347 ( 
.A(n_9792),
.B(n_8711),
.Y(n_10347)
);

NAND2xp5_ASAP7_75t_L g10348 ( 
.A(n_9244),
.B(n_8715),
.Y(n_10348)
);

INVx2_ASAP7_75t_L g10349 ( 
.A(n_9294),
.Y(n_10349)
);

AND2x2_ASAP7_75t_L g10350 ( 
.A(n_9760),
.B(n_9160),
.Y(n_10350)
);

INVx2_ASAP7_75t_L g10351 ( 
.A(n_9286),
.Y(n_10351)
);

INVx1_ASAP7_75t_L g10352 ( 
.A(n_9442),
.Y(n_10352)
);

BUFx3_ASAP7_75t_L g10353 ( 
.A(n_9722),
.Y(n_10353)
);

AND2x2_ASAP7_75t_L g10354 ( 
.A(n_9716),
.B(n_9160),
.Y(n_10354)
);

NAND2xp5_ASAP7_75t_L g10355 ( 
.A(n_9268),
.B(n_8725),
.Y(n_10355)
);

AND2x2_ASAP7_75t_L g10356 ( 
.A(n_9460),
.B(n_7235),
.Y(n_10356)
);

INVx2_ASAP7_75t_L g10357 ( 
.A(n_9731),
.Y(n_10357)
);

AND2x4_ASAP7_75t_L g10358 ( 
.A(n_9835),
.B(n_8484),
.Y(n_10358)
);

NAND2xp5_ASAP7_75t_L g10359 ( 
.A(n_9317),
.B(n_8727),
.Y(n_10359)
);

NOR2xp33_ASAP7_75t_L g10360 ( 
.A(n_9575),
.B(n_6050),
.Y(n_10360)
);

INVx2_ASAP7_75t_L g10361 ( 
.A(n_9666),
.Y(n_10361)
);

INVx2_ASAP7_75t_L g10362 ( 
.A(n_9304),
.Y(n_10362)
);

INVx2_ASAP7_75t_L g10363 ( 
.A(n_9799),
.Y(n_10363)
);

INVx2_ASAP7_75t_L g10364 ( 
.A(n_9803),
.Y(n_10364)
);

INVx1_ASAP7_75t_L g10365 ( 
.A(n_9500),
.Y(n_10365)
);

INVx2_ASAP7_75t_L g10366 ( 
.A(n_9594),
.Y(n_10366)
);

AND2x2_ASAP7_75t_L g10367 ( 
.A(n_9599),
.B(n_7235),
.Y(n_10367)
);

AND2x4_ASAP7_75t_SL g10368 ( 
.A(n_9745),
.B(n_6352),
.Y(n_10368)
);

HB1xp67_ASAP7_75t_L g10369 ( 
.A(n_9369),
.Y(n_10369)
);

INVxp67_ASAP7_75t_SL g10370 ( 
.A(n_9412),
.Y(n_10370)
);

INVx2_ASAP7_75t_L g10371 ( 
.A(n_9585),
.Y(n_10371)
);

INVx1_ASAP7_75t_L g10372 ( 
.A(n_9541),
.Y(n_10372)
);

INVx1_ASAP7_75t_L g10373 ( 
.A(n_9711),
.Y(n_10373)
);

INVx1_ASAP7_75t_L g10374 ( 
.A(n_9765),
.Y(n_10374)
);

INVx1_ASAP7_75t_L g10375 ( 
.A(n_9777),
.Y(n_10375)
);

INVx3_ASAP7_75t_L g10376 ( 
.A(n_9758),
.Y(n_10376)
);

INVx1_ASAP7_75t_L g10377 ( 
.A(n_9410),
.Y(n_10377)
);

NAND2xp5_ASAP7_75t_L g10378 ( 
.A(n_9399),
.B(n_8737),
.Y(n_10378)
);

AND2x2_ASAP7_75t_L g10379 ( 
.A(n_9609),
.B(n_7250),
.Y(n_10379)
);

BUFx2_ASAP7_75t_L g10380 ( 
.A(n_9593),
.Y(n_10380)
);

NOR2xp67_ASAP7_75t_L g10381 ( 
.A(n_9219),
.B(n_8254),
.Y(n_10381)
);

BUFx6f_ASAP7_75t_L g10382 ( 
.A(n_9782),
.Y(n_10382)
);

BUFx2_ASAP7_75t_L g10383 ( 
.A(n_9644),
.Y(n_10383)
);

NAND2x1_ASAP7_75t_L g10384 ( 
.A(n_9468),
.B(n_9080),
.Y(n_10384)
);

AND2x2_ASAP7_75t_L g10385 ( 
.A(n_9486),
.B(n_7250),
.Y(n_10385)
);

BUFx2_ASAP7_75t_L g10386 ( 
.A(n_9644),
.Y(n_10386)
);

AOI222xp33_ASAP7_75t_L g10387 ( 
.A1(n_9307),
.A2(n_8548),
.B1(n_8543),
.B2(n_8554),
.C1(n_8545),
.C2(n_8539),
.Y(n_10387)
);

HB1xp67_ASAP7_75t_L g10388 ( 
.A(n_9548),
.Y(n_10388)
);

AND2x2_ASAP7_75t_L g10389 ( 
.A(n_9619),
.B(n_7250),
.Y(n_10389)
);

NAND2xp5_ASAP7_75t_L g10390 ( 
.A(n_9297),
.B(n_8755),
.Y(n_10390)
);

INVxp67_ASAP7_75t_SL g10391 ( 
.A(n_9326),
.Y(n_10391)
);

AND2x2_ASAP7_75t_L g10392 ( 
.A(n_9625),
.B(n_7284),
.Y(n_10392)
);

AND2x4_ASAP7_75t_L g10393 ( 
.A(n_9745),
.B(n_8484),
.Y(n_10393)
);

INVx2_ASAP7_75t_L g10394 ( 
.A(n_9784),
.Y(n_10394)
);

INVxp67_ASAP7_75t_SL g10395 ( 
.A(n_9414),
.Y(n_10395)
);

AND2x2_ASAP7_75t_L g10396 ( 
.A(n_9630),
.B(n_7284),
.Y(n_10396)
);

INVx4_ASAP7_75t_L g10397 ( 
.A(n_9826),
.Y(n_10397)
);

AND2x2_ASAP7_75t_L g10398 ( 
.A(n_9637),
.B(n_7284),
.Y(n_10398)
);

INVx1_ASAP7_75t_L g10399 ( 
.A(n_9407),
.Y(n_10399)
);

INVx1_ASAP7_75t_L g10400 ( 
.A(n_9299),
.Y(n_10400)
);

AO21x2_ASAP7_75t_L g10401 ( 
.A1(n_9533),
.A2(n_8410),
.B(n_8400),
.Y(n_10401)
);

AND2x2_ASAP7_75t_L g10402 ( 
.A(n_9720),
.B(n_8231),
.Y(n_10402)
);

INVx1_ASAP7_75t_SL g10403 ( 
.A(n_9694),
.Y(n_10403)
);

INVx1_ASAP7_75t_L g10404 ( 
.A(n_9396),
.Y(n_10404)
);

HB1xp67_ASAP7_75t_L g10405 ( 
.A(n_9564),
.Y(n_10405)
);

INVxp67_ASAP7_75t_SL g10406 ( 
.A(n_9418),
.Y(n_10406)
);

INVx2_ASAP7_75t_L g10407 ( 
.A(n_9249),
.Y(n_10407)
);

INVx3_ASAP7_75t_L g10408 ( 
.A(n_9397),
.Y(n_10408)
);

BUFx2_ASAP7_75t_L g10409 ( 
.A(n_9323),
.Y(n_10409)
);

AND2x4_ASAP7_75t_L g10410 ( 
.A(n_9675),
.B(n_8484),
.Y(n_10410)
);

INVx2_ASAP7_75t_L g10411 ( 
.A(n_9562),
.Y(n_10411)
);

BUFx3_ASAP7_75t_L g10412 ( 
.A(n_9696),
.Y(n_10412)
);

INVx1_ASAP7_75t_L g10413 ( 
.A(n_9402),
.Y(n_10413)
);

INVx2_ASAP7_75t_L g10414 ( 
.A(n_9566),
.Y(n_10414)
);

NAND2xp5_ASAP7_75t_L g10415 ( 
.A(n_9748),
.B(n_8762),
.Y(n_10415)
);

AND2x2_ASAP7_75t_L g10416 ( 
.A(n_9726),
.B(n_8231),
.Y(n_10416)
);

OR2x2_ASAP7_75t_L g10417 ( 
.A(n_9569),
.B(n_8763),
.Y(n_10417)
);

HB1xp67_ASAP7_75t_L g10418 ( 
.A(n_9504),
.Y(n_10418)
);

BUFx3_ASAP7_75t_L g10419 ( 
.A(n_9696),
.Y(n_10419)
);

INVx2_ASAP7_75t_L g10420 ( 
.A(n_9200),
.Y(n_10420)
);

INVx2_ASAP7_75t_L g10421 ( 
.A(n_9578),
.Y(n_10421)
);

INVx1_ASAP7_75t_L g10422 ( 
.A(n_9671),
.Y(n_10422)
);

INVx2_ASAP7_75t_L g10423 ( 
.A(n_9578),
.Y(n_10423)
);

BUFx3_ASAP7_75t_L g10424 ( 
.A(n_9682),
.Y(n_10424)
);

INVx2_ASAP7_75t_L g10425 ( 
.A(n_9462),
.Y(n_10425)
);

INVx1_ASAP7_75t_L g10426 ( 
.A(n_9319),
.Y(n_10426)
);

AND2x4_ASAP7_75t_L g10427 ( 
.A(n_9681),
.B(n_8508),
.Y(n_10427)
);

INVx1_ASAP7_75t_L g10428 ( 
.A(n_9371),
.Y(n_10428)
);

AND2x2_ASAP7_75t_L g10429 ( 
.A(n_9750),
.B(n_9767),
.Y(n_10429)
);

INVx2_ASAP7_75t_L g10430 ( 
.A(n_9387),
.Y(n_10430)
);

NAND2xp5_ASAP7_75t_L g10431 ( 
.A(n_9232),
.B(n_8766),
.Y(n_10431)
);

INVx1_ASAP7_75t_L g10432 ( 
.A(n_9394),
.Y(n_10432)
);

INVx1_ASAP7_75t_L g10433 ( 
.A(n_9744),
.Y(n_10433)
);

INVx1_ASAP7_75t_L g10434 ( 
.A(n_9512),
.Y(n_10434)
);

INVx1_ASAP7_75t_L g10435 ( 
.A(n_9274),
.Y(n_10435)
);

AND2x2_ASAP7_75t_L g10436 ( 
.A(n_9769),
.B(n_8249),
.Y(n_10436)
);

INVx1_ASAP7_75t_L g10437 ( 
.A(n_9423),
.Y(n_10437)
);

OR2x2_ASAP7_75t_L g10438 ( 
.A(n_9746),
.B(n_8768),
.Y(n_10438)
);

INVx1_ASAP7_75t_L g10439 ( 
.A(n_9449),
.Y(n_10439)
);

AOI22xp33_ASAP7_75t_L g10440 ( 
.A1(n_9413),
.A2(n_8797),
.B1(n_8805),
.B2(n_8779),
.Y(n_10440)
);

NOR2x1p5_ASAP7_75t_L g10441 ( 
.A(n_9647),
.B(n_8218),
.Y(n_10441)
);

INVx2_ASAP7_75t_L g10442 ( 
.A(n_9240),
.Y(n_10442)
);

BUFx2_ASAP7_75t_L g10443 ( 
.A(n_9433),
.Y(n_10443)
);

INVx1_ASAP7_75t_L g10444 ( 
.A(n_9455),
.Y(n_10444)
);

AND2x4_ASAP7_75t_L g10445 ( 
.A(n_9473),
.B(n_8508),
.Y(n_10445)
);

AND2x2_ASAP7_75t_L g10446 ( 
.A(n_9775),
.B(n_8249),
.Y(n_10446)
);

OR2x2_ASAP7_75t_L g10447 ( 
.A(n_9355),
.B(n_8770),
.Y(n_10447)
);

AND2x2_ASAP7_75t_L g10448 ( 
.A(n_9788),
.B(n_8349),
.Y(n_10448)
);

AND2x2_ASAP7_75t_L g10449 ( 
.A(n_9794),
.B(n_8349),
.Y(n_10449)
);

AND2x2_ASAP7_75t_L g10450 ( 
.A(n_9808),
.B(n_8558),
.Y(n_10450)
);

AND2x4_ASAP7_75t_L g10451 ( 
.A(n_9478),
.B(n_8508),
.Y(n_10451)
);

BUFx2_ASAP7_75t_L g10452 ( 
.A(n_9790),
.Y(n_10452)
);

INVx1_ASAP7_75t_L g10453 ( 
.A(n_9269),
.Y(n_10453)
);

NAND2xp5_ASAP7_75t_L g10454 ( 
.A(n_9724),
.B(n_8775),
.Y(n_10454)
);

AND2x4_ASAP7_75t_L g10455 ( 
.A(n_9480),
.B(n_8570),
.Y(n_10455)
);

INVx2_ASAP7_75t_L g10456 ( 
.A(n_9762),
.Y(n_10456)
);

AND2x2_ASAP7_75t_L g10457 ( 
.A(n_9818),
.B(n_8558),
.Y(n_10457)
);

BUFx3_ASAP7_75t_L g10458 ( 
.A(n_9308),
.Y(n_10458)
);

INVx1_ASAP7_75t_L g10459 ( 
.A(n_9378),
.Y(n_10459)
);

INVx2_ASAP7_75t_L g10460 ( 
.A(n_9807),
.Y(n_10460)
);

AND2x2_ASAP7_75t_L g10461 ( 
.A(n_9820),
.B(n_8795),
.Y(n_10461)
);

INVx2_ASAP7_75t_L g10462 ( 
.A(n_9812),
.Y(n_10462)
);

AND2x2_ASAP7_75t_L g10463 ( 
.A(n_9831),
.B(n_8795),
.Y(n_10463)
);

INVx2_ASAP7_75t_L g10464 ( 
.A(n_9804),
.Y(n_10464)
);

NOR2xp33_ASAP7_75t_L g10465 ( 
.A(n_9196),
.B(n_6050),
.Y(n_10465)
);

NAND2xp5_ASAP7_75t_L g10466 ( 
.A(n_9476),
.B(n_8776),
.Y(n_10466)
);

INVx2_ASAP7_75t_L g10467 ( 
.A(n_9804),
.Y(n_10467)
);

BUFx2_ASAP7_75t_L g10468 ( 
.A(n_9790),
.Y(n_10468)
);

AND2x2_ASAP7_75t_L g10469 ( 
.A(n_9841),
.B(n_8877),
.Y(n_10469)
);

OR2x2_ASAP7_75t_L g10470 ( 
.A(n_9236),
.B(n_8780),
.Y(n_10470)
);

NAND3xp33_ASAP7_75t_L g10471 ( 
.A(n_9611),
.B(n_8662),
.C(n_8620),
.Y(n_10471)
);

HB1xp67_ASAP7_75t_L g10472 ( 
.A(n_9487),
.Y(n_10472)
);

AND2x4_ASAP7_75t_L g10473 ( 
.A(n_9485),
.B(n_8570),
.Y(n_10473)
);

AND2x2_ASAP7_75t_L g10474 ( 
.A(n_9738),
.B(n_8877),
.Y(n_10474)
);

INVx2_ASAP7_75t_L g10475 ( 
.A(n_9408),
.Y(n_10475)
);

INVxp67_ASAP7_75t_L g10476 ( 
.A(n_9311),
.Y(n_10476)
);

INVx1_ASAP7_75t_L g10477 ( 
.A(n_9420),
.Y(n_10477)
);

INVx1_ASAP7_75t_L g10478 ( 
.A(n_9427),
.Y(n_10478)
);

AND2x2_ASAP7_75t_L g10479 ( 
.A(n_9683),
.B(n_8877),
.Y(n_10479)
);

AND2x4_ASAP7_75t_L g10480 ( 
.A(n_9491),
.B(n_8570),
.Y(n_10480)
);

INVx2_ASAP7_75t_L g10481 ( 
.A(n_9779),
.Y(n_10481)
);

INVxp67_ASAP7_75t_L g10482 ( 
.A(n_9267),
.Y(n_10482)
);

BUFx2_ASAP7_75t_L g10483 ( 
.A(n_9305),
.Y(n_10483)
);

INVxp67_ASAP7_75t_L g10484 ( 
.A(n_9479),
.Y(n_10484)
);

AOI22xp5_ASAP7_75t_L g10485 ( 
.A1(n_10295),
.A2(n_9418),
.B1(n_9173),
.B2(n_9214),
.Y(n_10485)
);

AOI22xp33_ASAP7_75t_SL g10486 ( 
.A1(n_10408),
.A2(n_9496),
.B1(n_9632),
.B2(n_9613),
.Y(n_10486)
);

NAND2xp5_ASAP7_75t_L g10487 ( 
.A(n_9883),
.B(n_9265),
.Y(n_10487)
);

INVx1_ASAP7_75t_L g10488 ( 
.A(n_9921),
.Y(n_10488)
);

OR2x2_ASAP7_75t_L g10489 ( 
.A(n_9949),
.B(n_9604),
.Y(n_10489)
);

INVx2_ASAP7_75t_L g10490 ( 
.A(n_9951),
.Y(n_10490)
);

AND2x2_ASAP7_75t_L g10491 ( 
.A(n_9857),
.B(n_9662),
.Y(n_10491)
);

INVx1_ASAP7_75t_L g10492 ( 
.A(n_9921),
.Y(n_10492)
);

INVx1_ASAP7_75t_L g10493 ( 
.A(n_10231),
.Y(n_10493)
);

INVx1_ASAP7_75t_L g10494 ( 
.A(n_10231),
.Y(n_10494)
);

INVx5_ASAP7_75t_L g10495 ( 
.A(n_9907),
.Y(n_10495)
);

AND2x4_ASAP7_75t_L g10496 ( 
.A(n_9892),
.B(n_9502),
.Y(n_10496)
);

OR2x2_ASAP7_75t_L g10497 ( 
.A(n_10047),
.B(n_8782),
.Y(n_10497)
);

INVx2_ASAP7_75t_L g10498 ( 
.A(n_9951),
.Y(n_10498)
);

INVx1_ASAP7_75t_L g10499 ( 
.A(n_10238),
.Y(n_10499)
);

OR2x2_ASAP7_75t_L g10500 ( 
.A(n_9851),
.B(n_8784),
.Y(n_10500)
);

AND2x2_ASAP7_75t_L g10501 ( 
.A(n_9861),
.B(n_9662),
.Y(n_10501)
);

INVx1_ASAP7_75t_L g10502 ( 
.A(n_10238),
.Y(n_10502)
);

INVx1_ASAP7_75t_L g10503 ( 
.A(n_10249),
.Y(n_10503)
);

AND2x2_ASAP7_75t_L g10504 ( 
.A(n_9922),
.B(n_9603),
.Y(n_10504)
);

NOR2xp67_ASAP7_75t_L g10505 ( 
.A(n_10002),
.B(n_9795),
.Y(n_10505)
);

INVx2_ASAP7_75t_L g10506 ( 
.A(n_9951),
.Y(n_10506)
);

OR2x2_ASAP7_75t_L g10507 ( 
.A(n_9855),
.B(n_8786),
.Y(n_10507)
);

HB1xp67_ASAP7_75t_L g10508 ( 
.A(n_9997),
.Y(n_10508)
);

NAND2xp5_ASAP7_75t_L g10509 ( 
.A(n_9883),
.B(n_9261),
.Y(n_10509)
);

AOI22xp33_ASAP7_75t_L g10510 ( 
.A1(n_10037),
.A2(n_9597),
.B1(n_9471),
.B2(n_9314),
.Y(n_10510)
);

INVx1_ASAP7_75t_L g10511 ( 
.A(n_10249),
.Y(n_10511)
);

INVx1_ASAP7_75t_L g10512 ( 
.A(n_10251),
.Y(n_10512)
);

AND2x2_ASAP7_75t_L g10513 ( 
.A(n_9922),
.B(n_9482),
.Y(n_10513)
);

OR2x2_ASAP7_75t_L g10514 ( 
.A(n_9967),
.B(n_8787),
.Y(n_10514)
);

INVx1_ASAP7_75t_L g10515 ( 
.A(n_10251),
.Y(n_10515)
);

INVx1_ASAP7_75t_L g10516 ( 
.A(n_10039),
.Y(n_10516)
);

INVxp67_ASAP7_75t_L g10517 ( 
.A(n_10183),
.Y(n_10517)
);

NAND2xp5_ASAP7_75t_L g10518 ( 
.A(n_10117),
.B(n_9614),
.Y(n_10518)
);

AND2x2_ASAP7_75t_L g10519 ( 
.A(n_9900),
.B(n_8902),
.Y(n_10519)
);

INVx1_ASAP7_75t_L g10520 ( 
.A(n_10039),
.Y(n_10520)
);

NAND2xp5_ASAP7_75t_L g10521 ( 
.A(n_10117),
.B(n_9753),
.Y(n_10521)
);

AND2x2_ASAP7_75t_L g10522 ( 
.A(n_9872),
.B(n_8906),
.Y(n_10522)
);

INVx1_ASAP7_75t_L g10523 ( 
.A(n_10054),
.Y(n_10523)
);

INVx1_ASAP7_75t_L g10524 ( 
.A(n_10054),
.Y(n_10524)
);

HB1xp67_ASAP7_75t_L g10525 ( 
.A(n_10018),
.Y(n_10525)
);

INVx1_ASAP7_75t_L g10526 ( 
.A(n_10107),
.Y(n_10526)
);

NOR3xp33_ASAP7_75t_L g10527 ( 
.A(n_10132),
.B(n_10476),
.C(n_9945),
.Y(n_10527)
);

OR2x2_ASAP7_75t_L g10528 ( 
.A(n_9977),
.B(n_8788),
.Y(n_10528)
);

AND2x2_ASAP7_75t_L g10529 ( 
.A(n_9872),
.B(n_8906),
.Y(n_10529)
);

BUFx3_ASAP7_75t_L g10530 ( 
.A(n_9906),
.Y(n_10530)
);

HB1xp67_ASAP7_75t_L g10531 ( 
.A(n_10130),
.Y(n_10531)
);

INVxp67_ASAP7_75t_SL g10532 ( 
.A(n_9945),
.Y(n_10532)
);

AOI22xp33_ASAP7_75t_L g10533 ( 
.A1(n_10037),
.A2(n_10300),
.B1(n_10295),
.B2(n_10418),
.Y(n_10533)
);

INVxp67_ASAP7_75t_SL g10534 ( 
.A(n_9876),
.Y(n_10534)
);

AND2x4_ASAP7_75t_SL g10535 ( 
.A(n_9907),
.B(n_6179),
.Y(n_10535)
);

NAND2xp5_ASAP7_75t_L g10536 ( 
.A(n_10143),
.B(n_9306),
.Y(n_10536)
);

AND2x4_ASAP7_75t_L g10537 ( 
.A(n_9892),
.B(n_9505),
.Y(n_10537)
);

INVxp67_ASAP7_75t_SL g10538 ( 
.A(n_9876),
.Y(n_10538)
);

INVx1_ASAP7_75t_L g10539 ( 
.A(n_9867),
.Y(n_10539)
);

AND2x2_ASAP7_75t_L g10540 ( 
.A(n_10001),
.B(n_8914),
.Y(n_10540)
);

INVx1_ASAP7_75t_L g10541 ( 
.A(n_9867),
.Y(n_10541)
);

NAND2xp5_ASAP7_75t_L g10542 ( 
.A(n_10143),
.B(n_9761),
.Y(n_10542)
);

HB1xp67_ASAP7_75t_L g10543 ( 
.A(n_10136),
.Y(n_10543)
);

AOI22xp33_ASAP7_75t_L g10544 ( 
.A1(n_10300),
.A2(n_9503),
.B1(n_9264),
.B2(n_9257),
.Y(n_10544)
);

INVx2_ASAP7_75t_L g10545 ( 
.A(n_10001),
.Y(n_10545)
);

INVx4_ASAP7_75t_R g10546 ( 
.A(n_9885),
.Y(n_10546)
);

INVx2_ASAP7_75t_L g10547 ( 
.A(n_9978),
.Y(n_10547)
);

INVx1_ASAP7_75t_SL g10548 ( 
.A(n_9906),
.Y(n_10548)
);

NOR2xp33_ASAP7_75t_L g10549 ( 
.A(n_9885),
.B(n_6069),
.Y(n_10549)
);

NAND2xp5_ASAP7_75t_L g10550 ( 
.A(n_9915),
.B(n_9279),
.Y(n_10550)
);

AND2x2_ASAP7_75t_L g10551 ( 
.A(n_9978),
.B(n_9881),
.Y(n_10551)
);

AND2x2_ASAP7_75t_L g10552 ( 
.A(n_9881),
.B(n_8914),
.Y(n_10552)
);

NAND2xp67_ASAP7_75t_L g10553 ( 
.A(n_9962),
.B(n_9576),
.Y(n_10553)
);

NOR2xp33_ASAP7_75t_L g10554 ( 
.A(n_9873),
.B(n_6069),
.Y(n_10554)
);

AND2x4_ASAP7_75t_L g10555 ( 
.A(n_9929),
.B(n_9511),
.Y(n_10555)
);

INVx1_ASAP7_75t_L g10556 ( 
.A(n_9896),
.Y(n_10556)
);

OR2x2_ASAP7_75t_L g10557 ( 
.A(n_9970),
.B(n_8789),
.Y(n_10557)
);

AOI22xp33_ASAP7_75t_L g10558 ( 
.A1(n_10418),
.A2(n_9174),
.B1(n_9356),
.B2(n_9227),
.Y(n_10558)
);

INVx1_ASAP7_75t_L g10559 ( 
.A(n_9896),
.Y(n_10559)
);

INVx2_ASAP7_75t_L g10560 ( 
.A(n_10060),
.Y(n_10560)
);

INVx1_ASAP7_75t_L g10561 ( 
.A(n_9898),
.Y(n_10561)
);

HB1xp67_ASAP7_75t_L g10562 ( 
.A(n_10136),
.Y(n_10562)
);

INVxp67_ASAP7_75t_SL g10563 ( 
.A(n_9905),
.Y(n_10563)
);

AND2x2_ASAP7_75t_L g10564 ( 
.A(n_9905),
.B(n_9565),
.Y(n_10564)
);

BUFx2_ASAP7_75t_SL g10565 ( 
.A(n_10161),
.Y(n_10565)
);

INVx1_ASAP7_75t_L g10566 ( 
.A(n_9898),
.Y(n_10566)
);

AND2x2_ASAP7_75t_L g10567 ( 
.A(n_9931),
.B(n_9574),
.Y(n_10567)
);

AND2x2_ASAP7_75t_L g10568 ( 
.A(n_10011),
.B(n_9514),
.Y(n_10568)
);

INVx5_ASAP7_75t_L g10569 ( 
.A(n_10161),
.Y(n_10569)
);

NAND2xp5_ASAP7_75t_L g10570 ( 
.A(n_9847),
.B(n_9801),
.Y(n_10570)
);

INVx2_ASAP7_75t_L g10571 ( 
.A(n_10060),
.Y(n_10571)
);

INVx2_ASAP7_75t_L g10572 ( 
.A(n_10060),
.Y(n_10572)
);

AND2x2_ASAP7_75t_L g10573 ( 
.A(n_10011),
.B(n_9517),
.Y(n_10573)
);

NAND2xp5_ASAP7_75t_L g10574 ( 
.A(n_10482),
.B(n_9817),
.Y(n_10574)
);

NAND2xp5_ASAP7_75t_L g10575 ( 
.A(n_10482),
.B(n_9459),
.Y(n_10575)
);

AND2x2_ASAP7_75t_L g10576 ( 
.A(n_9854),
.B(n_9528),
.Y(n_10576)
);

AOI22xp33_ASAP7_75t_L g10577 ( 
.A1(n_10388),
.A2(n_9778),
.B1(n_9797),
.B2(n_9739),
.Y(n_10577)
);

INVx2_ASAP7_75t_L g10578 ( 
.A(n_10147),
.Y(n_10578)
);

INVx1_ASAP7_75t_L g10579 ( 
.A(n_9952),
.Y(n_10579)
);

HB1xp67_ASAP7_75t_L g10580 ( 
.A(n_10472),
.Y(n_10580)
);

AND2x4_ASAP7_75t_L g10581 ( 
.A(n_9929),
.B(n_9530),
.Y(n_10581)
);

AO22x1_ASAP7_75t_L g10582 ( 
.A1(n_10391),
.A2(n_10370),
.B1(n_10406),
.B2(n_10472),
.Y(n_10582)
);

INVx1_ASAP7_75t_SL g10583 ( 
.A(n_10089),
.Y(n_10583)
);

NAND2xp5_ASAP7_75t_L g10584 ( 
.A(n_10165),
.B(n_8790),
.Y(n_10584)
);

AND2x2_ASAP7_75t_L g10585 ( 
.A(n_9864),
.B(n_9532),
.Y(n_10585)
);

NOR2x1_ASAP7_75t_SL g10586 ( 
.A(n_10065),
.B(n_5936),
.Y(n_10586)
);

INVx1_ASAP7_75t_L g10587 ( 
.A(n_9952),
.Y(n_10587)
);

INVx2_ASAP7_75t_SL g10588 ( 
.A(n_10065),
.Y(n_10588)
);

OAI22x1_ASAP7_75t_L g10589 ( 
.A1(n_10248),
.A2(n_6169),
.B1(n_6171),
.B2(n_6152),
.Y(n_10589)
);

INVx1_ASAP7_75t_L g10590 ( 
.A(n_9958),
.Y(n_10590)
);

AND2x2_ASAP7_75t_L g10591 ( 
.A(n_9930),
.B(n_9545),
.Y(n_10591)
);

INVx2_ASAP7_75t_L g10592 ( 
.A(n_10147),
.Y(n_10592)
);

INVx1_ASAP7_75t_L g10593 ( 
.A(n_9958),
.Y(n_10593)
);

INVx2_ASAP7_75t_L g10594 ( 
.A(n_10147),
.Y(n_10594)
);

INVx2_ASAP7_75t_L g10595 ( 
.A(n_10004),
.Y(n_10595)
);

HB1xp67_ASAP7_75t_L g10596 ( 
.A(n_9893),
.Y(n_10596)
);

NAND2x1p5_ASAP7_75t_L g10597 ( 
.A(n_9993),
.B(n_9046),
.Y(n_10597)
);

INVx1_ASAP7_75t_L g10598 ( 
.A(n_9964),
.Y(n_10598)
);

NAND2xp5_ASAP7_75t_L g10599 ( 
.A(n_10165),
.B(n_8799),
.Y(n_10599)
);

AOI22xp33_ASAP7_75t_L g10600 ( 
.A1(n_10388),
.A2(n_10405),
.B1(n_10467),
.B2(n_10464),
.Y(n_10600)
);

AND2x4_ASAP7_75t_L g10601 ( 
.A(n_10065),
.B(n_9908),
.Y(n_10601)
);

OAI22xp5_ASAP7_75t_L g10602 ( 
.A1(n_10225),
.A2(n_9617),
.B1(n_9687),
.B2(n_9561),
.Y(n_10602)
);

OAI22xp5_ASAP7_75t_SL g10603 ( 
.A1(n_10038),
.A2(n_6171),
.B1(n_6185),
.B2(n_6182),
.Y(n_10603)
);

INVx1_ASAP7_75t_L g10604 ( 
.A(n_9964),
.Y(n_10604)
);

INVx1_ASAP7_75t_L g10605 ( 
.A(n_9998),
.Y(n_10605)
);

HB1xp67_ASAP7_75t_L g10606 ( 
.A(n_10008),
.Y(n_10606)
);

AND2x4_ASAP7_75t_SL g10607 ( 
.A(n_9911),
.B(n_6179),
.Y(n_10607)
);

AND2x2_ASAP7_75t_L g10608 ( 
.A(n_9862),
.B(n_9547),
.Y(n_10608)
);

AND2x4_ASAP7_75t_L g10609 ( 
.A(n_10065),
.B(n_9568),
.Y(n_10609)
);

AND2x4_ASAP7_75t_L g10610 ( 
.A(n_9914),
.B(n_9579),
.Y(n_10610)
);

AND2x2_ASAP7_75t_L g10611 ( 
.A(n_10268),
.B(n_9580),
.Y(n_10611)
);

AND2x2_ASAP7_75t_L g10612 ( 
.A(n_10278),
.B(n_9583),
.Y(n_10612)
);

HB1xp67_ASAP7_75t_L g10613 ( 
.A(n_10008),
.Y(n_10613)
);

BUFx2_ASAP7_75t_L g10614 ( 
.A(n_9965),
.Y(n_10614)
);

AND2x4_ASAP7_75t_L g10615 ( 
.A(n_9879),
.B(n_9592),
.Y(n_10615)
);

INVx1_ASAP7_75t_L g10616 ( 
.A(n_10107),
.Y(n_10616)
);

NOR2x1_ASAP7_75t_SL g10617 ( 
.A(n_10339),
.B(n_5936),
.Y(n_10617)
);

INVx1_ASAP7_75t_L g10618 ( 
.A(n_9998),
.Y(n_10618)
);

AND2x2_ASAP7_75t_L g10619 ( 
.A(n_10283),
.B(n_9757),
.Y(n_10619)
);

INVx1_ASAP7_75t_L g10620 ( 
.A(n_10007),
.Y(n_10620)
);

AND2x4_ASAP7_75t_L g10621 ( 
.A(n_9879),
.B(n_8722),
.Y(n_10621)
);

INVx2_ASAP7_75t_L g10622 ( 
.A(n_10004),
.Y(n_10622)
);

AND2x2_ASAP7_75t_L g10623 ( 
.A(n_9965),
.B(n_9692),
.Y(n_10623)
);

BUFx2_ASAP7_75t_L g10624 ( 
.A(n_10210),
.Y(n_10624)
);

INVx1_ASAP7_75t_L g10625 ( 
.A(n_10007),
.Y(n_10625)
);

OR2x2_ASAP7_75t_L g10626 ( 
.A(n_9846),
.B(n_8803),
.Y(n_10626)
);

INVx1_ASAP7_75t_L g10627 ( 
.A(n_10010),
.Y(n_10627)
);

NOR2x1_ASAP7_75t_L g10628 ( 
.A(n_10142),
.B(n_9669),
.Y(n_10628)
);

AND2x2_ASAP7_75t_L g10629 ( 
.A(n_10221),
.B(n_9706),
.Y(n_10629)
);

INVx2_ASAP7_75t_L g10630 ( 
.A(n_10142),
.Y(n_10630)
);

HB1xp67_ASAP7_75t_L g10631 ( 
.A(n_9850),
.Y(n_10631)
);

NOR2xp33_ASAP7_75t_L g10632 ( 
.A(n_10089),
.B(n_5936),
.Y(n_10632)
);

INVx1_ASAP7_75t_L g10633 ( 
.A(n_10010),
.Y(n_10633)
);

AND2x2_ASAP7_75t_L g10634 ( 
.A(n_10181),
.B(n_10098),
.Y(n_10634)
);

AND2x2_ASAP7_75t_L g10635 ( 
.A(n_10100),
.B(n_9322),
.Y(n_10635)
);

AND2x2_ASAP7_75t_L g10636 ( 
.A(n_9966),
.B(n_9601),
.Y(n_10636)
);

AOI22xp33_ASAP7_75t_L g10637 ( 
.A1(n_10405),
.A2(n_9223),
.B1(n_9275),
.B2(n_9457),
.Y(n_10637)
);

AND2x4_ASAP7_75t_L g10638 ( 
.A(n_10160),
.B(n_8254),
.Y(n_10638)
);

INVx2_ASAP7_75t_L g10639 ( 
.A(n_10160),
.Y(n_10639)
);

AND2x2_ASAP7_75t_L g10640 ( 
.A(n_9969),
.B(n_6182),
.Y(n_10640)
);

INVx1_ASAP7_75t_L g10641 ( 
.A(n_9902),
.Y(n_10641)
);

AND2x2_ASAP7_75t_L g10642 ( 
.A(n_9972),
.B(n_6185),
.Y(n_10642)
);

NAND2xp5_ASAP7_75t_L g10643 ( 
.A(n_10476),
.B(n_8804),
.Y(n_10643)
);

INVx2_ASAP7_75t_L g10644 ( 
.A(n_9938),
.Y(n_10644)
);

INVx1_ASAP7_75t_L g10645 ( 
.A(n_9902),
.Y(n_10645)
);

INVx2_ASAP7_75t_L g10646 ( 
.A(n_9938),
.Y(n_10646)
);

AOI22xp33_ASAP7_75t_L g10647 ( 
.A1(n_10412),
.A2(n_10419),
.B1(n_10406),
.B2(n_10408),
.Y(n_10647)
);

INVx2_ASAP7_75t_L g10648 ( 
.A(n_9888),
.Y(n_10648)
);

AND2x2_ASAP7_75t_L g10649 ( 
.A(n_10176),
.B(n_6288),
.Y(n_10649)
);

INVx1_ASAP7_75t_L g10650 ( 
.A(n_9995),
.Y(n_10650)
);

INVx1_ASAP7_75t_L g10651 ( 
.A(n_10036),
.Y(n_10651)
);

NAND2xp5_ASAP7_75t_L g10652 ( 
.A(n_10085),
.B(n_8811),
.Y(n_10652)
);

OR2x2_ASAP7_75t_L g10653 ( 
.A(n_9852),
.B(n_8814),
.Y(n_10653)
);

INVx1_ASAP7_75t_L g10654 ( 
.A(n_9853),
.Y(n_10654)
);

INVx2_ASAP7_75t_L g10655 ( 
.A(n_9888),
.Y(n_10655)
);

OR2x2_ASAP7_75t_L g10656 ( 
.A(n_9852),
.B(n_8816),
.Y(n_10656)
);

AND2x2_ASAP7_75t_L g10657 ( 
.A(n_10176),
.B(n_6288),
.Y(n_10657)
);

AND2x2_ASAP7_75t_L g10658 ( 
.A(n_9925),
.B(n_6340),
.Y(n_10658)
);

INVx3_ASAP7_75t_L g10659 ( 
.A(n_10310),
.Y(n_10659)
);

AND2x2_ASAP7_75t_L g10660 ( 
.A(n_9917),
.B(n_6340),
.Y(n_10660)
);

AND2x2_ASAP7_75t_L g10661 ( 
.A(n_9955),
.B(n_6349),
.Y(n_10661)
);

OR2x2_ASAP7_75t_L g10662 ( 
.A(n_9926),
.B(n_9961),
.Y(n_10662)
);

AND2x4_ASAP7_75t_SL g10663 ( 
.A(n_10183),
.B(n_10081),
.Y(n_10663)
);

AND2x4_ASAP7_75t_L g10664 ( 
.A(n_9863),
.B(n_8254),
.Y(n_10664)
);

INVx1_ASAP7_75t_L g10665 ( 
.A(n_9859),
.Y(n_10665)
);

INVxp67_ASAP7_75t_SL g10666 ( 
.A(n_10081),
.Y(n_10666)
);

INVxp67_ASAP7_75t_SL g10667 ( 
.A(n_9848),
.Y(n_10667)
);

HB1xp67_ASAP7_75t_L g10668 ( 
.A(n_9891),
.Y(n_10668)
);

INVx1_ASAP7_75t_L g10669 ( 
.A(n_9860),
.Y(n_10669)
);

INVx2_ASAP7_75t_L g10670 ( 
.A(n_9863),
.Y(n_10670)
);

AND2x4_ASAP7_75t_L g10671 ( 
.A(n_10061),
.B(n_6349),
.Y(n_10671)
);

INVx2_ASAP7_75t_L g10672 ( 
.A(n_9954),
.Y(n_10672)
);

BUFx2_ASAP7_75t_SL g10673 ( 
.A(n_10203),
.Y(n_10673)
);

INVx2_ASAP7_75t_L g10674 ( 
.A(n_9991),
.Y(n_10674)
);

AND2x2_ASAP7_75t_SL g10675 ( 
.A(n_10409),
.B(n_10443),
.Y(n_10675)
);

INVx2_ASAP7_75t_L g10676 ( 
.A(n_9991),
.Y(n_10676)
);

NAND2xp5_ASAP7_75t_L g10677 ( 
.A(n_10085),
.B(n_8823),
.Y(n_10677)
);

INVx2_ASAP7_75t_L g10678 ( 
.A(n_10112),
.Y(n_10678)
);

INVx1_ASAP7_75t_SL g10679 ( 
.A(n_10210),
.Y(n_10679)
);

INVx2_ASAP7_75t_L g10680 ( 
.A(n_10125),
.Y(n_10680)
);

NAND2xp5_ASAP7_75t_L g10681 ( 
.A(n_10370),
.B(n_8838),
.Y(n_10681)
);

INVx1_ASAP7_75t_L g10682 ( 
.A(n_9868),
.Y(n_10682)
);

INVx1_ASAP7_75t_L g10683 ( 
.A(n_9871),
.Y(n_10683)
);

AND2x2_ASAP7_75t_L g10684 ( 
.A(n_10331),
.B(n_9635),
.Y(n_10684)
);

AOI22xp33_ASAP7_75t_L g10685 ( 
.A1(n_10412),
.A2(n_10419),
.B1(n_10425),
.B2(n_10456),
.Y(n_10685)
);

OR2x2_ASAP7_75t_L g10686 ( 
.A(n_9926),
.B(n_8841),
.Y(n_10686)
);

NAND2xp5_ASAP7_75t_L g10687 ( 
.A(n_10453),
.B(n_8842),
.Y(n_10687)
);

AND2x2_ASAP7_75t_L g10688 ( 
.A(n_9856),
.B(n_9577),
.Y(n_10688)
);

OR2x2_ASAP7_75t_L g10689 ( 
.A(n_9961),
.B(n_8843),
.Y(n_10689)
);

AND2x2_ASAP7_75t_L g10690 ( 
.A(n_9856),
.B(n_8847),
.Y(n_10690)
);

NAND3xp33_ASAP7_75t_L g10691 ( 
.A(n_10260),
.B(n_9743),
.C(n_9590),
.Y(n_10691)
);

NAND2xp5_ASAP7_75t_L g10692 ( 
.A(n_10391),
.B(n_8854),
.Y(n_10692)
);

INVx1_ASAP7_75t_L g10693 ( 
.A(n_9875),
.Y(n_10693)
);

AND2x2_ASAP7_75t_L g10694 ( 
.A(n_9886),
.B(n_8857),
.Y(n_10694)
);

HB1xp67_ASAP7_75t_L g10695 ( 
.A(n_9941),
.Y(n_10695)
);

INVx1_ASAP7_75t_L g10696 ( 
.A(n_9878),
.Y(n_10696)
);

INVx2_ASAP7_75t_L g10697 ( 
.A(n_9865),
.Y(n_10697)
);

NAND2xp5_ASAP7_75t_L g10698 ( 
.A(n_10260),
.B(n_8861),
.Y(n_10698)
);

INVx1_ASAP7_75t_L g10699 ( 
.A(n_9880),
.Y(n_10699)
);

NOR2xp33_ASAP7_75t_L g10700 ( 
.A(n_10203),
.B(n_5936),
.Y(n_10700)
);

BUFx3_ASAP7_75t_L g10701 ( 
.A(n_9985),
.Y(n_10701)
);

INVx3_ASAP7_75t_SL g10702 ( 
.A(n_10186),
.Y(n_10702)
);

AND2x2_ASAP7_75t_L g10703 ( 
.A(n_10096),
.B(n_8864),
.Y(n_10703)
);

AND2x2_ASAP7_75t_L g10704 ( 
.A(n_10096),
.B(n_9956),
.Y(n_10704)
);

INVx1_ASAP7_75t_L g10705 ( 
.A(n_9882),
.Y(n_10705)
);

AND2x2_ASAP7_75t_L g10706 ( 
.A(n_9957),
.B(n_8866),
.Y(n_10706)
);

INVx2_ASAP7_75t_L g10707 ( 
.A(n_9866),
.Y(n_10707)
);

INVx5_ASAP7_75t_L g10708 ( 
.A(n_10126),
.Y(n_10708)
);

INVx2_ASAP7_75t_L g10709 ( 
.A(n_9870),
.Y(n_10709)
);

AND2x2_ASAP7_75t_L g10710 ( 
.A(n_9980),
.B(n_8868),
.Y(n_10710)
);

AND2x2_ASAP7_75t_L g10711 ( 
.A(n_9984),
.B(n_8870),
.Y(n_10711)
);

HB1xp67_ASAP7_75t_L g10712 ( 
.A(n_9874),
.Y(n_10712)
);

INVx1_ASAP7_75t_L g10713 ( 
.A(n_9884),
.Y(n_10713)
);

INVx2_ASAP7_75t_L g10714 ( 
.A(n_10072),
.Y(n_10714)
);

AND2x4_ASAP7_75t_SL g10715 ( 
.A(n_9869),
.B(n_6665),
.Y(n_10715)
);

AND2x2_ASAP7_75t_L g10716 ( 
.A(n_10320),
.B(n_8872),
.Y(n_10716)
);

AND2x2_ASAP7_75t_L g10717 ( 
.A(n_9986),
.B(n_8875),
.Y(n_10717)
);

INVx1_ASAP7_75t_L g10718 ( 
.A(n_9887),
.Y(n_10718)
);

INVx1_ASAP7_75t_L g10719 ( 
.A(n_10114),
.Y(n_10719)
);

INVx1_ASAP7_75t_L g10720 ( 
.A(n_10114),
.Y(n_10720)
);

AND2x2_ASAP7_75t_L g10721 ( 
.A(n_9989),
.B(n_8882),
.Y(n_10721)
);

NAND2xp5_ASAP7_75t_L g10722 ( 
.A(n_10038),
.B(n_8883),
.Y(n_10722)
);

INVxp67_ASAP7_75t_L g10723 ( 
.A(n_10178),
.Y(n_10723)
);

OAI22xp33_ASAP7_75t_L g10724 ( 
.A1(n_10032),
.A2(n_9567),
.B1(n_9406),
.B2(n_9332),
.Y(n_10724)
);

OR2x2_ASAP7_75t_L g10725 ( 
.A(n_10400),
.B(n_8884),
.Y(n_10725)
);

AND2x2_ASAP7_75t_L g10726 ( 
.A(n_9992),
.B(n_8888),
.Y(n_10726)
);

AND2x2_ASAP7_75t_L g10727 ( 
.A(n_10358),
.B(n_8891),
.Y(n_10727)
);

INVx1_ASAP7_75t_L g10728 ( 
.A(n_9940),
.Y(n_10728)
);

OR2x2_ASAP7_75t_L g10729 ( 
.A(n_10254),
.B(n_8892),
.Y(n_10729)
);

AND2x4_ASAP7_75t_SL g10730 ( 
.A(n_9897),
.B(n_6665),
.Y(n_10730)
);

BUFx2_ASAP7_75t_L g10731 ( 
.A(n_10358),
.Y(n_10731)
);

INVx1_ASAP7_75t_L g10732 ( 
.A(n_10124),
.Y(n_10732)
);

INVx1_ASAP7_75t_SL g10733 ( 
.A(n_10252),
.Y(n_10733)
);

AND2x2_ASAP7_75t_L g10734 ( 
.A(n_10243),
.B(n_10265),
.Y(n_10734)
);

INVx1_ASAP7_75t_L g10735 ( 
.A(n_10124),
.Y(n_10735)
);

BUFx2_ASAP7_75t_L g10736 ( 
.A(n_10274),
.Y(n_10736)
);

AND2x2_ASAP7_75t_L g10737 ( 
.A(n_10266),
.B(n_8893),
.Y(n_10737)
);

INVx1_ASAP7_75t_L g10738 ( 
.A(n_10250),
.Y(n_10738)
);

AND2x2_ASAP7_75t_L g10739 ( 
.A(n_9903),
.B(n_8896),
.Y(n_10739)
);

AND2x2_ASAP7_75t_L g10740 ( 
.A(n_10267),
.B(n_8905),
.Y(n_10740)
);

INVx1_ASAP7_75t_L g10741 ( 
.A(n_10250),
.Y(n_10741)
);

AND2x2_ASAP7_75t_L g10742 ( 
.A(n_9975),
.B(n_8907),
.Y(n_10742)
);

AND2x2_ASAP7_75t_L g10743 ( 
.A(n_10015),
.B(n_8922),
.Y(n_10743)
);

AOI22xp5_ASAP7_75t_L g10744 ( 
.A1(n_10032),
.A2(n_9383),
.B1(n_9389),
.B2(n_9357),
.Y(n_10744)
);

INVx1_ASAP7_75t_L g10745 ( 
.A(n_10369),
.Y(n_10745)
);

INVx1_ASAP7_75t_L g10746 ( 
.A(n_10369),
.Y(n_10746)
);

AND2x2_ASAP7_75t_L g10747 ( 
.A(n_10015),
.B(n_8932),
.Y(n_10747)
);

NAND2xp5_ASAP7_75t_L g10748 ( 
.A(n_9858),
.B(n_10483),
.Y(n_10748)
);

HB1xp67_ASAP7_75t_L g10749 ( 
.A(n_10276),
.Y(n_10749)
);

AND2x2_ASAP7_75t_L g10750 ( 
.A(n_10410),
.B(n_8937),
.Y(n_10750)
);

OR2x2_ASAP7_75t_L g10751 ( 
.A(n_9996),
.B(n_8939),
.Y(n_10751)
);

AND2x2_ASAP7_75t_L g10752 ( 
.A(n_10410),
.B(n_8942),
.Y(n_10752)
);

AND2x2_ASAP7_75t_L g10753 ( 
.A(n_10427),
.B(n_8946),
.Y(n_10753)
);

INVx2_ASAP7_75t_SL g10754 ( 
.A(n_10252),
.Y(n_10754)
);

INVx1_ASAP7_75t_L g10755 ( 
.A(n_9889),
.Y(n_10755)
);

INVxp67_ASAP7_75t_L g10756 ( 
.A(n_10048),
.Y(n_10756)
);

INVx2_ASAP7_75t_L g10757 ( 
.A(n_10072),
.Y(n_10757)
);

OAI22xp5_ASAP7_75t_L g10758 ( 
.A1(n_10225),
.A2(n_9623),
.B1(n_9652),
.B2(n_9352),
.Y(n_10758)
);

INVx1_ASAP7_75t_L g10759 ( 
.A(n_9895),
.Y(n_10759)
);

AND2x2_ASAP7_75t_L g10760 ( 
.A(n_10427),
.B(n_8950),
.Y(n_10760)
);

INVx2_ASAP7_75t_L g10761 ( 
.A(n_10208),
.Y(n_10761)
);

AND2x2_ASAP7_75t_L g10762 ( 
.A(n_10000),
.B(n_8952),
.Y(n_10762)
);

INVx1_ASAP7_75t_L g10763 ( 
.A(n_10034),
.Y(n_10763)
);

INVx1_ASAP7_75t_L g10764 ( 
.A(n_10034),
.Y(n_10764)
);

INVx1_ASAP7_75t_L g10765 ( 
.A(n_9983),
.Y(n_10765)
);

AND2x2_ASAP7_75t_L g10766 ( 
.A(n_10229),
.B(n_8954),
.Y(n_10766)
);

INVx1_ASAP7_75t_L g10767 ( 
.A(n_9983),
.Y(n_10767)
);

INVx1_ASAP7_75t_L g10768 ( 
.A(n_10315),
.Y(n_10768)
);

AND2x4_ASAP7_75t_L g10769 ( 
.A(n_10126),
.B(n_8608),
.Y(n_10769)
);

AND2x2_ASAP7_75t_L g10770 ( 
.A(n_10057),
.B(n_10090),
.Y(n_10770)
);

INVx1_ASAP7_75t_L g10771 ( 
.A(n_10315),
.Y(n_10771)
);

AND2x2_ASAP7_75t_L g10772 ( 
.A(n_10057),
.B(n_8959),
.Y(n_10772)
);

INVx2_ASAP7_75t_L g10773 ( 
.A(n_10213),
.Y(n_10773)
);

AND2x4_ASAP7_75t_L g10774 ( 
.A(n_10134),
.B(n_8608),
.Y(n_10774)
);

INVx1_ASAP7_75t_L g10775 ( 
.A(n_10323),
.Y(n_10775)
);

AND2x2_ASAP7_75t_L g10776 ( 
.A(n_10092),
.B(n_8960),
.Y(n_10776)
);

INVx2_ASAP7_75t_L g10777 ( 
.A(n_10217),
.Y(n_10777)
);

INVx1_ASAP7_75t_L g10778 ( 
.A(n_10325),
.Y(n_10778)
);

AND2x2_ASAP7_75t_L g10779 ( 
.A(n_10282),
.B(n_8961),
.Y(n_10779)
);

INVx2_ASAP7_75t_L g10780 ( 
.A(n_10215),
.Y(n_10780)
);

INVx1_ASAP7_75t_L g10781 ( 
.A(n_9979),
.Y(n_10781)
);

BUFx3_ASAP7_75t_L g10782 ( 
.A(n_10218),
.Y(n_10782)
);

AND2x2_ASAP7_75t_L g10783 ( 
.A(n_10322),
.B(n_8964),
.Y(n_10783)
);

AND2x2_ASAP7_75t_L g10784 ( 
.A(n_10322),
.B(n_8966),
.Y(n_10784)
);

NOR2xp33_ASAP7_75t_L g10785 ( 
.A(n_10134),
.B(n_6406),
.Y(n_10785)
);

INVx1_ASAP7_75t_L g10786 ( 
.A(n_9979),
.Y(n_10786)
);

NOR2x1p5_ASAP7_75t_L g10787 ( 
.A(n_9960),
.B(n_6406),
.Y(n_10787)
);

INVx1_ASAP7_75t_L g10788 ( 
.A(n_10013),
.Y(n_10788)
);

AND2x2_ASAP7_75t_L g10789 ( 
.A(n_10163),
.B(n_8967),
.Y(n_10789)
);

INVx3_ASAP7_75t_L g10790 ( 
.A(n_10310),
.Y(n_10790)
);

NAND2xp5_ASAP7_75t_L g10791 ( 
.A(n_9848),
.B(n_8971),
.Y(n_10791)
);

INVx1_ASAP7_75t_L g10792 ( 
.A(n_10013),
.Y(n_10792)
);

AOI22xp33_ASAP7_75t_L g10793 ( 
.A1(n_10127),
.A2(n_9426),
.B1(n_9464),
.B2(n_9456),
.Y(n_10793)
);

NAND2xp5_ASAP7_75t_L g10794 ( 
.A(n_9973),
.B(n_8977),
.Y(n_10794)
);

INVx1_ASAP7_75t_L g10795 ( 
.A(n_10242),
.Y(n_10795)
);

CKINVDCx20_ASAP7_75t_R g10796 ( 
.A(n_10269),
.Y(n_10796)
);

AOI22xp33_ASAP7_75t_L g10797 ( 
.A1(n_10127),
.A2(n_9339),
.B1(n_9345),
.B2(n_9342),
.Y(n_10797)
);

AND2x2_ASAP7_75t_L g10798 ( 
.A(n_10163),
.B(n_8983),
.Y(n_10798)
);

INVx2_ASAP7_75t_L g10799 ( 
.A(n_10062),
.Y(n_10799)
);

NAND2xp5_ASAP7_75t_L g10800 ( 
.A(n_9981),
.B(n_8998),
.Y(n_10800)
);

INVx2_ASAP7_75t_L g10801 ( 
.A(n_10071),
.Y(n_10801)
);

OR2x2_ASAP7_75t_L g10802 ( 
.A(n_10313),
.B(n_9014),
.Y(n_10802)
);

INVx2_ASAP7_75t_L g10803 ( 
.A(n_10074),
.Y(n_10803)
);

INVx2_ASAP7_75t_L g10804 ( 
.A(n_10075),
.Y(n_10804)
);

INVx2_ASAP7_75t_L g10805 ( 
.A(n_10080),
.Y(n_10805)
);

AOI21xp33_ASAP7_75t_L g10806 ( 
.A1(n_10437),
.A2(n_9438),
.B(n_9416),
.Y(n_10806)
);

INVx1_ASAP7_75t_L g10807 ( 
.A(n_9999),
.Y(n_10807)
);

AND2x2_ASAP7_75t_L g10808 ( 
.A(n_10247),
.B(n_9017),
.Y(n_10808)
);

INVx1_ASAP7_75t_L g10809 ( 
.A(n_10006),
.Y(n_10809)
);

HB1xp67_ASAP7_75t_L g10810 ( 
.A(n_10276),
.Y(n_10810)
);

AND2x2_ASAP7_75t_L g10811 ( 
.A(n_10247),
.B(n_9030),
.Y(n_10811)
);

NAND2xp5_ASAP7_75t_L g10812 ( 
.A(n_9988),
.B(n_9031),
.Y(n_10812)
);

AOI22xp33_ASAP7_75t_SL g10813 ( 
.A1(n_10383),
.A2(n_9838),
.B1(n_9737),
.B2(n_9540),
.Y(n_10813)
);

AND2x2_ASAP7_75t_L g10814 ( 
.A(n_10202),
.B(n_9032),
.Y(n_10814)
);

NOR2xp33_ASAP7_75t_L g10815 ( 
.A(n_10188),
.B(n_10206),
.Y(n_10815)
);

AND2x2_ASAP7_75t_L g10816 ( 
.A(n_10046),
.B(n_9033),
.Y(n_10816)
);

AND2x4_ASAP7_75t_L g10817 ( 
.A(n_10188),
.B(n_8622),
.Y(n_10817)
);

INVx1_ASAP7_75t_L g10818 ( 
.A(n_10246),
.Y(n_10818)
);

HB1xp67_ASAP7_75t_L g10819 ( 
.A(n_10279),
.Y(n_10819)
);

INVx2_ASAP7_75t_L g10820 ( 
.A(n_10191),
.Y(n_10820)
);

INVx1_ASAP7_75t_L g10821 ( 
.A(n_10171),
.Y(n_10821)
);

INVx3_ASAP7_75t_L g10822 ( 
.A(n_9849),
.Y(n_10822)
);

AND2x2_ASAP7_75t_L g10823 ( 
.A(n_10280),
.B(n_9036),
.Y(n_10823)
);

OR2x2_ASAP7_75t_L g10824 ( 
.A(n_10313),
.B(n_9045),
.Y(n_10824)
);

AND2x2_ASAP7_75t_L g10825 ( 
.A(n_9918),
.B(n_9047),
.Y(n_10825)
);

NAND2xp5_ASAP7_75t_L g10826 ( 
.A(n_10378),
.B(n_9053),
.Y(n_10826)
);

INVx2_ASAP7_75t_L g10827 ( 
.A(n_10196),
.Y(n_10827)
);

INVx1_ASAP7_75t_L g10828 ( 
.A(n_10292),
.Y(n_10828)
);

INVx1_ASAP7_75t_L g10829 ( 
.A(n_10294),
.Y(n_10829)
);

INVx2_ASAP7_75t_L g10830 ( 
.A(n_10211),
.Y(n_10830)
);

INVx1_ASAP7_75t_L g10831 ( 
.A(n_10026),
.Y(n_10831)
);

AND2x2_ASAP7_75t_L g10832 ( 
.A(n_10052),
.B(n_9056),
.Y(n_10832)
);

HB1xp67_ASAP7_75t_L g10833 ( 
.A(n_10279),
.Y(n_10833)
);

AND2x2_ASAP7_75t_L g10834 ( 
.A(n_10055),
.B(n_9058),
.Y(n_10834)
);

OR2x2_ASAP7_75t_L g10835 ( 
.A(n_10431),
.B(n_10348),
.Y(n_10835)
);

INVx1_ASAP7_75t_L g10836 ( 
.A(n_10067),
.Y(n_10836)
);

INVx1_ASAP7_75t_L g10837 ( 
.A(n_10086),
.Y(n_10837)
);

AND2x2_ASAP7_75t_L g10838 ( 
.A(n_10284),
.B(n_9062),
.Y(n_10838)
);

NOR2x1p5_ASAP7_75t_L g10839 ( 
.A(n_10206),
.B(n_6419),
.Y(n_10839)
);

OR2x2_ASAP7_75t_L g10840 ( 
.A(n_10431),
.B(n_9063),
.Y(n_10840)
);

AND2x4_ASAP7_75t_L g10841 ( 
.A(n_10204),
.B(n_8622),
.Y(n_10841)
);

AND2x2_ASAP7_75t_L g10842 ( 
.A(n_9877),
.B(n_10340),
.Y(n_10842)
);

NOR2xp33_ASAP7_75t_L g10843 ( 
.A(n_10269),
.B(n_6419),
.Y(n_10843)
);

OR2x2_ASAP7_75t_L g10844 ( 
.A(n_10348),
.B(n_9066),
.Y(n_10844)
);

INVx2_ASAP7_75t_L g10845 ( 
.A(n_10212),
.Y(n_10845)
);

INVx1_ASAP7_75t_L g10846 ( 
.A(n_9899),
.Y(n_10846)
);

INVx3_ASAP7_75t_L g10847 ( 
.A(n_10180),
.Y(n_10847)
);

NAND2xp5_ASAP7_75t_L g10848 ( 
.A(n_10378),
.B(n_9067),
.Y(n_10848)
);

AND2x2_ASAP7_75t_L g10849 ( 
.A(n_10150),
.B(n_9069),
.Y(n_10849)
);

BUFx2_ASAP7_75t_L g10850 ( 
.A(n_10274),
.Y(n_10850)
);

AND2x2_ASAP7_75t_L g10851 ( 
.A(n_10152),
.B(n_9070),
.Y(n_10851)
);

NAND2x1p5_ASAP7_75t_SL g10852 ( 
.A(n_10029),
.B(n_8413),
.Y(n_10852)
);

AND2x2_ASAP7_75t_L g10853 ( 
.A(n_10156),
.B(n_9073),
.Y(n_10853)
);

INVx1_ASAP7_75t_L g10854 ( 
.A(n_9901),
.Y(n_10854)
);

INVx1_ASAP7_75t_L g10855 ( 
.A(n_9909),
.Y(n_10855)
);

NAND2xp5_ASAP7_75t_L g10856 ( 
.A(n_10159),
.B(n_9074),
.Y(n_10856)
);

HB1xp67_ASAP7_75t_L g10857 ( 
.A(n_10220),
.Y(n_10857)
);

INVx2_ASAP7_75t_L g10858 ( 
.A(n_10288),
.Y(n_10858)
);

INVx2_ASAP7_75t_L g10859 ( 
.A(n_10290),
.Y(n_10859)
);

OR2x2_ASAP7_75t_L g10860 ( 
.A(n_10017),
.B(n_9075),
.Y(n_10860)
);

BUFx2_ASAP7_75t_SL g10861 ( 
.A(n_10105),
.Y(n_10861)
);

OR2x2_ASAP7_75t_L g10862 ( 
.A(n_10137),
.B(n_9076),
.Y(n_10862)
);

INVx2_ASAP7_75t_L g10863 ( 
.A(n_10341),
.Y(n_10863)
);

INVx1_ASAP7_75t_L g10864 ( 
.A(n_9912),
.Y(n_10864)
);

INVx1_ASAP7_75t_L g10865 ( 
.A(n_9913),
.Y(n_10865)
);

INVx3_ASAP7_75t_L g10866 ( 
.A(n_9971),
.Y(n_10866)
);

INVx1_ASAP7_75t_SL g10867 ( 
.A(n_10087),
.Y(n_10867)
);

AND2x4_ASAP7_75t_SL g10868 ( 
.A(n_10113),
.B(n_6665),
.Y(n_10868)
);

INVx1_ASAP7_75t_L g10869 ( 
.A(n_9916),
.Y(n_10869)
);

INVx2_ASAP7_75t_L g10870 ( 
.A(n_10223),
.Y(n_10870)
);

NAND2xp5_ASAP7_75t_L g10871 ( 
.A(n_10164),
.B(n_9081),
.Y(n_10871)
);

NAND2xp5_ASAP7_75t_L g10872 ( 
.A(n_10053),
.B(n_9082),
.Y(n_10872)
);

INVx2_ASAP7_75t_L g10873 ( 
.A(n_10226),
.Y(n_10873)
);

INVx1_ASAP7_75t_L g10874 ( 
.A(n_9919),
.Y(n_10874)
);

INVx2_ASAP7_75t_L g10875 ( 
.A(n_10235),
.Y(n_10875)
);

BUFx3_ASAP7_75t_L g10876 ( 
.A(n_10123),
.Y(n_10876)
);

OAI22xp5_ASAP7_75t_L g10877 ( 
.A1(n_10227),
.A2(n_9640),
.B1(n_9445),
.B2(n_9195),
.Y(n_10877)
);

INVx1_ASAP7_75t_L g10878 ( 
.A(n_9923),
.Y(n_10878)
);

INVx1_ASAP7_75t_L g10879 ( 
.A(n_9933),
.Y(n_10879)
);

AND2x2_ASAP7_75t_L g10880 ( 
.A(n_10157),
.B(n_9083),
.Y(n_10880)
);

INVx1_ASAP7_75t_L g10881 ( 
.A(n_9934),
.Y(n_10881)
);

AND2x2_ASAP7_75t_L g10882 ( 
.A(n_10174),
.B(n_9084),
.Y(n_10882)
);

AOI22xp33_ASAP7_75t_L g10883 ( 
.A1(n_10371),
.A2(n_9328),
.B1(n_9325),
.B2(n_9169),
.Y(n_10883)
);

NAND2xp5_ASAP7_75t_L g10884 ( 
.A(n_10053),
.B(n_9088),
.Y(n_10884)
);

OR2x2_ASAP7_75t_L g10885 ( 
.A(n_10137),
.B(n_9089),
.Y(n_10885)
);

AND2x4_ASAP7_75t_L g10886 ( 
.A(n_10003),
.B(n_9090),
.Y(n_10886)
);

NAND2xp5_ASAP7_75t_L g10887 ( 
.A(n_10435),
.B(n_9092),
.Y(n_10887)
);

INVx2_ASAP7_75t_L g10888 ( 
.A(n_10240),
.Y(n_10888)
);

INVx2_ASAP7_75t_SL g10889 ( 
.A(n_10172),
.Y(n_10889)
);

AND2x2_ASAP7_75t_L g10890 ( 
.A(n_10350),
.B(n_9095),
.Y(n_10890)
);

NAND2xp5_ASAP7_75t_L g10891 ( 
.A(n_10104),
.B(n_9099),
.Y(n_10891)
);

AND2x2_ASAP7_75t_L g10892 ( 
.A(n_10354),
.B(n_9104),
.Y(n_10892)
);

INVx2_ASAP7_75t_L g10893 ( 
.A(n_10241),
.Y(n_10893)
);

NOR2x1_ASAP7_75t_SL g10894 ( 
.A(n_10339),
.B(n_9783),
.Y(n_10894)
);

AND2x2_ASAP7_75t_L g10895 ( 
.A(n_10162),
.B(n_10190),
.Y(n_10895)
);

BUFx2_ASAP7_75t_L g10896 ( 
.A(n_9971),
.Y(n_10896)
);

AND2x2_ASAP7_75t_L g10897 ( 
.A(n_10021),
.B(n_9108),
.Y(n_10897)
);

INVx2_ASAP7_75t_L g10898 ( 
.A(n_10244),
.Y(n_10898)
);

INVx1_ASAP7_75t_L g10899 ( 
.A(n_9936),
.Y(n_10899)
);

INVx1_ASAP7_75t_L g10900 ( 
.A(n_9942),
.Y(n_10900)
);

AOI22xp33_ASAP7_75t_L g10901 ( 
.A1(n_10227),
.A2(n_9657),
.B1(n_9659),
.B2(n_9392),
.Y(n_10901)
);

AND2x2_ASAP7_75t_L g10902 ( 
.A(n_10024),
.B(n_9112),
.Y(n_10902)
);

INVx2_ASAP7_75t_L g10903 ( 
.A(n_10245),
.Y(n_10903)
);

AND2x4_ASAP7_75t_SL g10904 ( 
.A(n_10012),
.B(n_6665),
.Y(n_10904)
);

AND2x2_ASAP7_75t_L g10905 ( 
.A(n_10385),
.B(n_9114),
.Y(n_10905)
);

AND2x2_ASAP7_75t_L g10906 ( 
.A(n_10356),
.B(n_9118),
.Y(n_10906)
);

INVx1_ASAP7_75t_L g10907 ( 
.A(n_10311),
.Y(n_10907)
);

INVx1_ASAP7_75t_L g10908 ( 
.A(n_9946),
.Y(n_10908)
);

INVx1_ASAP7_75t_L g10909 ( 
.A(n_9947),
.Y(n_10909)
);

AND2x4_ASAP7_75t_L g10910 ( 
.A(n_10169),
.B(n_9119),
.Y(n_10910)
);

AND2x2_ASAP7_75t_L g10911 ( 
.A(n_10028),
.B(n_9123),
.Y(n_10911)
);

NOR2xp33_ASAP7_75t_L g10912 ( 
.A(n_10289),
.B(n_9733),
.Y(n_10912)
);

OR2x2_ASAP7_75t_L g10913 ( 
.A(n_10338),
.B(n_10343),
.Y(n_10913)
);

OR2x2_ASAP7_75t_L g10914 ( 
.A(n_10338),
.B(n_9126),
.Y(n_10914)
);

NAND2xp5_ASAP7_75t_L g10915 ( 
.A(n_10104),
.B(n_9128),
.Y(n_10915)
);

INVx1_ASAP7_75t_L g10916 ( 
.A(n_9950),
.Y(n_10916)
);

BUFx8_ASAP7_75t_L g10917 ( 
.A(n_10111),
.Y(n_10917)
);

INVx2_ASAP7_75t_L g10918 ( 
.A(n_10189),
.Y(n_10918)
);

BUFx2_ASAP7_75t_L g10919 ( 
.A(n_10445),
.Y(n_10919)
);

BUFx3_ASAP7_75t_L g10920 ( 
.A(n_10330),
.Y(n_10920)
);

INVx3_ASAP7_75t_R g10921 ( 
.A(n_10393),
.Y(n_10921)
);

INVx1_ASAP7_75t_L g10922 ( 
.A(n_9959),
.Y(n_10922)
);

AND2x2_ASAP7_75t_L g10923 ( 
.A(n_10030),
.B(n_9130),
.Y(n_10923)
);

AND2x2_ASAP7_75t_L g10924 ( 
.A(n_10040),
.B(n_9136),
.Y(n_10924)
);

AND2x2_ASAP7_75t_L g10925 ( 
.A(n_10321),
.B(n_9139),
.Y(n_10925)
);

BUFx2_ASAP7_75t_L g10926 ( 
.A(n_10445),
.Y(n_10926)
);

INVx1_ASAP7_75t_L g10927 ( 
.A(n_9963),
.Y(n_10927)
);

INVx2_ASAP7_75t_L g10928 ( 
.A(n_9943),
.Y(n_10928)
);

AND2x2_ASAP7_75t_L g10929 ( 
.A(n_10304),
.B(n_9147),
.Y(n_10929)
);

INVx1_ASAP7_75t_SL g10930 ( 
.A(n_10172),
.Y(n_10930)
);

AND2x2_ASAP7_75t_L g10931 ( 
.A(n_10317),
.B(n_9154),
.Y(n_10931)
);

INVx2_ASAP7_75t_L g10932 ( 
.A(n_9944),
.Y(n_10932)
);

INVx1_ASAP7_75t_L g10933 ( 
.A(n_9968),
.Y(n_10933)
);

AND2x2_ASAP7_75t_L g10934 ( 
.A(n_10131),
.B(n_10144),
.Y(n_10934)
);

AND2x2_ASAP7_75t_L g10935 ( 
.A(n_9953),
.B(n_9158),
.Y(n_10935)
);

AND2x2_ASAP7_75t_L g10936 ( 
.A(n_10324),
.B(n_9161),
.Y(n_10936)
);

AND2x4_ASAP7_75t_L g10937 ( 
.A(n_10451),
.B(n_10455),
.Y(n_10937)
);

INVx1_ASAP7_75t_L g10938 ( 
.A(n_9974),
.Y(n_10938)
);

AND2x2_ASAP7_75t_L g10939 ( 
.A(n_9904),
.B(n_6496),
.Y(n_10939)
);

AND2x2_ASAP7_75t_L g10940 ( 
.A(n_9924),
.B(n_6496),
.Y(n_10940)
);

INVxp67_ASAP7_75t_L g10941 ( 
.A(n_10289),
.Y(n_10941)
);

INVx2_ASAP7_75t_L g10942 ( 
.A(n_10451),
.Y(n_10942)
);

NAND2xp5_ASAP7_75t_L g10943 ( 
.A(n_10362),
.B(n_9203),
.Y(n_10943)
);

AND2x2_ASAP7_75t_L g10944 ( 
.A(n_9927),
.B(n_6496),
.Y(n_10944)
);

HB1xp67_ASAP7_75t_L g10945 ( 
.A(n_10386),
.Y(n_10945)
);

INVx2_ASAP7_75t_L g10946 ( 
.A(n_10455),
.Y(n_10946)
);

AND2x4_ASAP7_75t_L g10947 ( 
.A(n_10473),
.B(n_9698),
.Y(n_10947)
);

BUFx2_ASAP7_75t_L g10948 ( 
.A(n_10473),
.Y(n_10948)
);

INVx2_ASAP7_75t_L g10949 ( 
.A(n_10480),
.Y(n_10949)
);

INVx1_ASAP7_75t_L g10950 ( 
.A(n_9976),
.Y(n_10950)
);

AND2x2_ASAP7_75t_L g10951 ( 
.A(n_9932),
.B(n_9937),
.Y(n_10951)
);

INVx1_ASAP7_75t_L g10952 ( 
.A(n_9982),
.Y(n_10952)
);

INVx2_ASAP7_75t_L g10953 ( 
.A(n_10480),
.Y(n_10953)
);

AND2x2_ASAP7_75t_L g10954 ( 
.A(n_9939),
.B(n_6496),
.Y(n_10954)
);

AOI221xp5_ASAP7_75t_L g10955 ( 
.A1(n_10484),
.A2(n_9494),
.B1(n_9344),
.B2(n_9590),
.C(n_9587),
.Y(n_10955)
);

INVx1_ASAP7_75t_L g10956 ( 
.A(n_9987),
.Y(n_10956)
);

INVx1_ASAP7_75t_L g10957 ( 
.A(n_9994),
.Y(n_10957)
);

AND2x2_ASAP7_75t_L g10958 ( 
.A(n_10328),
.B(n_6496),
.Y(n_10958)
);

INVx1_ASAP7_75t_L g10959 ( 
.A(n_10005),
.Y(n_10959)
);

AND2x2_ASAP7_75t_L g10960 ( 
.A(n_10367),
.B(n_6528),
.Y(n_10960)
);

BUFx3_ASAP7_75t_L g10961 ( 
.A(n_10330),
.Y(n_10961)
);

AND2x2_ASAP7_75t_L g10962 ( 
.A(n_10379),
.B(n_10424),
.Y(n_10962)
);

INVx1_ASAP7_75t_L g10963 ( 
.A(n_10019),
.Y(n_10963)
);

INVx2_ASAP7_75t_L g10964 ( 
.A(n_10043),
.Y(n_10964)
);

INVx1_ASAP7_75t_L g10965 ( 
.A(n_10020),
.Y(n_10965)
);

AOI22xp33_ASAP7_75t_L g10966 ( 
.A1(n_10442),
.A2(n_9331),
.B1(n_9787),
.B2(n_9774),
.Y(n_10966)
);

INVx1_ASAP7_75t_L g10967 ( 
.A(n_10016),
.Y(n_10967)
);

INVx1_ASAP7_75t_L g10968 ( 
.A(n_10233),
.Y(n_10968)
);

AND2x4_ASAP7_75t_SL g10969 ( 
.A(n_10393),
.B(n_6847),
.Y(n_10969)
);

NAND2xp5_ASAP7_75t_L g10970 ( 
.A(n_10179),
.B(n_6806),
.Y(n_10970)
);

NAND2xp5_ASAP7_75t_L g10971 ( 
.A(n_10484),
.B(n_6806),
.Y(n_10971)
);

HB1xp67_ASAP7_75t_L g10972 ( 
.A(n_10141),
.Y(n_10972)
);

INVx2_ASAP7_75t_SL g10973 ( 
.A(n_10207),
.Y(n_10973)
);

INVx2_ASAP7_75t_L g10974 ( 
.A(n_10120),
.Y(n_10974)
);

INVx2_ASAP7_75t_L g10975 ( 
.A(n_10177),
.Y(n_10975)
);

AND2x4_ASAP7_75t_SL g10976 ( 
.A(n_10301),
.B(n_6847),
.Y(n_10976)
);

AND2x2_ASAP7_75t_L g10977 ( 
.A(n_10424),
.B(n_6528),
.Y(n_10977)
);

INVx4_ASAP7_75t_L g10978 ( 
.A(n_10368),
.Y(n_10978)
);

NAND2xp5_ASAP7_75t_L g10979 ( 
.A(n_10403),
.B(n_10023),
.Y(n_10979)
);

AND2x2_ASAP7_75t_L g10980 ( 
.A(n_10083),
.B(n_6528),
.Y(n_10980)
);

INVx1_ASAP7_75t_L g10981 ( 
.A(n_10234),
.Y(n_10981)
);

NOR2x1p5_ASAP7_75t_L g10982 ( 
.A(n_10458),
.B(n_8449),
.Y(n_10982)
);

INVx1_ASAP7_75t_L g10983 ( 
.A(n_10236),
.Y(n_10983)
);

INVx2_ASAP7_75t_L g10984 ( 
.A(n_10095),
.Y(n_10984)
);

NOR2xp33_ASAP7_75t_L g10985 ( 
.A(n_10397),
.B(n_8054),
.Y(n_10985)
);

INVx1_ASAP7_75t_L g10986 ( 
.A(n_10261),
.Y(n_10986)
);

NAND2x1p5_ASAP7_75t_SL g10987 ( 
.A(n_10133),
.B(n_8413),
.Y(n_10987)
);

AND2x2_ASAP7_75t_L g10988 ( 
.A(n_10389),
.B(n_6528),
.Y(n_10988)
);

AOI22xp33_ASAP7_75t_L g10989 ( 
.A1(n_10357),
.A2(n_9805),
.B1(n_9815),
.B2(n_9822),
.Y(n_10989)
);

INVxp67_ASAP7_75t_SL g10990 ( 
.A(n_10277),
.Y(n_10990)
);

BUFx2_ASAP7_75t_L g10991 ( 
.A(n_10232),
.Y(n_10991)
);

INVx2_ASAP7_75t_L g10992 ( 
.A(n_10293),
.Y(n_10992)
);

NAND2xp33_ASAP7_75t_R g10993 ( 
.A(n_10452),
.B(n_6266),
.Y(n_10993)
);

INVx3_ASAP7_75t_L g10994 ( 
.A(n_10232),
.Y(n_10994)
);

AND2x2_ASAP7_75t_L g10995 ( 
.A(n_10392),
.B(n_6528),
.Y(n_10995)
);

INVx2_ASAP7_75t_L g10996 ( 
.A(n_10170),
.Y(n_10996)
);

AND2x2_ASAP7_75t_L g10997 ( 
.A(n_10396),
.B(n_6584),
.Y(n_10997)
);

INVxp67_ASAP7_75t_L g10998 ( 
.A(n_10380),
.Y(n_10998)
);

AND2x4_ASAP7_75t_L g10999 ( 
.A(n_10301),
.B(n_9702),
.Y(n_10999)
);

INVx3_ASAP7_75t_L g11000 ( 
.A(n_10286),
.Y(n_11000)
);

INVx1_ASAP7_75t_SL g11001 ( 
.A(n_10403),
.Y(n_11001)
);

INVx1_ASAP7_75t_L g11002 ( 
.A(n_10319),
.Y(n_11002)
);

AND2x4_ASAP7_75t_L g11003 ( 
.A(n_10368),
.B(n_9703),
.Y(n_11003)
);

OR2x2_ASAP7_75t_L g11004 ( 
.A(n_10343),
.B(n_6852),
.Y(n_11004)
);

INVx1_ASAP7_75t_L g11005 ( 
.A(n_10327),
.Y(n_11005)
);

INVx2_ASAP7_75t_L g11006 ( 
.A(n_10173),
.Y(n_11006)
);

AND2x2_ASAP7_75t_L g11007 ( 
.A(n_10398),
.B(n_6584),
.Y(n_11007)
);

BUFx3_ASAP7_75t_L g11008 ( 
.A(n_10353),
.Y(n_11008)
);

INVx2_ASAP7_75t_L g11009 ( 
.A(n_10033),
.Y(n_11009)
);

INVx1_ASAP7_75t_L g11010 ( 
.A(n_10327),
.Y(n_11010)
);

OR2x2_ASAP7_75t_L g11011 ( 
.A(n_10128),
.B(n_6852),
.Y(n_11011)
);

BUFx6f_ASAP7_75t_L g11012 ( 
.A(n_10353),
.Y(n_11012)
);

NAND2xp5_ASAP7_75t_L g11013 ( 
.A(n_10041),
.B(n_8554),
.Y(n_11013)
);

AND2x2_ASAP7_75t_L g11014 ( 
.A(n_10429),
.B(n_10479),
.Y(n_11014)
);

AND2x4_ASAP7_75t_L g11015 ( 
.A(n_10286),
.B(n_10458),
.Y(n_11015)
);

OR2x2_ASAP7_75t_L g11016 ( 
.A(n_10138),
.B(n_6852),
.Y(n_11016)
);

INVx1_ASAP7_75t_L g11017 ( 
.A(n_10228),
.Y(n_11017)
);

INVx1_ASAP7_75t_L g11018 ( 
.A(n_10228),
.Y(n_11018)
);

INVx2_ASAP7_75t_L g11019 ( 
.A(n_10042),
.Y(n_11019)
);

INVx1_ASAP7_75t_L g11020 ( 
.A(n_10264),
.Y(n_11020)
);

AOI22xp33_ASAP7_75t_L g11021 ( 
.A1(n_10377),
.A2(n_8662),
.B1(n_9292),
.B2(n_8805),
.Y(n_11021)
);

INVx3_ASAP7_75t_L g11022 ( 
.A(n_10401),
.Y(n_11022)
);

AND2x2_ASAP7_75t_L g11023 ( 
.A(n_10360),
.B(n_10361),
.Y(n_11023)
);

INVx1_ASAP7_75t_SL g11024 ( 
.A(n_10237),
.Y(n_11024)
);

AND2x2_ASAP7_75t_L g11025 ( 
.A(n_10360),
.B(n_6584),
.Y(n_11025)
);

INVx1_ASAP7_75t_L g11026 ( 
.A(n_10264),
.Y(n_11026)
);

NAND2xp5_ASAP7_75t_L g11027 ( 
.A(n_10051),
.B(n_8564),
.Y(n_11027)
);

AND2x2_ASAP7_75t_L g11028 ( 
.A(n_10481),
.B(n_6584),
.Y(n_11028)
);

INVx2_ASAP7_75t_L g11029 ( 
.A(n_10530),
.Y(n_11029)
);

INVx1_ASAP7_75t_L g11030 ( 
.A(n_10525),
.Y(n_11030)
);

AND2x2_ASAP7_75t_L g11031 ( 
.A(n_10535),
.B(n_10397),
.Y(n_11031)
);

NAND2xp5_ASAP7_75t_L g11032 ( 
.A(n_10614),
.B(n_10411),
.Y(n_11032)
);

AND2x2_ASAP7_75t_L g11033 ( 
.A(n_10624),
.B(n_10363),
.Y(n_11033)
);

INVx2_ASAP7_75t_L g11034 ( 
.A(n_11015),
.Y(n_11034)
);

BUFx2_ASAP7_75t_L g11035 ( 
.A(n_10532),
.Y(n_11035)
);

INVx1_ASAP7_75t_L g11036 ( 
.A(n_10508),
.Y(n_11036)
);

INVx1_ASAP7_75t_L g11037 ( 
.A(n_10531),
.Y(n_11037)
);

AND2x2_ASAP7_75t_L g11038 ( 
.A(n_11015),
.B(n_10364),
.Y(n_11038)
);

INVx1_ASAP7_75t_L g11039 ( 
.A(n_10543),
.Y(n_11039)
);

INVxp67_ASAP7_75t_SL g11040 ( 
.A(n_10580),
.Y(n_11040)
);

INVx1_ASAP7_75t_L g11041 ( 
.A(n_10562),
.Y(n_11041)
);

INVx2_ASAP7_75t_L g11042 ( 
.A(n_11012),
.Y(n_11042)
);

INVx2_ASAP7_75t_L g11043 ( 
.A(n_11012),
.Y(n_11043)
);

INVx1_ASAP7_75t_L g11044 ( 
.A(n_10606),
.Y(n_11044)
);

BUFx2_ASAP7_75t_L g11045 ( 
.A(n_10749),
.Y(n_11045)
);

INVx2_ASAP7_75t_L g11046 ( 
.A(n_11012),
.Y(n_11046)
);

AND2x2_ASAP7_75t_L g11047 ( 
.A(n_10607),
.B(n_10460),
.Y(n_11047)
);

AND2x2_ASAP7_75t_L g11048 ( 
.A(n_10548),
.B(n_10842),
.Y(n_11048)
);

INVx2_ASAP7_75t_L g11049 ( 
.A(n_10731),
.Y(n_11049)
);

AND2x2_ASAP7_75t_L g11050 ( 
.A(n_10673),
.B(n_10462),
.Y(n_11050)
);

AND2x2_ASAP7_75t_L g11051 ( 
.A(n_10679),
.B(n_10441),
.Y(n_11051)
);

INVx1_ASAP7_75t_L g11052 ( 
.A(n_10613),
.Y(n_11052)
);

OR2x2_ASAP7_75t_L g11053 ( 
.A(n_11001),
.B(n_10184),
.Y(n_11053)
);

NAND2xp5_ASAP7_75t_L g11054 ( 
.A(n_10582),
.B(n_10414),
.Y(n_11054)
);

AND2x2_ASAP7_75t_L g11055 ( 
.A(n_10962),
.B(n_10214),
.Y(n_11055)
);

BUFx6f_ASAP7_75t_L g11056 ( 
.A(n_10495),
.Y(n_11056)
);

NAND2xp5_ASAP7_75t_L g11057 ( 
.A(n_10675),
.B(n_10459),
.Y(n_11057)
);

OR2x2_ASAP7_75t_L g11058 ( 
.A(n_11024),
.B(n_10355),
.Y(n_11058)
);

INVx2_ASAP7_75t_L g11059 ( 
.A(n_10937),
.Y(n_11059)
);

INVx1_ASAP7_75t_L g11060 ( 
.A(n_10972),
.Y(n_11060)
);

INVx5_ASAP7_75t_L g11061 ( 
.A(n_10495),
.Y(n_11061)
);

BUFx2_ASAP7_75t_L g11062 ( 
.A(n_10810),
.Y(n_11062)
);

AND2x2_ASAP7_75t_L g11063 ( 
.A(n_10704),
.B(n_10175),
.Y(n_11063)
);

INVx1_ASAP7_75t_L g11064 ( 
.A(n_10488),
.Y(n_11064)
);

AND2x2_ASAP7_75t_L g11065 ( 
.A(n_10623),
.B(n_10182),
.Y(n_11065)
);

INVx1_ASAP7_75t_L g11066 ( 
.A(n_10488),
.Y(n_11066)
);

AND2x2_ASAP7_75t_L g11067 ( 
.A(n_10504),
.B(n_10185),
.Y(n_11067)
);

AO21x2_ASAP7_75t_L g11068 ( 
.A1(n_10763),
.A2(n_10395),
.B(n_10044),
.Y(n_11068)
);

HB1xp67_ASAP7_75t_L g11069 ( 
.A(n_10919),
.Y(n_11069)
);

INVx4_ASAP7_75t_L g11070 ( 
.A(n_10495),
.Y(n_11070)
);

INVx1_ASAP7_75t_L g11071 ( 
.A(n_10492),
.Y(n_11071)
);

NAND2x1_ASAP7_75t_L g11072 ( 
.A(n_11022),
.B(n_10628),
.Y(n_11072)
);

AND2x2_ASAP7_75t_L g11073 ( 
.A(n_10513),
.B(n_10187),
.Y(n_11073)
);

AND2x2_ASAP7_75t_L g11074 ( 
.A(n_10702),
.B(n_10193),
.Y(n_11074)
);

HB1xp67_ASAP7_75t_L g11075 ( 
.A(n_10926),
.Y(n_11075)
);

HB1xp67_ASAP7_75t_L g11076 ( 
.A(n_10948),
.Y(n_11076)
);

INVx2_ASAP7_75t_SL g11077 ( 
.A(n_10546),
.Y(n_11077)
);

AOI22xp33_ASAP7_75t_L g11078 ( 
.A1(n_10510),
.A2(n_10395),
.B1(n_10399),
.B2(n_10404),
.Y(n_11078)
);

HB1xp67_ASAP7_75t_L g11079 ( 
.A(n_10819),
.Y(n_11079)
);

AO21x2_ASAP7_75t_L g11080 ( 
.A1(n_10763),
.A2(n_10044),
.B(n_9910),
.Y(n_11080)
);

NAND2xp5_ASAP7_75t_L g11081 ( 
.A(n_10920),
.B(n_10961),
.Y(n_11081)
);

HB1xp67_ASAP7_75t_L g11082 ( 
.A(n_10833),
.Y(n_11082)
);

HB1xp67_ASAP7_75t_L g11083 ( 
.A(n_10644),
.Y(n_11083)
);

AND2x2_ASAP7_75t_L g11084 ( 
.A(n_10551),
.B(n_10194),
.Y(n_11084)
);

INVx1_ASAP7_75t_L g11085 ( 
.A(n_10492),
.Y(n_11085)
);

AND2x2_ASAP7_75t_L g11086 ( 
.A(n_10522),
.B(n_10195),
.Y(n_11086)
);

INVx2_ASAP7_75t_L g11087 ( 
.A(n_10937),
.Y(n_11087)
);

AND2x2_ASAP7_75t_L g11088 ( 
.A(n_10529),
.B(n_10198),
.Y(n_11088)
);

NAND3xp33_ASAP7_75t_SL g11089 ( 
.A(n_10955),
.B(n_10248),
.C(n_10387),
.Y(n_11089)
);

AND2x4_ASAP7_75t_L g11090 ( 
.A(n_10601),
.B(n_10200),
.Y(n_11090)
);

OR2x2_ASAP7_75t_L g11091 ( 
.A(n_10695),
.B(n_10355),
.Y(n_11091)
);

INVx1_ASAP7_75t_L g11092 ( 
.A(n_10579),
.Y(n_11092)
);

HB1xp67_ASAP7_75t_L g11093 ( 
.A(n_10646),
.Y(n_11093)
);

INVx1_ASAP7_75t_L g11094 ( 
.A(n_10587),
.Y(n_11094)
);

INVxp67_ASAP7_75t_L g11095 ( 
.A(n_10554),
.Y(n_11095)
);

AND2x2_ASAP7_75t_L g11096 ( 
.A(n_10583),
.B(n_10465),
.Y(n_11096)
);

AND2x2_ASAP7_75t_SL g11097 ( 
.A(n_10835),
.B(n_10428),
.Y(n_11097)
);

OR2x6_ASAP7_75t_L g11098 ( 
.A(n_10565),
.B(n_10314),
.Y(n_11098)
);

AND2x2_ASAP7_75t_L g11099 ( 
.A(n_10734),
.B(n_10465),
.Y(n_11099)
);

AND2x2_ASAP7_75t_L g11100 ( 
.A(n_10660),
.B(n_10474),
.Y(n_11100)
);

AND2x2_ASAP7_75t_L g11101 ( 
.A(n_10661),
.B(n_10063),
.Y(n_11101)
);

OR2x6_ASAP7_75t_L g11102 ( 
.A(n_10861),
.B(n_10595),
.Y(n_11102)
);

INVx1_ASAP7_75t_SL g11103 ( 
.A(n_10796),
.Y(n_11103)
);

NAND2xp5_ASAP7_75t_L g11104 ( 
.A(n_11008),
.B(n_10990),
.Y(n_11104)
);

OR2x2_ASAP7_75t_L g11105 ( 
.A(n_10964),
.B(n_10025),
.Y(n_11105)
);

AOI22xp33_ASAP7_75t_L g11106 ( 
.A1(n_10913),
.A2(n_10413),
.B1(n_10422),
.B2(n_10366),
.Y(n_11106)
);

INVx1_ASAP7_75t_L g11107 ( 
.A(n_10590),
.Y(n_11107)
);

INVx2_ASAP7_75t_L g11108 ( 
.A(n_10659),
.Y(n_11108)
);

BUFx3_ASAP7_75t_L g11109 ( 
.A(n_10917),
.Y(n_11109)
);

INVx2_ASAP7_75t_L g11110 ( 
.A(n_10659),
.Y(n_11110)
);

NAND2xp5_ASAP7_75t_L g11111 ( 
.A(n_10716),
.B(n_10151),
.Y(n_11111)
);

AND2x4_ASAP7_75t_L g11112 ( 
.A(n_10601),
.B(n_10070),
.Y(n_11112)
);

AND2x2_ASAP7_75t_L g11113 ( 
.A(n_10982),
.B(n_10076),
.Y(n_11113)
);

AND2x2_ASAP7_75t_L g11114 ( 
.A(n_10658),
.B(n_10078),
.Y(n_11114)
);

INVx1_ASAP7_75t_L g11115 ( 
.A(n_10593),
.Y(n_11115)
);

INVx2_ASAP7_75t_L g11116 ( 
.A(n_10790),
.Y(n_11116)
);

AND2x2_ASAP7_75t_L g11117 ( 
.A(n_10567),
.B(n_10088),
.Y(n_11117)
);

INVx2_ASAP7_75t_L g11118 ( 
.A(n_10790),
.Y(n_11118)
);

AND2x2_ASAP7_75t_L g11119 ( 
.A(n_10733),
.B(n_10094),
.Y(n_11119)
);

INVx2_ASAP7_75t_L g11120 ( 
.A(n_10736),
.Y(n_11120)
);

BUFx2_ASAP7_75t_L g11121 ( 
.A(n_10852),
.Y(n_11121)
);

OAI221xp5_ASAP7_75t_L g11122 ( 
.A1(n_10486),
.A2(n_10440),
.B1(n_10082),
.B2(n_10468),
.C(n_10149),
.Y(n_11122)
);

INVx2_ASAP7_75t_L g11123 ( 
.A(n_10850),
.Y(n_11123)
);

AND2x4_ASAP7_75t_L g11124 ( 
.A(n_10701),
.B(n_10108),
.Y(n_11124)
);

AND2x2_ASAP7_75t_L g11125 ( 
.A(n_10770),
.B(n_10115),
.Y(n_11125)
);

INVx2_ASAP7_75t_L g11126 ( 
.A(n_10994),
.Y(n_11126)
);

NAND2xp5_ASAP7_75t_L g11127 ( 
.A(n_10779),
.B(n_10151),
.Y(n_11127)
);

INVx2_ASAP7_75t_L g11128 ( 
.A(n_10994),
.Y(n_11128)
);

INVx3_ASAP7_75t_L g11129 ( 
.A(n_10822),
.Y(n_11129)
);

HB1xp67_ASAP7_75t_L g11130 ( 
.A(n_10782),
.Y(n_11130)
);

AND2x2_ASAP7_75t_L g11131 ( 
.A(n_10636),
.B(n_10116),
.Y(n_11131)
);

OAI221xp5_ASAP7_75t_L g11132 ( 
.A1(n_10577),
.A2(n_10485),
.B1(n_10793),
.B2(n_10544),
.C(n_10691),
.Y(n_11132)
);

AND2x2_ASAP7_75t_L g11133 ( 
.A(n_10754),
.B(n_9935),
.Y(n_11133)
);

INVx3_ASAP7_75t_L g11134 ( 
.A(n_10822),
.Y(n_11134)
);

INVx1_ASAP7_75t_L g11135 ( 
.A(n_10598),
.Y(n_11135)
);

AND2x2_ASAP7_75t_L g11136 ( 
.A(n_10608),
.B(n_9935),
.Y(n_11136)
);

OR2x2_ASAP7_75t_L g11137 ( 
.A(n_10974),
.B(n_10263),
.Y(n_11137)
);

CKINVDCx5p33_ASAP7_75t_R g11138 ( 
.A(n_10663),
.Y(n_11138)
);

OR2x2_ASAP7_75t_L g11139 ( 
.A(n_10984),
.B(n_10470),
.Y(n_11139)
);

OR2x2_ASAP7_75t_L g11140 ( 
.A(n_10979),
.B(n_10197),
.Y(n_11140)
);

HB1xp67_ASAP7_75t_L g11141 ( 
.A(n_10942),
.Y(n_11141)
);

AND2x4_ASAP7_75t_L g11142 ( 
.A(n_10534),
.B(n_10027),
.Y(n_11142)
);

INVx1_ASAP7_75t_L g11143 ( 
.A(n_10604),
.Y(n_11143)
);

AND2x2_ASAP7_75t_L g11144 ( 
.A(n_10843),
.B(n_10634),
.Y(n_11144)
);

AND2x2_ASAP7_75t_L g11145 ( 
.A(n_10649),
.B(n_10402),
.Y(n_11145)
);

INVx2_ASAP7_75t_L g11146 ( 
.A(n_10866),
.Y(n_11146)
);

INVx1_ASAP7_75t_L g11147 ( 
.A(n_10605),
.Y(n_11147)
);

HB1xp67_ASAP7_75t_L g11148 ( 
.A(n_10946),
.Y(n_11148)
);

INVx1_ASAP7_75t_L g11149 ( 
.A(n_10618),
.Y(n_11149)
);

AND2x2_ASAP7_75t_L g11150 ( 
.A(n_10657),
.B(n_10416),
.Y(n_11150)
);

INVx1_ASAP7_75t_L g11151 ( 
.A(n_10620),
.Y(n_11151)
);

HB1xp67_ASAP7_75t_L g11152 ( 
.A(n_10949),
.Y(n_11152)
);

INVx2_ASAP7_75t_L g11153 ( 
.A(n_10866),
.Y(n_11153)
);

INVx1_ASAP7_75t_L g11154 ( 
.A(n_10625),
.Y(n_11154)
);

INVx1_ASAP7_75t_L g11155 ( 
.A(n_10627),
.Y(n_11155)
);

AND2x4_ASAP7_75t_L g11156 ( 
.A(n_10538),
.B(n_10563),
.Y(n_11156)
);

INVx5_ASAP7_75t_L g11157 ( 
.A(n_10569),
.Y(n_11157)
);

INVx2_ASAP7_75t_L g11158 ( 
.A(n_11000),
.Y(n_11158)
);

INVx3_ASAP7_75t_L g11159 ( 
.A(n_10847),
.Y(n_11159)
);

AND2x2_ASAP7_75t_L g11160 ( 
.A(n_10591),
.B(n_10436),
.Y(n_11160)
);

BUFx2_ASAP7_75t_L g11161 ( 
.A(n_10667),
.Y(n_11161)
);

INVx1_ASAP7_75t_L g11162 ( 
.A(n_10633),
.Y(n_11162)
);

AND2x2_ASAP7_75t_L g11163 ( 
.A(n_10629),
.B(n_10446),
.Y(n_11163)
);

NOR2x1_ASAP7_75t_L g11164 ( 
.A(n_10764),
.B(n_10471),
.Y(n_11164)
);

AND2x2_ASAP7_75t_L g11165 ( 
.A(n_10585),
.B(n_10448),
.Y(n_11165)
);

INVx2_ASAP7_75t_L g11166 ( 
.A(n_11000),
.Y(n_11166)
);

OR2x2_ASAP7_75t_L g11167 ( 
.A(n_10891),
.B(n_10035),
.Y(n_11167)
);

INVx2_ASAP7_75t_L g11168 ( 
.A(n_10896),
.Y(n_11168)
);

INVx3_ASAP7_75t_L g11169 ( 
.A(n_10847),
.Y(n_11169)
);

NAND2xp33_ASAP7_75t_SL g11170 ( 
.A(n_10921),
.B(n_10359),
.Y(n_11170)
);

HB1xp67_ASAP7_75t_L g11171 ( 
.A(n_10953),
.Y(n_11171)
);

INVx2_ASAP7_75t_L g11172 ( 
.A(n_10991),
.Y(n_11172)
);

INVx3_ASAP7_75t_L g11173 ( 
.A(n_10664),
.Y(n_11173)
);

INVx2_ASAP7_75t_L g11174 ( 
.A(n_10977),
.Y(n_11174)
);

INVx2_ASAP7_75t_L g11175 ( 
.A(n_10670),
.Y(n_11175)
);

OR2x2_ASAP7_75t_L g11176 ( 
.A(n_10915),
.B(n_10035),
.Y(n_11176)
);

INVx1_ASAP7_75t_SL g11177 ( 
.A(n_10748),
.Y(n_11177)
);

INVx2_ASAP7_75t_L g11178 ( 
.A(n_10615),
.Y(n_11178)
);

CKINVDCx20_ASAP7_75t_R g11179 ( 
.A(n_10603),
.Y(n_11179)
);

AND2x2_ASAP7_75t_L g11180 ( 
.A(n_10622),
.B(n_10449),
.Y(n_11180)
);

NOR2xp67_ASAP7_75t_L g11181 ( 
.A(n_10569),
.B(n_10381),
.Y(n_11181)
);

INVx2_ASAP7_75t_L g11182 ( 
.A(n_10615),
.Y(n_11182)
);

INVx1_ASAP7_75t_L g11183 ( 
.A(n_10765),
.Y(n_11183)
);

INVx1_ASAP7_75t_L g11184 ( 
.A(n_10765),
.Y(n_11184)
);

AND2x2_ASAP7_75t_L g11185 ( 
.A(n_10640),
.B(n_10450),
.Y(n_11185)
);

AND2x2_ASAP7_75t_L g11186 ( 
.A(n_10642),
.B(n_10457),
.Y(n_11186)
);

INVx1_ASAP7_75t_L g11187 ( 
.A(n_10767),
.Y(n_11187)
);

INVx2_ASAP7_75t_L g11188 ( 
.A(n_10876),
.Y(n_11188)
);

AND2x2_ASAP7_75t_L g11189 ( 
.A(n_10610),
.B(n_10461),
.Y(n_11189)
);

AOI22xp33_ASAP7_75t_L g11190 ( 
.A1(n_10533),
.A2(n_10216),
.B1(n_10434),
.B2(n_10432),
.Y(n_11190)
);

INVx1_ASAP7_75t_L g11191 ( 
.A(n_10767),
.Y(n_11191)
);

INVx1_ASAP7_75t_L g11192 ( 
.A(n_10641),
.Y(n_11192)
);

HB1xp67_ASAP7_75t_L g11193 ( 
.A(n_10756),
.Y(n_11193)
);

AND2x2_ASAP7_75t_L g11194 ( 
.A(n_10610),
.B(n_10463),
.Y(n_11194)
);

AND2x2_ASAP7_75t_L g11195 ( 
.A(n_10858),
.B(n_10469),
.Y(n_11195)
);

NAND2xp5_ASAP7_75t_L g11196 ( 
.A(n_10740),
.B(n_10155),
.Y(n_11196)
);

INVxp67_ASAP7_75t_L g11197 ( 
.A(n_10549),
.Y(n_11197)
);

INVx3_ASAP7_75t_L g11198 ( 
.A(n_10664),
.Y(n_11198)
);

HB1xp67_ASAP7_75t_L g11199 ( 
.A(n_10780),
.Y(n_11199)
);

AND2x2_ASAP7_75t_L g11200 ( 
.A(n_10859),
.B(n_10344),
.Y(n_11200)
);

AND2x2_ASAP7_75t_L g11201 ( 
.A(n_10496),
.B(n_10009),
.Y(n_11201)
);

AOI22xp5_ASAP7_75t_L g11202 ( 
.A1(n_10744),
.A2(n_10149),
.B1(n_10440),
.B2(n_10097),
.Y(n_11202)
);

AOI22xp5_ASAP7_75t_SL g11203 ( 
.A1(n_10998),
.A2(n_10155),
.B1(n_10359),
.B2(n_9910),
.Y(n_11203)
);

AOI22xp33_ASAP7_75t_L g11204 ( 
.A1(n_10912),
.A2(n_10439),
.B1(n_10444),
.B2(n_10433),
.Y(n_11204)
);

AND2x2_ASAP7_75t_L g11205 ( 
.A(n_10496),
.B(n_10009),
.Y(n_11205)
);

OAI22xp5_ASAP7_75t_L g11206 ( 
.A1(n_10602),
.A2(n_10381),
.B1(n_10298),
.B2(n_10384),
.Y(n_11206)
);

CKINVDCx6p67_ASAP7_75t_R g11207 ( 
.A(n_10569),
.Y(n_11207)
);

AND2x2_ASAP7_75t_L g11208 ( 
.A(n_10537),
.B(n_10009),
.Y(n_11208)
);

BUFx2_ASAP7_75t_L g11209 ( 
.A(n_10764),
.Y(n_11209)
);

AND2x4_ASAP7_75t_L g11210 ( 
.A(n_10839),
.B(n_10031),
.Y(n_11210)
);

INVx2_ASAP7_75t_L g11211 ( 
.A(n_10537),
.Y(n_11211)
);

INVx2_ASAP7_75t_L g11212 ( 
.A(n_10609),
.Y(n_11212)
);

INVx1_ASAP7_75t_L g11213 ( 
.A(n_10645),
.Y(n_11213)
);

NAND2xp33_ASAP7_75t_L g11214 ( 
.A(n_10527),
.B(n_10056),
.Y(n_11214)
);

INVx2_ASAP7_75t_SL g11215 ( 
.A(n_10917),
.Y(n_11215)
);

INVx2_ASAP7_75t_L g11216 ( 
.A(n_10609),
.Y(n_11216)
);

OAI22xp5_ASAP7_75t_L g11217 ( 
.A1(n_10813),
.A2(n_10298),
.B1(n_10438),
.B2(n_10466),
.Y(n_11217)
);

AOI22xp33_ASAP7_75t_L g11218 ( 
.A1(n_11021),
.A2(n_10420),
.B1(n_10478),
.B2(n_10477),
.Y(n_11218)
);

INVx1_ASAP7_75t_L g11219 ( 
.A(n_10728),
.Y(n_11219)
);

INVx2_ASAP7_75t_L g11220 ( 
.A(n_10588),
.Y(n_11220)
);

BUFx6f_ASAP7_75t_L g11221 ( 
.A(n_10708),
.Y(n_11221)
);

HB1xp67_ASAP7_75t_L g11222 ( 
.A(n_10668),
.Y(n_11222)
);

INVx2_ASAP7_75t_L g11223 ( 
.A(n_10708),
.Y(n_11223)
);

NAND2xp5_ASAP7_75t_L g11224 ( 
.A(n_10596),
.B(n_10475),
.Y(n_11224)
);

NOR2x1_ASAP7_75t_L g11225 ( 
.A(n_11022),
.B(n_10471),
.Y(n_11225)
);

INVxp67_ASAP7_75t_SL g11226 ( 
.A(n_10945),
.Y(n_11226)
);

HB1xp67_ASAP7_75t_L g11227 ( 
.A(n_10545),
.Y(n_11227)
);

AND2x4_ASAP7_75t_L g11228 ( 
.A(n_10787),
.B(n_10045),
.Y(n_11228)
);

OAI221xp5_ASAP7_75t_L g11229 ( 
.A1(n_10637),
.A2(n_10082),
.B1(n_10303),
.B2(n_9894),
.C(n_10230),
.Y(n_11229)
);

HB1xp67_ASAP7_75t_L g11230 ( 
.A(n_10547),
.Y(n_11230)
);

AND2x2_ASAP7_75t_L g11231 ( 
.A(n_10688),
.B(n_10417),
.Y(n_11231)
);

NAND2xp5_ASAP7_75t_L g11232 ( 
.A(n_10838),
.B(n_10239),
.Y(n_11232)
);

INVx1_ASAP7_75t_L g11233 ( 
.A(n_10728),
.Y(n_11233)
);

INVx1_ASAP7_75t_L g11234 ( 
.A(n_10556),
.Y(n_11234)
);

AND2x4_ASAP7_75t_L g11235 ( 
.A(n_10671),
.B(n_10049),
.Y(n_11235)
);

INVx1_ASAP7_75t_L g11236 ( 
.A(n_10559),
.Y(n_11236)
);

OAI211xp5_ASAP7_75t_SL g11237 ( 
.A1(n_10574),
.A2(n_10387),
.B(n_10316),
.C(n_10230),
.Y(n_11237)
);

INVxp67_ASAP7_75t_SL g11238 ( 
.A(n_10894),
.Y(n_11238)
);

OR2x2_ASAP7_75t_L g11239 ( 
.A(n_10987),
.B(n_10239),
.Y(n_11239)
);

AND2x4_ASAP7_75t_L g11240 ( 
.A(n_10671),
.B(n_10058),
.Y(n_11240)
);

NAND2xp5_ASAP7_75t_L g11241 ( 
.A(n_10823),
.B(n_9894),
.Y(n_11241)
);

INVx2_ASAP7_75t_L g11242 ( 
.A(n_10708),
.Y(n_11242)
);

INVx1_ASAP7_75t_SL g11243 ( 
.A(n_10867),
.Y(n_11243)
);

INVx3_ASAP7_75t_L g11244 ( 
.A(n_10638),
.Y(n_11244)
);

INVx2_ASAP7_75t_L g11245 ( 
.A(n_10621),
.Y(n_11245)
);

INVx2_ASAP7_75t_L g11246 ( 
.A(n_10621),
.Y(n_11246)
);

INVx1_ASAP7_75t_L g11247 ( 
.A(n_10561),
.Y(n_11247)
);

OR2x2_ASAP7_75t_L g11248 ( 
.A(n_10497),
.B(n_10447),
.Y(n_11248)
);

OR2x6_ASAP7_75t_L g11249 ( 
.A(n_10490),
.B(n_10352),
.Y(n_11249)
);

INVx4_ASAP7_75t_L g11250 ( 
.A(n_10978),
.Y(n_11250)
);

AND2x2_ASAP7_75t_L g11251 ( 
.A(n_10491),
.B(n_10050),
.Y(n_11251)
);

INVx2_ASAP7_75t_L g11252 ( 
.A(n_10540),
.Y(n_11252)
);

AND2x2_ASAP7_75t_L g11253 ( 
.A(n_10501),
.B(n_10209),
.Y(n_11253)
);

OR2x2_ASAP7_75t_L g11254 ( 
.A(n_10489),
.B(n_10056),
.Y(n_11254)
);

BUFx3_ASAP7_75t_L g11255 ( 
.A(n_10632),
.Y(n_11255)
);

INVx1_ASAP7_75t_L g11256 ( 
.A(n_10566),
.Y(n_11256)
);

INVx1_ASAP7_75t_L g11257 ( 
.A(n_10631),
.Y(n_11257)
);

INVx3_ASAP7_75t_L g11258 ( 
.A(n_10638),
.Y(n_11258)
);

HB1xp67_ASAP7_75t_L g11259 ( 
.A(n_10712),
.Y(n_11259)
);

AND2x2_ASAP7_75t_L g11260 ( 
.A(n_10934),
.B(n_10201),
.Y(n_11260)
);

INVx4_ASAP7_75t_L g11261 ( 
.A(n_10978),
.Y(n_11261)
);

OR2x6_ASAP7_75t_L g11262 ( 
.A(n_10498),
.B(n_10365),
.Y(n_11262)
);

OR2x2_ASAP7_75t_L g11263 ( 
.A(n_10992),
.B(n_10103),
.Y(n_11263)
);

INVx1_ASAP7_75t_L g11264 ( 
.A(n_10503),
.Y(n_11264)
);

AND2x4_ASAP7_75t_L g11265 ( 
.A(n_10506),
.B(n_10059),
.Y(n_11265)
);

AND2x2_ASAP7_75t_L g11266 ( 
.A(n_10619),
.B(n_10205),
.Y(n_11266)
);

INVx1_ASAP7_75t_L g11267 ( 
.A(n_10503),
.Y(n_11267)
);

INVx2_ASAP7_75t_L g11268 ( 
.A(n_10555),
.Y(n_11268)
);

AND2x2_ASAP7_75t_L g11269 ( 
.A(n_10568),
.B(n_10097),
.Y(n_11269)
);

NOR2xp33_ASAP7_75t_SL g11270 ( 
.A(n_10666),
.B(n_7234),
.Y(n_11270)
);

INVx1_ASAP7_75t_L g11271 ( 
.A(n_10511),
.Y(n_11271)
);

BUFx3_ASAP7_75t_L g11272 ( 
.A(n_10785),
.Y(n_11272)
);

INVx1_ASAP7_75t_L g11273 ( 
.A(n_10511),
.Y(n_11273)
);

AOI221xp5_ASAP7_75t_L g11274 ( 
.A1(n_11005),
.A2(n_10192),
.B1(n_10390),
.B2(n_10415),
.C(n_10135),
.Y(n_11274)
);

BUFx2_ASAP7_75t_L g11275 ( 
.A(n_10745),
.Y(n_11275)
);

AND2x2_ASAP7_75t_L g11276 ( 
.A(n_10573),
.B(n_10064),
.Y(n_11276)
);

INVx3_ASAP7_75t_L g11277 ( 
.A(n_10555),
.Y(n_11277)
);

INVx1_ASAP7_75t_L g11278 ( 
.A(n_10512),
.Y(n_11278)
);

NAND2xp5_ASAP7_75t_L g11279 ( 
.A(n_10739),
.B(n_10103),
.Y(n_11279)
);

INVx1_ASAP7_75t_L g11280 ( 
.A(n_10512),
.Y(n_11280)
);

AND2x2_ASAP7_75t_L g11281 ( 
.A(n_10969),
.B(n_10519),
.Y(n_11281)
);

AND2x4_ASAP7_75t_L g11282 ( 
.A(n_10560),
.B(n_10066),
.Y(n_11282)
);

INVx2_ASAP7_75t_SL g11283 ( 
.A(n_10976),
.Y(n_11283)
);

AND2x4_ASAP7_75t_L g11284 ( 
.A(n_10571),
.B(n_10068),
.Y(n_11284)
);

AND2x2_ASAP7_75t_L g11285 ( 
.A(n_10895),
.B(n_10069),
.Y(n_11285)
);

INVx1_ASAP7_75t_L g11286 ( 
.A(n_10515),
.Y(n_11286)
);

OR2x2_ASAP7_75t_L g11287 ( 
.A(n_10651),
.B(n_10729),
.Y(n_11287)
);

AND2x4_ASAP7_75t_L g11288 ( 
.A(n_10572),
.B(n_10073),
.Y(n_11288)
);

AND2x4_ASAP7_75t_L g11289 ( 
.A(n_10578),
.B(n_10592),
.Y(n_11289)
);

INVx1_ASAP7_75t_L g11290 ( 
.A(n_10515),
.Y(n_11290)
);

INVx1_ASAP7_75t_L g11291 ( 
.A(n_10821),
.Y(n_11291)
);

INVxp67_ASAP7_75t_SL g11292 ( 
.A(n_10894),
.Y(n_11292)
);

INVx1_ASAP7_75t_L g11293 ( 
.A(n_10775),
.Y(n_11293)
);

INVx2_ASAP7_75t_L g11294 ( 
.A(n_10581),
.Y(n_11294)
);

INVx2_ASAP7_75t_SL g11295 ( 
.A(n_10581),
.Y(n_11295)
);

AND2x2_ASAP7_75t_L g11296 ( 
.A(n_10576),
.B(n_10077),
.Y(n_11296)
);

INVx1_ASAP7_75t_L g11297 ( 
.A(n_10775),
.Y(n_11297)
);

AND2x2_ASAP7_75t_L g11298 ( 
.A(n_10951),
.B(n_10079),
.Y(n_11298)
);

AND2x2_ASAP7_75t_L g11299 ( 
.A(n_10635),
.B(n_10084),
.Y(n_11299)
);

INVx2_ASAP7_75t_L g11300 ( 
.A(n_10841),
.Y(n_11300)
);

INVx1_ASAP7_75t_L g11301 ( 
.A(n_10778),
.Y(n_11301)
);

OR2x2_ASAP7_75t_L g11302 ( 
.A(n_10650),
.B(n_10454),
.Y(n_11302)
);

INVx2_ASAP7_75t_L g11303 ( 
.A(n_10841),
.Y(n_11303)
);

INVx1_ASAP7_75t_L g11304 ( 
.A(n_10778),
.Y(n_11304)
);

OR2x6_ASAP7_75t_L g11305 ( 
.A(n_10594),
.B(n_10372),
.Y(n_11305)
);

AOI22xp33_ASAP7_75t_SL g11306 ( 
.A1(n_10536),
.A2(n_10192),
.B1(n_10466),
.B2(n_10135),
.Y(n_11306)
);

INVx2_ASAP7_75t_L g11307 ( 
.A(n_10552),
.Y(n_11307)
);

NAND2xp5_ASAP7_75t_L g11308 ( 
.A(n_10694),
.B(n_10415),
.Y(n_11308)
);

AND2x2_ASAP7_75t_L g11309 ( 
.A(n_10611),
.B(n_10093),
.Y(n_11309)
);

INVx1_ASAP7_75t_L g11310 ( 
.A(n_10907),
.Y(n_11310)
);

BUFx2_ASAP7_75t_L g11311 ( 
.A(n_10745),
.Y(n_11311)
);

BUFx3_ASAP7_75t_L g11312 ( 
.A(n_10678),
.Y(n_11312)
);

OR2x2_ASAP7_75t_L g11313 ( 
.A(n_10967),
.B(n_10454),
.Y(n_11313)
);

INVx1_ASAP7_75t_L g11314 ( 
.A(n_10907),
.Y(n_11314)
);

INVx1_ASAP7_75t_L g11315 ( 
.A(n_11002),
.Y(n_11315)
);

INVx2_ASAP7_75t_L g11316 ( 
.A(n_10507),
.Y(n_11316)
);

INVx2_ASAP7_75t_L g11317 ( 
.A(n_10557),
.Y(n_11317)
);

INVx1_ASAP7_75t_SL g11318 ( 
.A(n_11014),
.Y(n_11318)
);

INVx1_ASAP7_75t_L g11319 ( 
.A(n_11002),
.Y(n_11319)
);

INVx1_ASAP7_75t_L g11320 ( 
.A(n_10986),
.Y(n_11320)
);

INVx1_ASAP7_75t_L g11321 ( 
.A(n_10968),
.Y(n_11321)
);

AND2x2_ASAP7_75t_L g11322 ( 
.A(n_10612),
.B(n_10099),
.Y(n_11322)
);

BUFx2_ASAP7_75t_L g11323 ( 
.A(n_10746),
.Y(n_11323)
);

AND2x2_ASAP7_75t_L g11324 ( 
.A(n_10762),
.B(n_10101),
.Y(n_11324)
);

INVx1_ASAP7_75t_L g11325 ( 
.A(n_10981),
.Y(n_11325)
);

INVx1_ASAP7_75t_L g11326 ( 
.A(n_10983),
.Y(n_11326)
);

HB1xp67_ASAP7_75t_L g11327 ( 
.A(n_10857),
.Y(n_11327)
);

NAND2xp5_ASAP7_75t_L g11328 ( 
.A(n_10925),
.B(n_10303),
.Y(n_11328)
);

HB1xp67_ASAP7_75t_L g11329 ( 
.A(n_10517),
.Y(n_11329)
);

INVx1_ASAP7_75t_L g11330 ( 
.A(n_10539),
.Y(n_11330)
);

AND2x4_ASAP7_75t_L g11331 ( 
.A(n_10586),
.B(n_10102),
.Y(n_11331)
);

INVx1_ASAP7_75t_L g11332 ( 
.A(n_10541),
.Y(n_11332)
);

NOR2xp33_ASAP7_75t_R g11333 ( 
.A(n_10985),
.B(n_8054),
.Y(n_11333)
);

AND2x2_ASAP7_75t_L g11334 ( 
.A(n_10766),
.B(n_10106),
.Y(n_11334)
);

NAND2xp5_ASAP7_75t_L g11335 ( 
.A(n_10929),
.B(n_10931),
.Y(n_11335)
);

INVx3_ASAP7_75t_SL g11336 ( 
.A(n_10973),
.Y(n_11336)
);

INVx1_ASAP7_75t_L g11337 ( 
.A(n_10795),
.Y(n_11337)
);

HB1xp67_ASAP7_75t_L g11338 ( 
.A(n_10723),
.Y(n_11338)
);

AND2x2_ASAP7_75t_L g11339 ( 
.A(n_10684),
.B(n_10109),
.Y(n_11339)
);

INVx2_ASAP7_75t_L g11340 ( 
.A(n_10500),
.Y(n_11340)
);

NAND2xp5_ASAP7_75t_L g11341 ( 
.A(n_10936),
.B(n_10890),
.Y(n_11341)
);

INVx1_ASAP7_75t_L g11342 ( 
.A(n_10795),
.Y(n_11342)
);

INVx2_ASAP7_75t_L g11343 ( 
.A(n_10958),
.Y(n_11343)
);

HB1xp67_ASAP7_75t_L g11344 ( 
.A(n_10630),
.Y(n_11344)
);

NAND2xp5_ASAP7_75t_L g11345 ( 
.A(n_10706),
.B(n_10110),
.Y(n_11345)
);

INVx1_ASAP7_75t_L g11346 ( 
.A(n_10516),
.Y(n_11346)
);

AND2x2_ASAP7_75t_L g11347 ( 
.A(n_11023),
.B(n_10892),
.Y(n_11347)
);

AND2x4_ASAP7_75t_L g11348 ( 
.A(n_10586),
.B(n_10118),
.Y(n_11348)
);

INVx1_ASAP7_75t_L g11349 ( 
.A(n_10516),
.Y(n_11349)
);

INVx1_ASAP7_75t_L g11350 ( 
.A(n_10520),
.Y(n_11350)
);

AND2x2_ASAP7_75t_L g11351 ( 
.A(n_10863),
.B(n_10119),
.Y(n_11351)
);

NAND2xp5_ASAP7_75t_L g11352 ( 
.A(n_10910),
.B(n_10121),
.Y(n_11352)
);

HB1xp67_ASAP7_75t_L g11353 ( 
.A(n_10639),
.Y(n_11353)
);

INVx1_ASAP7_75t_L g11354 ( 
.A(n_10520),
.Y(n_11354)
);

NAND2xp5_ASAP7_75t_L g11355 ( 
.A(n_10910),
.B(n_10122),
.Y(n_11355)
);

AO21x2_ASAP7_75t_L g11356 ( 
.A1(n_10493),
.A2(n_10499),
.B(n_10494),
.Y(n_11356)
);

OR2x2_ASAP7_75t_L g11357 ( 
.A(n_10725),
.B(n_10390),
.Y(n_11357)
);

INVx5_ASAP7_75t_L g11358 ( 
.A(n_10714),
.Y(n_11358)
);

OR2x2_ASAP7_75t_L g11359 ( 
.A(n_10831),
.B(n_10836),
.Y(n_11359)
);

INVx1_ASAP7_75t_L g11360 ( 
.A(n_10523),
.Y(n_11360)
);

INVx2_ASAP7_75t_L g11361 ( 
.A(n_10727),
.Y(n_11361)
);

AOI22xp33_ASAP7_75t_L g11362 ( 
.A1(n_11005),
.A2(n_11017),
.B1(n_11018),
.B2(n_11010),
.Y(n_11362)
);

AND2x2_ASAP7_75t_L g11363 ( 
.A(n_10617),
.B(n_10129),
.Y(n_11363)
);

INVx1_ASAP7_75t_L g11364 ( 
.A(n_10523),
.Y(n_11364)
);

INVx2_ASAP7_75t_L g11365 ( 
.A(n_10889),
.Y(n_11365)
);

BUFx3_ASAP7_75t_L g11366 ( 
.A(n_10680),
.Y(n_11366)
);

BUFx2_ASAP7_75t_L g11367 ( 
.A(n_10746),
.Y(n_11367)
);

INVx1_ASAP7_75t_L g11368 ( 
.A(n_10524),
.Y(n_11368)
);

INVx2_ASAP7_75t_L g11369 ( 
.A(n_10750),
.Y(n_11369)
);

INVx1_ASAP7_75t_L g11370 ( 
.A(n_10524),
.Y(n_11370)
);

AND2x2_ASAP7_75t_L g11371 ( 
.A(n_10617),
.B(n_10139),
.Y(n_11371)
);

NAND2xp5_ASAP7_75t_SL g11372 ( 
.A(n_10505),
.B(n_9636),
.Y(n_11372)
);

OR2x2_ASAP7_75t_L g11373 ( 
.A(n_10837),
.B(n_10291),
.Y(n_11373)
);

NOR2xp33_ASAP7_75t_L g11374 ( 
.A(n_10700),
.B(n_10140),
.Y(n_11374)
);

BUFx6f_ASAP7_75t_L g11375 ( 
.A(n_11010),
.Y(n_11375)
);

INVx1_ASAP7_75t_L g11376 ( 
.A(n_10732),
.Y(n_11376)
);

INVx1_ASAP7_75t_L g11377 ( 
.A(n_10732),
.Y(n_11377)
);

INVx2_ASAP7_75t_SL g11378 ( 
.A(n_10904),
.Y(n_11378)
);

OR2x2_ASAP7_75t_L g11379 ( 
.A(n_10653),
.B(n_10291),
.Y(n_11379)
);

OR2x2_ASAP7_75t_L g11380 ( 
.A(n_10656),
.B(n_10296),
.Y(n_11380)
);

AND2x2_ASAP7_75t_L g11381 ( 
.A(n_10799),
.B(n_10145),
.Y(n_11381)
);

AND2x2_ASAP7_75t_L g11382 ( 
.A(n_10801),
.B(n_10146),
.Y(n_11382)
);

AND2x2_ASAP7_75t_L g11383 ( 
.A(n_10803),
.B(n_10153),
.Y(n_11383)
);

INVx2_ASAP7_75t_L g11384 ( 
.A(n_10752),
.Y(n_11384)
);

INVx1_ASAP7_75t_L g11385 ( 
.A(n_10735),
.Y(n_11385)
);

INVxp67_ASAP7_75t_SL g11386 ( 
.A(n_10662),
.Y(n_11386)
);

INVx3_ASAP7_75t_L g11387 ( 
.A(n_11003),
.Y(n_11387)
);

INVxp67_ASAP7_75t_SL g11388 ( 
.A(n_10509),
.Y(n_11388)
);

OR2x2_ASAP7_75t_L g11389 ( 
.A(n_10514),
.B(n_10296),
.Y(n_11389)
);

INVx3_ASAP7_75t_L g11390 ( 
.A(n_10597),
.Y(n_11390)
);

AND2x2_ASAP7_75t_L g11391 ( 
.A(n_10804),
.B(n_10154),
.Y(n_11391)
);

INVx2_ASAP7_75t_L g11392 ( 
.A(n_10753),
.Y(n_11392)
);

INVx3_ASAP7_75t_L g11393 ( 
.A(n_10769),
.Y(n_11393)
);

AND2x2_ASAP7_75t_L g11394 ( 
.A(n_10805),
.B(n_10158),
.Y(n_11394)
);

AND2x2_ASAP7_75t_L g11395 ( 
.A(n_10905),
.B(n_10166),
.Y(n_11395)
);

INVx2_ASAP7_75t_L g11396 ( 
.A(n_10760),
.Y(n_11396)
);

INVx2_ASAP7_75t_L g11397 ( 
.A(n_10751),
.Y(n_11397)
);

AO21x2_ASAP7_75t_L g11398 ( 
.A1(n_10493),
.A2(n_9990),
.B(n_10148),
.Y(n_11398)
);

AND2x2_ASAP7_75t_L g11399 ( 
.A(n_10906),
.B(n_10564),
.Y(n_11399)
);

NAND2xp5_ASAP7_75t_L g11400 ( 
.A(n_10814),
.B(n_10168),
.Y(n_11400)
);

NAND2xp5_ASAP7_75t_L g11401 ( 
.A(n_10737),
.B(n_10407),
.Y(n_11401)
);

INVx1_ASAP7_75t_L g11402 ( 
.A(n_10735),
.Y(n_11402)
);

NAND2xp5_ASAP7_75t_L g11403 ( 
.A(n_10783),
.B(n_10346),
.Y(n_11403)
);

INVx3_ASAP7_75t_L g11404 ( 
.A(n_10769),
.Y(n_11404)
);

INVx1_ASAP7_75t_L g11405 ( 
.A(n_10738),
.Y(n_11405)
);

AND2x2_ASAP7_75t_L g11406 ( 
.A(n_10742),
.B(n_10287),
.Y(n_11406)
);

HB1xp67_ASAP7_75t_L g11407 ( 
.A(n_10768),
.Y(n_11407)
);

INVx3_ASAP7_75t_L g11408 ( 
.A(n_10774),
.Y(n_11408)
);

BUFx6f_ASAP7_75t_L g11409 ( 
.A(n_11017),
.Y(n_11409)
);

INVx1_ASAP7_75t_L g11410 ( 
.A(n_10738),
.Y(n_11410)
);

INVx1_ASAP7_75t_L g11411 ( 
.A(n_10741),
.Y(n_11411)
);

OAI221xp5_ASAP7_75t_L g11412 ( 
.A1(n_10575),
.A2(n_10199),
.B1(n_10347),
.B2(n_10316),
.C(n_10309),
.Y(n_11412)
);

INVx3_ASAP7_75t_L g11413 ( 
.A(n_10774),
.Y(n_11413)
);

NAND2x1_ASAP7_75t_L g11414 ( 
.A(n_11018),
.B(n_10257),
.Y(n_11414)
);

NAND2xp5_ASAP7_75t_L g11415 ( 
.A(n_10784),
.B(n_10346),
.Y(n_11415)
);

AND2x2_ASAP7_75t_L g11416 ( 
.A(n_10717),
.B(n_10346),
.Y(n_11416)
);

AND2x2_ASAP7_75t_L g11417 ( 
.A(n_10721),
.B(n_10299),
.Y(n_11417)
);

OR2x2_ASAP7_75t_L g11418 ( 
.A(n_10528),
.B(n_9890),
.Y(n_11418)
);

INVx1_ASAP7_75t_L g11419 ( 
.A(n_10741),
.Y(n_11419)
);

INVx2_ASAP7_75t_L g11420 ( 
.A(n_10947),
.Y(n_11420)
);

AND2x2_ASAP7_75t_L g11421 ( 
.A(n_10726),
.B(n_10308),
.Y(n_11421)
);

AND2x2_ASAP7_75t_L g11422 ( 
.A(n_10918),
.B(n_10091),
.Y(n_11422)
);

OR2x2_ASAP7_75t_L g11423 ( 
.A(n_10807),
.B(n_9920),
.Y(n_11423)
);

AND2x2_ASAP7_75t_L g11424 ( 
.A(n_10761),
.B(n_10091),
.Y(n_11424)
);

AND2x2_ASAP7_75t_L g11425 ( 
.A(n_10773),
.B(n_10091),
.Y(n_11425)
);

INVx2_ASAP7_75t_SL g11426 ( 
.A(n_10715),
.Y(n_11426)
);

OR2x2_ASAP7_75t_L g11427 ( 
.A(n_10809),
.B(n_9948),
.Y(n_11427)
);

HB1xp67_ASAP7_75t_L g11428 ( 
.A(n_10768),
.Y(n_11428)
);

NAND2xp5_ASAP7_75t_SL g11429 ( 
.A(n_10724),
.B(n_9600),
.Y(n_11429)
);

INVx1_ASAP7_75t_L g11430 ( 
.A(n_10996),
.Y(n_11430)
);

INVx2_ASAP7_75t_L g11431 ( 
.A(n_10947),
.Y(n_11431)
);

INVx2_ASAP7_75t_L g11432 ( 
.A(n_10648),
.Y(n_11432)
);

INVx1_ASAP7_75t_L g11433 ( 
.A(n_11006),
.Y(n_11433)
);

AND2x2_ASAP7_75t_L g11434 ( 
.A(n_10777),
.B(n_10329),
.Y(n_11434)
);

NAND2xp5_ASAP7_75t_L g11435 ( 
.A(n_10935),
.B(n_10421),
.Y(n_11435)
);

AND2x2_ASAP7_75t_L g11436 ( 
.A(n_10975),
.B(n_10199),
.Y(n_11436)
);

HB1xp67_ASAP7_75t_L g11437 ( 
.A(n_10771),
.Y(n_11437)
);

AND2x2_ASAP7_75t_L g11438 ( 
.A(n_10710),
.B(n_9928),
.Y(n_11438)
);

AOI22xp33_ASAP7_75t_L g11439 ( 
.A1(n_11020),
.A2(n_10423),
.B1(n_10373),
.B2(n_10375),
.Y(n_11439)
);

AO21x2_ASAP7_75t_L g11440 ( 
.A1(n_10494),
.A2(n_10022),
.B(n_10014),
.Y(n_11440)
);

AND2x2_ASAP7_75t_L g11441 ( 
.A(n_10711),
.B(n_10258),
.Y(n_11441)
);

NAND2xp5_ASAP7_75t_L g11442 ( 
.A(n_11009),
.B(n_10430),
.Y(n_11442)
);

AND2x4_ASAP7_75t_L g11443 ( 
.A(n_10697),
.B(n_10285),
.Y(n_11443)
);

AND2x2_ASAP7_75t_L g11444 ( 
.A(n_10930),
.B(n_10999),
.Y(n_11444)
);

AO21x2_ASAP7_75t_L g11445 ( 
.A1(n_10499),
.A2(n_10309),
.B(n_10332),
.Y(n_11445)
);

AOI22xp33_ASAP7_75t_L g11446 ( 
.A1(n_11020),
.A2(n_10374),
.B1(n_10426),
.B2(n_10351),
.Y(n_11446)
);

INVx1_ASAP7_75t_L g11447 ( 
.A(n_10828),
.Y(n_11447)
);

INVx1_ASAP7_75t_L g11448 ( 
.A(n_10829),
.Y(n_11448)
);

INVxp67_ASAP7_75t_SL g11449 ( 
.A(n_10518),
.Y(n_11449)
);

AND2x2_ASAP7_75t_L g11450 ( 
.A(n_10999),
.B(n_10297),
.Y(n_11450)
);

AND2x2_ASAP7_75t_L g11451 ( 
.A(n_10816),
.B(n_10401),
.Y(n_11451)
);

INVx1_ASAP7_75t_L g11452 ( 
.A(n_10818),
.Y(n_11452)
);

INVx1_ASAP7_75t_L g11453 ( 
.A(n_10502),
.Y(n_11453)
);

INVx1_ASAP7_75t_L g11454 ( 
.A(n_10502),
.Y(n_11454)
);

HB1xp67_ASAP7_75t_L g11455 ( 
.A(n_10771),
.Y(n_11455)
);

INVx1_ASAP7_75t_L g11456 ( 
.A(n_10652),
.Y(n_11456)
);

OR2x2_ASAP7_75t_L g11457 ( 
.A(n_10840),
.B(n_10347),
.Y(n_11457)
);

AND2x2_ASAP7_75t_L g11458 ( 
.A(n_10832),
.B(n_8831),
.Y(n_11458)
);

INVx2_ASAP7_75t_L g11459 ( 
.A(n_10655),
.Y(n_11459)
);

AND2x2_ASAP7_75t_L g11460 ( 
.A(n_10834),
.B(n_8831),
.Y(n_11460)
);

AOI221xp5_ASAP7_75t_L g11461 ( 
.A1(n_11026),
.A2(n_10342),
.B1(n_10337),
.B2(n_10333),
.C(n_10382),
.Y(n_11461)
);

INVx1_ASAP7_75t_L g11462 ( 
.A(n_10677),
.Y(n_11462)
);

AND2x2_ASAP7_75t_L g11463 ( 
.A(n_10849),
.B(n_9663),
.Y(n_11463)
);

INVx1_ASAP7_75t_L g11464 ( 
.A(n_10584),
.Y(n_11464)
);

AND2x2_ASAP7_75t_L g11465 ( 
.A(n_10851),
.B(n_6584),
.Y(n_11465)
);

AOI221xp5_ASAP7_75t_L g11466 ( 
.A1(n_11026),
.A2(n_10382),
.B1(n_10376),
.B2(n_10345),
.C(n_10349),
.Y(n_11466)
);

INVx2_ASAP7_75t_L g11467 ( 
.A(n_10703),
.Y(n_11467)
);

AND2x2_ASAP7_75t_L g11468 ( 
.A(n_10853),
.B(n_6598),
.Y(n_11468)
);

INVx2_ASAP7_75t_L g11469 ( 
.A(n_10743),
.Y(n_11469)
);

INVx2_ASAP7_75t_L g11470 ( 
.A(n_10747),
.Y(n_11470)
);

AOI211xp5_ASAP7_75t_L g11471 ( 
.A1(n_10758),
.A2(n_9755),
.B(n_10382),
.C(n_9766),
.Y(n_11471)
);

NAND2xp5_ASAP7_75t_L g11472 ( 
.A(n_11019),
.B(n_10345),
.Y(n_11472)
);

OAI33xp33_ASAP7_75t_L g11473 ( 
.A1(n_10781),
.A2(n_10222),
.A3(n_10224),
.B1(n_10219),
.B2(n_10255),
.B3(n_10253),
.Y(n_11473)
);

INVxp67_ASAP7_75t_L g11474 ( 
.A(n_10815),
.Y(n_11474)
);

INVx1_ASAP7_75t_L g11475 ( 
.A(n_10599),
.Y(n_11475)
);

HB1xp67_ASAP7_75t_L g11476 ( 
.A(n_10870),
.Y(n_11476)
);

INVx1_ASAP7_75t_L g11477 ( 
.A(n_10860),
.Y(n_11477)
);

INVxp67_ASAP7_75t_L g11478 ( 
.A(n_10589),
.Y(n_11478)
);

INVx1_ASAP7_75t_L g11479 ( 
.A(n_10626),
.Y(n_11479)
);

OR2x2_ASAP7_75t_L g11480 ( 
.A(n_10802),
.B(n_10376),
.Y(n_11480)
);

INVx2_ASAP7_75t_L g11481 ( 
.A(n_10674),
.Y(n_11481)
);

OAI211xp5_ASAP7_75t_SL g11482 ( 
.A1(n_10722),
.A2(n_10167),
.B(n_8467),
.C(n_8475),
.Y(n_11482)
);

INVx1_ASAP7_75t_L g11483 ( 
.A(n_10856),
.Y(n_11483)
);

BUFx3_ASAP7_75t_L g11484 ( 
.A(n_10707),
.Y(n_11484)
);

BUFx2_ASAP7_75t_L g11485 ( 
.A(n_10692),
.Y(n_11485)
);

OR2x2_ASAP7_75t_L g11486 ( 
.A(n_10824),
.B(n_10394),
.Y(n_11486)
);

OR2x6_ASAP7_75t_L g11487 ( 
.A(n_10873),
.B(n_7647),
.Y(n_11487)
);

AND2x2_ASAP7_75t_L g11488 ( 
.A(n_10880),
.B(n_6598),
.Y(n_11488)
);

AND2x2_ASAP7_75t_L g11489 ( 
.A(n_10776),
.B(n_6598),
.Y(n_11489)
);

AND2x4_ASAP7_75t_L g11490 ( 
.A(n_10709),
.B(n_8456),
.Y(n_11490)
);

NAND2xp5_ASAP7_75t_L g11491 ( 
.A(n_10690),
.B(n_10336),
.Y(n_11491)
);

NAND2xp5_ASAP7_75t_SL g11492 ( 
.A(n_11003),
.B(n_9747),
.Y(n_11492)
);

HB1xp67_ASAP7_75t_L g11493 ( 
.A(n_10875),
.Y(n_11493)
);

AND2x4_ASAP7_75t_L g11494 ( 
.A(n_10820),
.B(n_8467),
.Y(n_11494)
);

NAND4xp25_ASAP7_75t_L g11495 ( 
.A(n_10550),
.B(n_8420),
.C(n_8421),
.D(n_8467),
.Y(n_11495)
);

INVxp67_ASAP7_75t_L g11496 ( 
.A(n_10487),
.Y(n_11496)
);

NOR2x1_ASAP7_75t_SL g11497 ( 
.A(n_10757),
.B(n_10259),
.Y(n_11497)
);

INVx2_ASAP7_75t_L g11498 ( 
.A(n_10676),
.Y(n_11498)
);

AND2x2_ASAP7_75t_L g11499 ( 
.A(n_10868),
.B(n_6598),
.Y(n_11499)
);

AND2x2_ASAP7_75t_L g11500 ( 
.A(n_10825),
.B(n_6598),
.Y(n_11500)
);

AND2x2_ASAP7_75t_L g11501 ( 
.A(n_10941),
.B(n_6642),
.Y(n_11501)
);

AND2x2_ASAP7_75t_L g11502 ( 
.A(n_10808),
.B(n_6642),
.Y(n_11502)
);

AND2x4_ASAP7_75t_L g11503 ( 
.A(n_10827),
.B(n_8475),
.Y(n_11503)
);

AND2x2_ASAP7_75t_L g11504 ( 
.A(n_10811),
.B(n_6642),
.Y(n_11504)
);

AND2x2_ASAP7_75t_L g11505 ( 
.A(n_11103),
.B(n_10789),
.Y(n_11505)
);

AND2x2_ASAP7_75t_L g11506 ( 
.A(n_11077),
.B(n_10798),
.Y(n_11506)
);

INVx1_ASAP7_75t_L g11507 ( 
.A(n_11069),
.Y(n_11507)
);

INVx2_ASAP7_75t_L g11508 ( 
.A(n_11277),
.Y(n_11508)
);

AND2x2_ASAP7_75t_L g11509 ( 
.A(n_11048),
.B(n_10772),
.Y(n_11509)
);

AND2x4_ASAP7_75t_L g11510 ( 
.A(n_11109),
.B(n_10888),
.Y(n_11510)
);

HB1xp67_ASAP7_75t_L g11511 ( 
.A(n_11072),
.Y(n_11511)
);

INVx1_ASAP7_75t_L g11512 ( 
.A(n_11075),
.Y(n_11512)
);

NAND2xp5_ASAP7_75t_L g11513 ( 
.A(n_11253),
.B(n_10928),
.Y(n_11513)
);

INVx2_ASAP7_75t_L g11514 ( 
.A(n_11277),
.Y(n_11514)
);

NAND2x1_ASAP7_75t_SL g11515 ( 
.A(n_11076),
.B(n_10830),
.Y(n_11515)
);

NAND2xp5_ASAP7_75t_L g11516 ( 
.A(n_11251),
.B(n_10932),
.Y(n_11516)
);

INVx2_ASAP7_75t_L g11517 ( 
.A(n_11387),
.Y(n_11517)
);

AND2x2_ASAP7_75t_L g11518 ( 
.A(n_11318),
.B(n_10897),
.Y(n_11518)
);

HB1xp67_ASAP7_75t_L g11519 ( 
.A(n_11072),
.Y(n_11519)
);

AND2x2_ASAP7_75t_L g11520 ( 
.A(n_11399),
.B(n_11102),
.Y(n_11520)
);

INVx1_ASAP7_75t_L g11521 ( 
.A(n_11356),
.Y(n_11521)
);

AND2x4_ASAP7_75t_SL g11522 ( 
.A(n_11031),
.B(n_10893),
.Y(n_11522)
);

INVx2_ASAP7_75t_L g11523 ( 
.A(n_11221),
.Y(n_11523)
);

INVxp67_ASAP7_75t_L g11524 ( 
.A(n_11238),
.Y(n_11524)
);

INVx1_ASAP7_75t_L g11525 ( 
.A(n_11222),
.Y(n_11525)
);

NAND2xp5_ASAP7_75t_L g11526 ( 
.A(n_11231),
.B(n_10845),
.Y(n_11526)
);

BUFx2_ASAP7_75t_L g11527 ( 
.A(n_11225),
.Y(n_11527)
);

INVx1_ASAP7_75t_L g11528 ( 
.A(n_11141),
.Y(n_11528)
);

INVx2_ASAP7_75t_L g11529 ( 
.A(n_11221),
.Y(n_11529)
);

AND2x2_ASAP7_75t_L g11530 ( 
.A(n_11102),
.B(n_10902),
.Y(n_11530)
);

INVx2_ASAP7_75t_L g11531 ( 
.A(n_11221),
.Y(n_11531)
);

NAND2xp5_ASAP7_75t_L g11532 ( 
.A(n_11097),
.B(n_10672),
.Y(n_11532)
);

NAND2xp5_ASAP7_75t_L g11533 ( 
.A(n_11386),
.B(n_10886),
.Y(n_11533)
);

INVx2_ASAP7_75t_L g11534 ( 
.A(n_11295),
.Y(n_11534)
);

INVx2_ASAP7_75t_L g11535 ( 
.A(n_11129),
.Y(n_11535)
);

INVx1_ASAP7_75t_L g11536 ( 
.A(n_11148),
.Y(n_11536)
);

NAND2xp5_ASAP7_75t_L g11537 ( 
.A(n_11131),
.B(n_10886),
.Y(n_11537)
);

AND2x4_ASAP7_75t_L g11538 ( 
.A(n_11215),
.B(n_10898),
.Y(n_11538)
);

AND2x2_ASAP7_75t_L g11539 ( 
.A(n_11339),
.B(n_11028),
.Y(n_11539)
);

AND2x2_ASAP7_75t_L g11540 ( 
.A(n_11299),
.B(n_11444),
.Y(n_11540)
);

AND2x4_ASAP7_75t_L g11541 ( 
.A(n_11059),
.B(n_10903),
.Y(n_11541)
);

AND2x4_ASAP7_75t_L g11542 ( 
.A(n_11087),
.B(n_10654),
.Y(n_11542)
);

INVx1_ASAP7_75t_L g11543 ( 
.A(n_11152),
.Y(n_11543)
);

CKINVDCx16_ASAP7_75t_R g11544 ( 
.A(n_11050),
.Y(n_11544)
);

AND2x2_ASAP7_75t_L g11545 ( 
.A(n_11144),
.B(n_10730),
.Y(n_11545)
);

AND2x4_ASAP7_75t_L g11546 ( 
.A(n_11034),
.B(n_10665),
.Y(n_11546)
);

INVx1_ASAP7_75t_L g11547 ( 
.A(n_11171),
.Y(n_11547)
);

INVx1_ASAP7_75t_L g11548 ( 
.A(n_11259),
.Y(n_11548)
);

BUFx3_ASAP7_75t_L g11549 ( 
.A(n_11138),
.Y(n_11549)
);

OR2x2_ASAP7_75t_L g11550 ( 
.A(n_11254),
.B(n_10643),
.Y(n_11550)
);

AND2x2_ASAP7_75t_L g11551 ( 
.A(n_11163),
.B(n_10882),
.Y(n_11551)
);

INVx1_ASAP7_75t_L g11552 ( 
.A(n_11327),
.Y(n_11552)
);

NAND2xp5_ASAP7_75t_L g11553 ( 
.A(n_11296),
.B(n_11117),
.Y(n_11553)
);

INVx2_ASAP7_75t_L g11554 ( 
.A(n_11129),
.Y(n_11554)
);

INVx1_ASAP7_75t_L g11555 ( 
.A(n_11199),
.Y(n_11555)
);

NAND2xp5_ASAP7_75t_L g11556 ( 
.A(n_11266),
.B(n_11156),
.Y(n_11556)
);

INVx1_ASAP7_75t_L g11557 ( 
.A(n_11161),
.Y(n_11557)
);

INVx2_ASAP7_75t_L g11558 ( 
.A(n_11134),
.Y(n_11558)
);

INVx1_ASAP7_75t_L g11559 ( 
.A(n_11161),
.Y(n_11559)
);

AND2x4_ASAP7_75t_L g11560 ( 
.A(n_11124),
.B(n_10669),
.Y(n_11560)
);

INVx1_ASAP7_75t_L g11561 ( 
.A(n_11035),
.Y(n_11561)
);

AND2x2_ASAP7_75t_L g11562 ( 
.A(n_11347),
.B(n_10911),
.Y(n_11562)
);

AND2x4_ASAP7_75t_SL g11563 ( 
.A(n_11047),
.B(n_10682),
.Y(n_11563)
);

INVx1_ASAP7_75t_L g11564 ( 
.A(n_11035),
.Y(n_11564)
);

INVx2_ASAP7_75t_L g11565 ( 
.A(n_11134),
.Y(n_11565)
);

AND2x4_ASAP7_75t_L g11566 ( 
.A(n_11124),
.B(n_10683),
.Y(n_11566)
);

OR2x2_ASAP7_75t_L g11567 ( 
.A(n_11053),
.B(n_10887),
.Y(n_11567)
);

INVx1_ASAP7_75t_L g11568 ( 
.A(n_11375),
.Y(n_11568)
);

OR2x2_ASAP7_75t_L g11569 ( 
.A(n_11248),
.B(n_10872),
.Y(n_11569)
);

BUFx2_ASAP7_75t_L g11570 ( 
.A(n_11068),
.Y(n_11570)
);

INVx1_ASAP7_75t_L g11571 ( 
.A(n_11375),
.Y(n_11571)
);

OR2x2_ASAP7_75t_L g11572 ( 
.A(n_11111),
.B(n_10884),
.Y(n_11572)
);

OR2x2_ASAP7_75t_L g11573 ( 
.A(n_11196),
.B(n_10686),
.Y(n_11573)
);

INVx2_ASAP7_75t_L g11574 ( 
.A(n_11159),
.Y(n_11574)
);

INVx2_ASAP7_75t_L g11575 ( 
.A(n_11159),
.Y(n_11575)
);

INVx1_ASAP7_75t_L g11576 ( 
.A(n_11375),
.Y(n_11576)
);

AND2x2_ASAP7_75t_L g11577 ( 
.A(n_11260),
.B(n_10923),
.Y(n_11577)
);

NOR2xp67_ASAP7_75t_L g11578 ( 
.A(n_11061),
.B(n_10689),
.Y(n_11578)
);

NAND2xp5_ASAP7_75t_L g11579 ( 
.A(n_11156),
.B(n_10553),
.Y(n_11579)
);

INVx1_ASAP7_75t_L g11580 ( 
.A(n_11409),
.Y(n_11580)
);

OR2x2_ASAP7_75t_L g11581 ( 
.A(n_11091),
.B(n_10687),
.Y(n_11581)
);

OR2x2_ASAP7_75t_L g11582 ( 
.A(n_11389),
.B(n_11357),
.Y(n_11582)
);

BUFx2_ASAP7_75t_L g11583 ( 
.A(n_11445),
.Y(n_11583)
);

AND2x4_ASAP7_75t_SL g11584 ( 
.A(n_11029),
.B(n_10693),
.Y(n_11584)
);

OR2x2_ASAP7_75t_L g11585 ( 
.A(n_11241),
.B(n_10681),
.Y(n_11585)
);

NAND2xp5_ASAP7_75t_L g11586 ( 
.A(n_11065),
.B(n_10826),
.Y(n_11586)
);

AND2x4_ASAP7_75t_L g11587 ( 
.A(n_11125),
.B(n_10696),
.Y(n_11587)
);

NAND2xp5_ASAP7_75t_L g11588 ( 
.A(n_11485),
.B(n_10848),
.Y(n_11588)
);

INVx1_ASAP7_75t_L g11589 ( 
.A(n_11409),
.Y(n_11589)
);

AND2x4_ASAP7_75t_L g11590 ( 
.A(n_11098),
.B(n_10699),
.Y(n_11590)
);

INVx2_ASAP7_75t_L g11591 ( 
.A(n_11169),
.Y(n_11591)
);

OR2x2_ASAP7_75t_L g11592 ( 
.A(n_11127),
.B(n_10844),
.Y(n_11592)
);

INVx1_ASAP7_75t_SL g11593 ( 
.A(n_11038),
.Y(n_11593)
);

OR2x2_ASAP7_75t_L g11594 ( 
.A(n_11232),
.B(n_10914),
.Y(n_11594)
);

AND2x2_ASAP7_75t_L g11595 ( 
.A(n_11336),
.B(n_10924),
.Y(n_11595)
);

INVx2_ASAP7_75t_L g11596 ( 
.A(n_11169),
.Y(n_11596)
);

NAND2xp5_ASAP7_75t_L g11597 ( 
.A(n_11485),
.B(n_10698),
.Y(n_11597)
);

AND2x2_ASAP7_75t_L g11598 ( 
.A(n_11165),
.B(n_11025),
.Y(n_11598)
);

AND2x2_ASAP7_75t_L g11599 ( 
.A(n_11033),
.B(n_10960),
.Y(n_11599)
);

OR2x2_ASAP7_75t_L g11600 ( 
.A(n_11287),
.B(n_10862),
.Y(n_11600)
);

INVx1_ASAP7_75t_L g11601 ( 
.A(n_11409),
.Y(n_11601)
);

AND2x2_ASAP7_75t_L g11602 ( 
.A(n_11130),
.B(n_10705),
.Y(n_11602)
);

INVx1_ASAP7_75t_L g11603 ( 
.A(n_11045),
.Y(n_11603)
);

AND2x2_ASAP7_75t_L g11604 ( 
.A(n_11160),
.B(n_10713),
.Y(n_11604)
);

NAND2xp5_ASAP7_75t_SL g11605 ( 
.A(n_11121),
.B(n_10542),
.Y(n_11605)
);

AND2x2_ASAP7_75t_L g11606 ( 
.A(n_11309),
.B(n_10718),
.Y(n_11606)
);

AND2x2_ASAP7_75t_L g11607 ( 
.A(n_11322),
.B(n_10755),
.Y(n_11607)
);

AND2x2_ASAP7_75t_L g11608 ( 
.A(n_11119),
.B(n_10759),
.Y(n_11608)
);

AND2x2_ASAP7_75t_L g11609 ( 
.A(n_11133),
.B(n_10988),
.Y(n_11609)
);

AND2x2_ASAP7_75t_L g11610 ( 
.A(n_11063),
.B(n_10995),
.Y(n_11610)
);

INVx1_ASAP7_75t_L g11611 ( 
.A(n_11045),
.Y(n_11611)
);

INVx1_ASAP7_75t_L g11612 ( 
.A(n_11062),
.Y(n_11612)
);

BUFx2_ASAP7_75t_L g11613 ( 
.A(n_11062),
.Y(n_11613)
);

INVx1_ASAP7_75t_L g11614 ( 
.A(n_11420),
.Y(n_11614)
);

INVx3_ASAP7_75t_L g11615 ( 
.A(n_11112),
.Y(n_11615)
);

INVx1_ASAP7_75t_L g11616 ( 
.A(n_11431),
.Y(n_11616)
);

AOI22xp33_ASAP7_75t_L g11617 ( 
.A1(n_11237),
.A2(n_10600),
.B1(n_10647),
.B2(n_10521),
.Y(n_11617)
);

NAND2xp5_ASAP7_75t_L g11618 ( 
.A(n_11040),
.B(n_10781),
.Y(n_11618)
);

NAND2xp33_ASAP7_75t_R g11619 ( 
.A(n_11121),
.B(n_10786),
.Y(n_11619)
);

INVx1_ASAP7_75t_L g11620 ( 
.A(n_11268),
.Y(n_11620)
);

AND2x2_ASAP7_75t_L g11621 ( 
.A(n_11406),
.B(n_10997),
.Y(n_11621)
);

AND2x2_ASAP7_75t_L g11622 ( 
.A(n_11074),
.B(n_11007),
.Y(n_11622)
);

INVxp67_ASAP7_75t_SL g11623 ( 
.A(n_11164),
.Y(n_11623)
);

AND2x2_ASAP7_75t_L g11624 ( 
.A(n_11101),
.B(n_10939),
.Y(n_11624)
);

NAND2xp5_ASAP7_75t_SL g11625 ( 
.A(n_11239),
.B(n_10877),
.Y(n_11625)
);

AND2x2_ASAP7_75t_L g11626 ( 
.A(n_11276),
.B(n_10940),
.Y(n_11626)
);

INVx1_ASAP7_75t_L g11627 ( 
.A(n_11294),
.Y(n_11627)
);

NAND2xp5_ASAP7_75t_L g11628 ( 
.A(n_11226),
.B(n_10786),
.Y(n_11628)
);

INVx2_ASAP7_75t_SL g11629 ( 
.A(n_11098),
.Y(n_11629)
);

AND2x2_ASAP7_75t_L g11630 ( 
.A(n_11136),
.B(n_10944),
.Y(n_11630)
);

INVx1_ASAP7_75t_L g11631 ( 
.A(n_11193),
.Y(n_11631)
);

NAND2xp5_ASAP7_75t_L g11632 ( 
.A(n_11055),
.B(n_10788),
.Y(n_11632)
);

INVx1_ASAP7_75t_L g11633 ( 
.A(n_11476),
.Y(n_11633)
);

NAND2xp5_ASAP7_75t_L g11634 ( 
.A(n_11298),
.B(n_11285),
.Y(n_11634)
);

INVx2_ASAP7_75t_SL g11635 ( 
.A(n_11112),
.Y(n_11635)
);

INVx1_ASAP7_75t_L g11636 ( 
.A(n_11493),
.Y(n_11636)
);

AND2x4_ASAP7_75t_L g11637 ( 
.A(n_11211),
.B(n_10846),
.Y(n_11637)
);

AND2x2_ASAP7_75t_L g11638 ( 
.A(n_11067),
.B(n_10954),
.Y(n_11638)
);

HB1xp67_ASAP7_75t_L g11639 ( 
.A(n_11080),
.Y(n_11639)
);

NAND2xp5_ASAP7_75t_L g11640 ( 
.A(n_11395),
.B(n_10788),
.Y(n_11640)
);

INVx2_ASAP7_75t_L g11641 ( 
.A(n_11061),
.Y(n_11641)
);

AND2x2_ASAP7_75t_L g11642 ( 
.A(n_11145),
.B(n_10570),
.Y(n_11642)
);

OR2x2_ASAP7_75t_L g11643 ( 
.A(n_11243),
.B(n_10885),
.Y(n_11643)
);

INVx1_ASAP7_75t_L g11644 ( 
.A(n_11275),
.Y(n_11644)
);

INVx2_ASAP7_75t_L g11645 ( 
.A(n_11061),
.Y(n_11645)
);

AND2x2_ASAP7_75t_L g11646 ( 
.A(n_11150),
.B(n_10980),
.Y(n_11646)
);

INVx2_ASAP7_75t_L g11647 ( 
.A(n_11056),
.Y(n_11647)
);

INVxp67_ASAP7_75t_SL g11648 ( 
.A(n_11203),
.Y(n_11648)
);

AND2x2_ASAP7_75t_L g11649 ( 
.A(n_11292),
.B(n_10854),
.Y(n_11649)
);

INVxp67_ASAP7_75t_L g11650 ( 
.A(n_11201),
.Y(n_11650)
);

INVx1_ASAP7_75t_L g11651 ( 
.A(n_11275),
.Y(n_11651)
);

INVx1_ASAP7_75t_L g11652 ( 
.A(n_11311),
.Y(n_11652)
);

BUFx3_ASAP7_75t_L g11653 ( 
.A(n_11312),
.Y(n_11653)
);

AND2x2_ASAP7_75t_L g11654 ( 
.A(n_11114),
.B(n_10855),
.Y(n_11654)
);

AND2x2_ASAP7_75t_L g11655 ( 
.A(n_11180),
.B(n_10864),
.Y(n_11655)
);

AND2x2_ASAP7_75t_L g11656 ( 
.A(n_11188),
.B(n_10865),
.Y(n_11656)
);

INVx2_ASAP7_75t_L g11657 ( 
.A(n_11056),
.Y(n_11657)
);

AND2x4_ASAP7_75t_L g11658 ( 
.A(n_11366),
.B(n_10869),
.Y(n_11658)
);

AND2x2_ASAP7_75t_L g11659 ( 
.A(n_11049),
.B(n_10874),
.Y(n_11659)
);

OR2x2_ASAP7_75t_L g11660 ( 
.A(n_11105),
.B(n_10794),
.Y(n_11660)
);

INVxp67_ASAP7_75t_SL g11661 ( 
.A(n_11079),
.Y(n_11661)
);

AND2x2_ASAP7_75t_L g11662 ( 
.A(n_11168),
.B(n_11086),
.Y(n_11662)
);

INVx2_ASAP7_75t_L g11663 ( 
.A(n_11056),
.Y(n_11663)
);

INVx1_ASAP7_75t_L g11664 ( 
.A(n_11311),
.Y(n_11664)
);

NAND2xp5_ASAP7_75t_L g11665 ( 
.A(n_11334),
.B(n_10792),
.Y(n_11665)
);

OR2x2_ASAP7_75t_L g11666 ( 
.A(n_11167),
.B(n_10800),
.Y(n_11666)
);

INVx2_ASAP7_75t_L g11667 ( 
.A(n_11157),
.Y(n_11667)
);

AND2x2_ASAP7_75t_L g11668 ( 
.A(n_11088),
.B(n_10878),
.Y(n_11668)
);

AND2x4_ASAP7_75t_SL g11669 ( 
.A(n_11250),
.B(n_10879),
.Y(n_11669)
);

OR2x2_ASAP7_75t_L g11670 ( 
.A(n_11176),
.B(n_10812),
.Y(n_11670)
);

NAND2xp5_ASAP7_75t_L g11671 ( 
.A(n_11042),
.B(n_10792),
.Y(n_11671)
);

AND2x2_ASAP7_75t_L g11672 ( 
.A(n_11250),
.B(n_10881),
.Y(n_11672)
);

INVx1_ASAP7_75t_L g11673 ( 
.A(n_11323),
.Y(n_11673)
);

NAND2xp5_ASAP7_75t_L g11674 ( 
.A(n_11043),
.B(n_10899),
.Y(n_11674)
);

INVx1_ASAP7_75t_L g11675 ( 
.A(n_11323),
.Y(n_11675)
);

NAND2xp5_ASAP7_75t_L g11676 ( 
.A(n_11046),
.B(n_10900),
.Y(n_11676)
);

AND2x2_ASAP7_75t_L g11677 ( 
.A(n_11261),
.B(n_10908),
.Y(n_11677)
);

INVx1_ASAP7_75t_L g11678 ( 
.A(n_11367),
.Y(n_11678)
);

AND2x2_ASAP7_75t_L g11679 ( 
.A(n_11261),
.B(n_10909),
.Y(n_11679)
);

AND2x4_ASAP7_75t_L g11680 ( 
.A(n_11212),
.B(n_10916),
.Y(n_11680)
);

NAND2x1_ASAP7_75t_L g11681 ( 
.A(n_11367),
.B(n_10526),
.Y(n_11681)
);

AND2x2_ASAP7_75t_L g11682 ( 
.A(n_11185),
.B(n_10922),
.Y(n_11682)
);

INVx1_ASAP7_75t_L g11683 ( 
.A(n_11178),
.Y(n_11683)
);

INVx1_ASAP7_75t_L g11684 ( 
.A(n_11182),
.Y(n_11684)
);

OR2x2_ASAP7_75t_L g11685 ( 
.A(n_11137),
.B(n_10871),
.Y(n_11685)
);

HB1xp67_ASAP7_75t_L g11686 ( 
.A(n_11209),
.Y(n_11686)
);

INVx1_ASAP7_75t_L g11687 ( 
.A(n_11082),
.Y(n_11687)
);

NAND2xp5_ASAP7_75t_L g11688 ( 
.A(n_11073),
.B(n_10927),
.Y(n_11688)
);

AND2x2_ASAP7_75t_L g11689 ( 
.A(n_11186),
.B(n_10933),
.Y(n_11689)
);

NAND2xp5_ASAP7_75t_L g11690 ( 
.A(n_11324),
.B(n_10938),
.Y(n_11690)
);

AND2x2_ASAP7_75t_L g11691 ( 
.A(n_11083),
.B(n_10950),
.Y(n_11691)
);

AND2x2_ASAP7_75t_L g11692 ( 
.A(n_11093),
.B(n_10952),
.Y(n_11692)
);

OR2x2_ASAP7_75t_L g11693 ( 
.A(n_11177),
.B(n_10791),
.Y(n_11693)
);

AND2x2_ASAP7_75t_L g11694 ( 
.A(n_11100),
.B(n_10956),
.Y(n_11694)
);

OR2x2_ASAP7_75t_L g11695 ( 
.A(n_11140),
.B(n_11004),
.Y(n_11695)
);

INVx1_ASAP7_75t_L g11696 ( 
.A(n_11407),
.Y(n_11696)
);

INVx1_ASAP7_75t_L g11697 ( 
.A(n_11428),
.Y(n_11697)
);

BUFx2_ASAP7_75t_L g11698 ( 
.A(n_11209),
.Y(n_11698)
);

AND2x4_ASAP7_75t_L g11699 ( 
.A(n_11216),
.B(n_11484),
.Y(n_11699)
);

INVx1_ASAP7_75t_L g11700 ( 
.A(n_11437),
.Y(n_11700)
);

HB1xp67_ASAP7_75t_L g11701 ( 
.A(n_11205),
.Y(n_11701)
);

INVx1_ASAP7_75t_L g11702 ( 
.A(n_11455),
.Y(n_11702)
);

INVx1_ASAP7_75t_L g11703 ( 
.A(n_11224),
.Y(n_11703)
);

NAND2xp5_ASAP7_75t_L g11704 ( 
.A(n_11438),
.B(n_10957),
.Y(n_11704)
);

AND2x4_ASAP7_75t_SL g11705 ( 
.A(n_11207),
.B(n_10959),
.Y(n_11705)
);

NAND2xp5_ASAP7_75t_L g11706 ( 
.A(n_11200),
.B(n_10963),
.Y(n_11706)
);

AND2x2_ASAP7_75t_L g11707 ( 
.A(n_11084),
.B(n_10965),
.Y(n_11707)
);

INVx2_ASAP7_75t_L g11708 ( 
.A(n_11157),
.Y(n_11708)
);

INVx1_ASAP7_75t_L g11709 ( 
.A(n_11338),
.Y(n_11709)
);

OR2x2_ASAP7_75t_L g11710 ( 
.A(n_11302),
.B(n_11013),
.Y(n_11710)
);

AND2x4_ASAP7_75t_L g11711 ( 
.A(n_11108),
.B(n_11027),
.Y(n_11711)
);

NOR2x1_ASAP7_75t_SL g11712 ( 
.A(n_11157),
.B(n_10526),
.Y(n_11712)
);

NOR2xp33_ASAP7_75t_L g11713 ( 
.A(n_11081),
.B(n_10943),
.Y(n_11713)
);

NAND2xp5_ASAP7_75t_SL g11714 ( 
.A(n_11274),
.B(n_10817),
.Y(n_11714)
);

INVx1_ASAP7_75t_L g11715 ( 
.A(n_11329),
.Y(n_11715)
);

AND2x2_ASAP7_75t_L g11716 ( 
.A(n_11281),
.B(n_10817),
.Y(n_11716)
);

AND2x2_ASAP7_75t_L g11717 ( 
.A(n_11099),
.B(n_11195),
.Y(n_11717)
);

INVx1_ASAP7_75t_L g11718 ( 
.A(n_11227),
.Y(n_11718)
);

NAND2xp5_ASAP7_75t_L g11719 ( 
.A(n_11388),
.B(n_10558),
.Y(n_11719)
);

OR2x2_ASAP7_75t_L g11720 ( 
.A(n_11313),
.B(n_10971),
.Y(n_11720)
);

INVx2_ASAP7_75t_L g11721 ( 
.A(n_11393),
.Y(n_11721)
);

AND2x2_ASAP7_75t_L g11722 ( 
.A(n_11120),
.B(n_10616),
.Y(n_11722)
);

INVx2_ASAP7_75t_SL g11723 ( 
.A(n_11358),
.Y(n_11723)
);

INVx1_ASAP7_75t_L g11724 ( 
.A(n_11230),
.Y(n_11724)
);

INVxp67_ASAP7_75t_L g11725 ( 
.A(n_11208),
.Y(n_11725)
);

INVx2_ASAP7_75t_L g11726 ( 
.A(n_11393),
.Y(n_11726)
);

INVx1_ASAP7_75t_L g11727 ( 
.A(n_11104),
.Y(n_11727)
);

NAND2xp5_ASAP7_75t_L g11728 ( 
.A(n_11416),
.B(n_10685),
.Y(n_11728)
);

INVx1_ASAP7_75t_L g11729 ( 
.A(n_11139),
.Y(n_11729)
);

NAND2xp5_ASAP7_75t_L g11730 ( 
.A(n_11441),
.B(n_10901),
.Y(n_11730)
);

NOR2xp33_ASAP7_75t_L g11731 ( 
.A(n_11390),
.B(n_10806),
.Y(n_11731)
);

INVx2_ASAP7_75t_L g11732 ( 
.A(n_11404),
.Y(n_11732)
);

INVx2_ASAP7_75t_L g11733 ( 
.A(n_11404),
.Y(n_11733)
);

NAND2xp5_ASAP7_75t_L g11734 ( 
.A(n_11142),
.B(n_10797),
.Y(n_11734)
);

INVx1_ASAP7_75t_L g11735 ( 
.A(n_11414),
.Y(n_11735)
);

OAI22xp5_ASAP7_75t_L g11736 ( 
.A1(n_11306),
.A2(n_10883),
.B1(n_9712),
.B2(n_9710),
.Y(n_11736)
);

HB1xp67_ASAP7_75t_SL g11737 ( 
.A(n_11272),
.Y(n_11737)
);

OR2x2_ASAP7_75t_L g11738 ( 
.A(n_11308),
.B(n_10616),
.Y(n_11738)
);

NAND2xp5_ASAP7_75t_L g11739 ( 
.A(n_11142),
.B(n_10336),
.Y(n_11739)
);

INVx1_ASAP7_75t_L g11740 ( 
.A(n_11414),
.Y(n_11740)
);

AND2x2_ASAP7_75t_L g11741 ( 
.A(n_11123),
.B(n_10719),
.Y(n_11741)
);

OAI21xp5_ASAP7_75t_SL g11742 ( 
.A1(n_11217),
.A2(n_10720),
.B(n_10719),
.Y(n_11742)
);

INVx1_ASAP7_75t_L g11743 ( 
.A(n_11440),
.Y(n_11743)
);

INVx3_ASAP7_75t_L g11744 ( 
.A(n_11090),
.Y(n_11744)
);

INVx1_ASAP7_75t_L g11745 ( 
.A(n_11032),
.Y(n_11745)
);

OR2x2_ASAP7_75t_L g11746 ( 
.A(n_11257),
.B(n_11373),
.Y(n_11746)
);

NAND2xp5_ASAP7_75t_L g11747 ( 
.A(n_11335),
.B(n_10720),
.Y(n_11747)
);

INVx1_ASAP7_75t_L g11748 ( 
.A(n_11249),
.Y(n_11748)
);

AND2x2_ASAP7_75t_L g11749 ( 
.A(n_11110),
.B(n_8475),
.Y(n_11749)
);

INVx1_ASAP7_75t_L g11750 ( 
.A(n_11249),
.Y(n_11750)
);

NAND2xp5_ASAP7_75t_L g11751 ( 
.A(n_11341),
.B(n_10970),
.Y(n_11751)
);

AND2x2_ASAP7_75t_L g11752 ( 
.A(n_11116),
.B(n_8516),
.Y(n_11752)
);

INVx2_ASAP7_75t_L g11753 ( 
.A(n_11408),
.Y(n_11753)
);

AND2x2_ASAP7_75t_L g11754 ( 
.A(n_11118),
.B(n_11365),
.Y(n_11754)
);

NAND2xp5_ASAP7_75t_L g11755 ( 
.A(n_11344),
.B(n_11011),
.Y(n_11755)
);

AND2x4_ASAP7_75t_L g11756 ( 
.A(n_11146),
.B(n_8516),
.Y(n_11756)
);

HB1xp67_ASAP7_75t_L g11757 ( 
.A(n_11450),
.Y(n_11757)
);

INVx1_ASAP7_75t_SL g11758 ( 
.A(n_11189),
.Y(n_11758)
);

INVx1_ASAP7_75t_L g11759 ( 
.A(n_11262),
.Y(n_11759)
);

OR2x2_ASAP7_75t_L g11760 ( 
.A(n_11263),
.B(n_11016),
.Y(n_11760)
);

OR2x2_ASAP7_75t_L g11761 ( 
.A(n_11379),
.B(n_8564),
.Y(n_11761)
);

INVx1_ASAP7_75t_L g11762 ( 
.A(n_11262),
.Y(n_11762)
);

INVx2_ASAP7_75t_L g11763 ( 
.A(n_11408),
.Y(n_11763)
);

AND2x2_ASAP7_75t_L g11764 ( 
.A(n_11467),
.B(n_8516),
.Y(n_11764)
);

AND2x2_ASAP7_75t_L g11765 ( 
.A(n_11269),
.B(n_11096),
.Y(n_11765)
);

AND2x2_ASAP7_75t_L g11766 ( 
.A(n_11361),
.B(n_8524),
.Y(n_11766)
);

INVx1_ASAP7_75t_L g11767 ( 
.A(n_11305),
.Y(n_11767)
);

INVx1_ASAP7_75t_L g11768 ( 
.A(n_11305),
.Y(n_11768)
);

AND2x4_ASAP7_75t_L g11769 ( 
.A(n_11153),
.B(n_8524),
.Y(n_11769)
);

AND2x2_ASAP7_75t_L g11770 ( 
.A(n_11369),
.B(n_8524),
.Y(n_11770)
);

AND2x2_ASAP7_75t_L g11771 ( 
.A(n_11384),
.B(n_8557),
.Y(n_11771)
);

INVx1_ASAP7_75t_L g11772 ( 
.A(n_11398),
.Y(n_11772)
);

INVx1_ASAP7_75t_L g11773 ( 
.A(n_11480),
.Y(n_11773)
);

NAND2xp5_ASAP7_75t_L g11774 ( 
.A(n_11353),
.B(n_10966),
.Y(n_11774)
);

INVx1_ASAP7_75t_L g11775 ( 
.A(n_11486),
.Y(n_11775)
);

OR2x2_ASAP7_75t_L g11776 ( 
.A(n_11317),
.B(n_8565),
.Y(n_11776)
);

INVx1_ASAP7_75t_L g11777 ( 
.A(n_11044),
.Y(n_11777)
);

INVx1_ASAP7_75t_L g11778 ( 
.A(n_11052),
.Y(n_11778)
);

OR2x2_ASAP7_75t_L g11779 ( 
.A(n_11359),
.B(n_8565),
.Y(n_11779)
);

INVx2_ASAP7_75t_SL g11780 ( 
.A(n_11358),
.Y(n_11780)
);

INVx2_ASAP7_75t_L g11781 ( 
.A(n_11413),
.Y(n_11781)
);

BUFx2_ASAP7_75t_L g11782 ( 
.A(n_11170),
.Y(n_11782)
);

HB1xp67_ASAP7_75t_L g11783 ( 
.A(n_11194),
.Y(n_11783)
);

NAND2xp5_ASAP7_75t_L g11784 ( 
.A(n_11351),
.B(n_8568),
.Y(n_11784)
);

INVx1_ASAP7_75t_L g11785 ( 
.A(n_11036),
.Y(n_11785)
);

AND2x4_ASAP7_75t_L g11786 ( 
.A(n_11090),
.B(n_8557),
.Y(n_11786)
);

INVx3_ASAP7_75t_L g11787 ( 
.A(n_11235),
.Y(n_11787)
);

INVx1_ASAP7_75t_L g11788 ( 
.A(n_11037),
.Y(n_11788)
);

HB1xp67_ASAP7_75t_L g11789 ( 
.A(n_11413),
.Y(n_11789)
);

NAND2x1p5_ASAP7_75t_L g11790 ( 
.A(n_11390),
.B(n_6245),
.Y(n_11790)
);

INVx1_ASAP7_75t_L g11791 ( 
.A(n_11030),
.Y(n_11791)
);

AND2x2_ASAP7_75t_L g11792 ( 
.A(n_11392),
.B(n_8557),
.Y(n_11792)
);

INVx1_ASAP7_75t_L g11793 ( 
.A(n_11039),
.Y(n_11793)
);

AND2x2_ASAP7_75t_L g11794 ( 
.A(n_11396),
.B(n_8561),
.Y(n_11794)
);

INVx1_ASAP7_75t_L g11795 ( 
.A(n_11041),
.Y(n_11795)
);

INVx2_ASAP7_75t_L g11796 ( 
.A(n_11070),
.Y(n_11796)
);

AND2x4_ASAP7_75t_L g11797 ( 
.A(n_11235),
.B(n_8561),
.Y(n_11797)
);

AND2x2_ASAP7_75t_L g11798 ( 
.A(n_11469),
.B(n_8561),
.Y(n_11798)
);

AND2x2_ASAP7_75t_L g11799 ( 
.A(n_11470),
.B(n_8574),
.Y(n_11799)
);

OR2x2_ASAP7_75t_L g11800 ( 
.A(n_11316),
.B(n_8568),
.Y(n_11800)
);

INVx1_ASAP7_75t_L g11801 ( 
.A(n_11435),
.Y(n_11801)
);

AND2x2_ASAP7_75t_L g11802 ( 
.A(n_11252),
.B(n_8574),
.Y(n_11802)
);

INVx1_ASAP7_75t_L g11803 ( 
.A(n_11060),
.Y(n_11803)
);

NAND2xp5_ASAP7_75t_L g11804 ( 
.A(n_11265),
.B(n_8576),
.Y(n_11804)
);

NAND2xp5_ASAP7_75t_L g11805 ( 
.A(n_11265),
.B(n_8576),
.Y(n_11805)
);

OR2x2_ASAP7_75t_L g11806 ( 
.A(n_11340),
.B(n_8577),
.Y(n_11806)
);

BUFx3_ASAP7_75t_L g11807 ( 
.A(n_11172),
.Y(n_11807)
);

NAND2xp5_ASAP7_75t_L g11808 ( 
.A(n_11282),
.B(n_11284),
.Y(n_11808)
);

INVxp67_ASAP7_75t_SL g11809 ( 
.A(n_11057),
.Y(n_11809)
);

NAND2xp5_ASAP7_75t_L g11810 ( 
.A(n_11282),
.B(n_8577),
.Y(n_11810)
);

AND2x2_ASAP7_75t_L g11811 ( 
.A(n_11307),
.B(n_11487),
.Y(n_11811)
);

INVx1_ASAP7_75t_L g11812 ( 
.A(n_11442),
.Y(n_11812)
);

BUFx2_ASAP7_75t_L g11813 ( 
.A(n_11070),
.Y(n_11813)
);

INVx4_ASAP7_75t_L g11814 ( 
.A(n_11358),
.Y(n_11814)
);

AND2x2_ASAP7_75t_L g11815 ( 
.A(n_11487),
.B(n_8574),
.Y(n_11815)
);

INVx2_ASAP7_75t_L g11816 ( 
.A(n_11497),
.Y(n_11816)
);

AND2x2_ASAP7_75t_L g11817 ( 
.A(n_11436),
.B(n_8580),
.Y(n_11817)
);

OR2x2_ASAP7_75t_L g11818 ( 
.A(n_11477),
.B(n_11397),
.Y(n_11818)
);

NAND2xp5_ASAP7_75t_L g11819 ( 
.A(n_11284),
.B(n_11288),
.Y(n_11819)
);

INVx2_ASAP7_75t_L g11820 ( 
.A(n_11497),
.Y(n_11820)
);

INVx1_ASAP7_75t_L g11821 ( 
.A(n_11175),
.Y(n_11821)
);

INVx1_ASAP7_75t_L g11822 ( 
.A(n_11264),
.Y(n_11822)
);

NOR2xp33_ASAP7_75t_L g11823 ( 
.A(n_11270),
.B(n_8097),
.Y(n_11823)
);

INVx1_ASAP7_75t_L g11824 ( 
.A(n_11267),
.Y(n_11824)
);

INVx1_ASAP7_75t_L g11825 ( 
.A(n_11271),
.Y(n_11825)
);

AND2x2_ASAP7_75t_L g11826 ( 
.A(n_11417),
.B(n_8580),
.Y(n_11826)
);

AND2x2_ASAP7_75t_SL g11827 ( 
.A(n_11380),
.B(n_10262),
.Y(n_11827)
);

AND2x2_ASAP7_75t_L g11828 ( 
.A(n_11421),
.B(n_8580),
.Y(n_11828)
);

AND2x2_ASAP7_75t_L g11829 ( 
.A(n_11463),
.B(n_8420),
.Y(n_11829)
);

NAND2xp5_ASAP7_75t_L g11830 ( 
.A(n_11288),
.B(n_8578),
.Y(n_11830)
);

AND2x2_ASAP7_75t_L g11831 ( 
.A(n_11478),
.B(n_8421),
.Y(n_11831)
);

HB1xp67_ASAP7_75t_L g11832 ( 
.A(n_11422),
.Y(n_11832)
);

HB1xp67_ASAP7_75t_L g11833 ( 
.A(n_11424),
.Y(n_11833)
);

NAND2xp5_ASAP7_75t_L g11834 ( 
.A(n_11381),
.B(n_11382),
.Y(n_11834)
);

INVx1_ASAP7_75t_L g11835 ( 
.A(n_11273),
.Y(n_11835)
);

INVx1_ASAP7_75t_L g11836 ( 
.A(n_11278),
.Y(n_11836)
);

NAND2xp5_ASAP7_75t_L g11837 ( 
.A(n_11383),
.B(n_8578),
.Y(n_11837)
);

INVx2_ASAP7_75t_L g11838 ( 
.A(n_11300),
.Y(n_11838)
);

AND2x2_ASAP7_75t_L g11839 ( 
.A(n_11051),
.B(n_8579),
.Y(n_11839)
);

INVx1_ASAP7_75t_L g11840 ( 
.A(n_11280),
.Y(n_11840)
);

NAND2xp5_ASAP7_75t_L g11841 ( 
.A(n_11391),
.B(n_11394),
.Y(n_11841)
);

OR2x2_ASAP7_75t_L g11842 ( 
.A(n_11279),
.B(n_8579),
.Y(n_11842)
);

INVx1_ASAP7_75t_L g11843 ( 
.A(n_11286),
.Y(n_11843)
);

AND2x2_ASAP7_75t_L g11844 ( 
.A(n_11240),
.B(n_8589),
.Y(n_11844)
);

INVx2_ASAP7_75t_L g11845 ( 
.A(n_11303),
.Y(n_11845)
);

OR2x2_ASAP7_75t_L g11846 ( 
.A(n_11479),
.B(n_8589),
.Y(n_11846)
);

AND2x4_ASAP7_75t_SL g11847 ( 
.A(n_11240),
.B(n_6847),
.Y(n_11847)
);

AND2x4_ASAP7_75t_L g11848 ( 
.A(n_11126),
.B(n_11128),
.Y(n_11848)
);

OR2x2_ASAP7_75t_L g11849 ( 
.A(n_11054),
.B(n_8590),
.Y(n_11849)
);

INVx2_ASAP7_75t_SL g11850 ( 
.A(n_11289),
.Y(n_11850)
);

NAND2xp5_ASAP7_75t_L g11851 ( 
.A(n_11289),
.B(n_11451),
.Y(n_11851)
);

AND2x2_ASAP7_75t_L g11852 ( 
.A(n_11343),
.B(n_8590),
.Y(n_11852)
);

INVx2_ASAP7_75t_L g11853 ( 
.A(n_11244),
.Y(n_11853)
);

AND2x4_ASAP7_75t_L g11854 ( 
.A(n_11158),
.B(n_8594),
.Y(n_11854)
);

OAI21xp5_ASAP7_75t_L g11855 ( 
.A1(n_11206),
.A2(n_9106),
.B(n_8874),
.Y(n_11855)
);

INVx1_ASAP7_75t_L g11856 ( 
.A(n_11290),
.Y(n_11856)
);

BUFx2_ASAP7_75t_L g11857 ( 
.A(n_11403),
.Y(n_11857)
);

NAND2xp5_ASAP7_75t_SL g11858 ( 
.A(n_11181),
.B(n_8097),
.Y(n_11858)
);

NAND2x1p5_ASAP7_75t_L g11859 ( 
.A(n_11255),
.B(n_11166),
.Y(n_11859)
);

OR2x2_ASAP7_75t_L g11860 ( 
.A(n_11058),
.B(n_8594),
.Y(n_11860)
);

INVx1_ASAP7_75t_L g11861 ( 
.A(n_11346),
.Y(n_11861)
);

AND2x2_ASAP7_75t_L g11862 ( 
.A(n_11174),
.B(n_8607),
.Y(n_11862)
);

NAND2xp5_ASAP7_75t_L g11863 ( 
.A(n_11401),
.B(n_8607),
.Y(n_11863)
);

AND2x2_ASAP7_75t_L g11864 ( 
.A(n_11113),
.B(n_11501),
.Y(n_11864)
);

INVx2_ASAP7_75t_SL g11865 ( 
.A(n_11220),
.Y(n_11865)
);

AND2x4_ASAP7_75t_L g11866 ( 
.A(n_11228),
.B(n_8609),
.Y(n_11866)
);

HB1xp67_ASAP7_75t_L g11867 ( 
.A(n_11425),
.Y(n_11867)
);

NOR2xp67_ASAP7_75t_L g11868 ( 
.A(n_11244),
.B(n_8894),
.Y(n_11868)
);

AND2x2_ASAP7_75t_L g11869 ( 
.A(n_11095),
.B(n_8609),
.Y(n_11869)
);

AND2x2_ASAP7_75t_L g11870 ( 
.A(n_11228),
.B(n_8634),
.Y(n_11870)
);

INVx2_ASAP7_75t_L g11871 ( 
.A(n_11258),
.Y(n_11871)
);

INVx1_ASAP7_75t_L g11872 ( 
.A(n_11349),
.Y(n_11872)
);

NAND2xp5_ASAP7_75t_L g11873 ( 
.A(n_11449),
.B(n_8634),
.Y(n_11873)
);

INVxp67_ASAP7_75t_L g11874 ( 
.A(n_11328),
.Y(n_11874)
);

NOR2x1_ASAP7_75t_L g11875 ( 
.A(n_11214),
.B(n_10271),
.Y(n_11875)
);

NOR2xp67_ASAP7_75t_L g11876 ( 
.A(n_11258),
.B(n_8894),
.Y(n_11876)
);

INVx1_ASAP7_75t_L g11877 ( 
.A(n_11350),
.Y(n_11877)
);

AND2x4_ASAP7_75t_L g11878 ( 
.A(n_11173),
.B(n_8894),
.Y(n_11878)
);

INVx1_ASAP7_75t_L g11879 ( 
.A(n_11354),
.Y(n_11879)
);

AND2x2_ASAP7_75t_L g11880 ( 
.A(n_11474),
.B(n_7334),
.Y(n_11880)
);

AND2x4_ASAP7_75t_L g11881 ( 
.A(n_11173),
.B(n_8901),
.Y(n_11881)
);

AND2x2_ASAP7_75t_L g11882 ( 
.A(n_11197),
.B(n_7334),
.Y(n_11882)
);

INVx3_ASAP7_75t_L g11883 ( 
.A(n_11198),
.Y(n_11883)
);

AND2x2_ASAP7_75t_L g11884 ( 
.A(n_11283),
.B(n_7334),
.Y(n_11884)
);

INVx1_ASAP7_75t_L g11885 ( 
.A(n_11360),
.Y(n_11885)
);

AND2x2_ASAP7_75t_L g11886 ( 
.A(n_11198),
.B(n_7392),
.Y(n_11886)
);

INVx1_ASAP7_75t_L g11887 ( 
.A(n_11364),
.Y(n_11887)
);

BUFx2_ASAP7_75t_L g11888 ( 
.A(n_11415),
.Y(n_11888)
);

OR2x2_ASAP7_75t_L g11889 ( 
.A(n_11423),
.B(n_8422),
.Y(n_11889)
);

AND2x2_ASAP7_75t_L g11890 ( 
.A(n_11210),
.B(n_7392),
.Y(n_11890)
);

AND2x2_ASAP7_75t_L g11891 ( 
.A(n_11210),
.B(n_11378),
.Y(n_11891)
);

INVx1_ASAP7_75t_L g11892 ( 
.A(n_11368),
.Y(n_11892)
);

INVx1_ASAP7_75t_L g11893 ( 
.A(n_11370),
.Y(n_11893)
);

AND2x2_ASAP7_75t_L g11894 ( 
.A(n_11434),
.B(n_7392),
.Y(n_11894)
);

OR2x2_ASAP7_75t_L g11895 ( 
.A(n_11427),
.B(n_8422),
.Y(n_11895)
);

INVx1_ASAP7_75t_L g11896 ( 
.A(n_11352),
.Y(n_11896)
);

INVx1_ASAP7_75t_L g11897 ( 
.A(n_11355),
.Y(n_11897)
);

AND2x2_ASAP7_75t_L g11898 ( 
.A(n_11426),
.B(n_8423),
.Y(n_11898)
);

AND2x2_ASAP7_75t_L g11899 ( 
.A(n_11502),
.B(n_8423),
.Y(n_11899)
);

INVx1_ASAP7_75t_L g11900 ( 
.A(n_11443),
.Y(n_11900)
);

INVx2_ASAP7_75t_L g11901 ( 
.A(n_11443),
.Y(n_11901)
);

AND2x2_ASAP7_75t_SL g11902 ( 
.A(n_11457),
.B(n_10989),
.Y(n_11902)
);

INVx2_ASAP7_75t_L g11903 ( 
.A(n_11465),
.Y(n_11903)
);

AND2x2_ASAP7_75t_L g11904 ( 
.A(n_11504),
.B(n_8425),
.Y(n_11904)
);

AND2x2_ASAP7_75t_L g11905 ( 
.A(n_11500),
.B(n_8425),
.Y(n_11905)
);

INVx1_ASAP7_75t_L g11906 ( 
.A(n_11345),
.Y(n_11906)
);

AND2x2_ASAP7_75t_L g11907 ( 
.A(n_11363),
.B(n_8444),
.Y(n_11907)
);

AND2x2_ASAP7_75t_L g11908 ( 
.A(n_11371),
.B(n_8444),
.Y(n_11908)
);

INVx1_ASAP7_75t_L g11909 ( 
.A(n_11064),
.Y(n_11909)
);

INVx2_ASAP7_75t_SL g11910 ( 
.A(n_11432),
.Y(n_11910)
);

NAND3xp33_ASAP7_75t_L g11911 ( 
.A(n_11122),
.B(n_10993),
.C(n_10167),
.Y(n_11911)
);

NAND2xp5_ASAP7_75t_L g11912 ( 
.A(n_11483),
.B(n_6852),
.Y(n_11912)
);

OR2x2_ASAP7_75t_L g11913 ( 
.A(n_11418),
.B(n_11400),
.Y(n_11913)
);

INVx1_ASAP7_75t_L g11914 ( 
.A(n_11066),
.Y(n_11914)
);

OR2x2_ASAP7_75t_L g11915 ( 
.A(n_11491),
.B(n_8458),
.Y(n_11915)
);

HB1xp67_ASAP7_75t_L g11916 ( 
.A(n_11245),
.Y(n_11916)
);

AND2x2_ASAP7_75t_L g11917 ( 
.A(n_11374),
.B(n_8458),
.Y(n_11917)
);

NAND2xp5_ASAP7_75t_L g11918 ( 
.A(n_11456),
.B(n_6852),
.Y(n_11918)
);

INVx2_ASAP7_75t_L g11919 ( 
.A(n_11468),
.Y(n_11919)
);

AND2x2_ASAP7_75t_L g11920 ( 
.A(n_11246),
.B(n_8459),
.Y(n_11920)
);

AND2x2_ASAP7_75t_L g11921 ( 
.A(n_11488),
.B(n_8459),
.Y(n_11921)
);

INVx3_ASAP7_75t_L g11922 ( 
.A(n_11331),
.Y(n_11922)
);

AND2x2_ASAP7_75t_L g11923 ( 
.A(n_11489),
.B(n_8468),
.Y(n_11923)
);

NAND2xp5_ASAP7_75t_L g11924 ( 
.A(n_11462),
.B(n_6852),
.Y(n_11924)
);

INVx1_ASAP7_75t_L g11925 ( 
.A(n_11071),
.Y(n_11925)
);

INVx1_ASAP7_75t_L g11926 ( 
.A(n_11085),
.Y(n_11926)
);

AND2x2_ASAP7_75t_L g11927 ( 
.A(n_11464),
.B(n_8468),
.Y(n_11927)
);

AND2x2_ASAP7_75t_L g11928 ( 
.A(n_11475),
.B(n_8490),
.Y(n_11928)
);

INVx1_ASAP7_75t_L g11929 ( 
.A(n_11453),
.Y(n_11929)
);

INVx2_ASAP7_75t_L g11930 ( 
.A(n_11490),
.Y(n_11930)
);

INVx2_ASAP7_75t_L g11931 ( 
.A(n_11490),
.Y(n_11931)
);

NAND2xp5_ASAP7_75t_L g11932 ( 
.A(n_11466),
.B(n_6852),
.Y(n_11932)
);

AND2x2_ASAP7_75t_L g11933 ( 
.A(n_11331),
.B(n_11348),
.Y(n_11933)
);

INVx1_ASAP7_75t_L g11934 ( 
.A(n_11454),
.Y(n_11934)
);

INVx1_ASAP7_75t_L g11935 ( 
.A(n_11183),
.Y(n_11935)
);

INVx2_ASAP7_75t_L g11936 ( 
.A(n_11494),
.Y(n_11936)
);

INVx1_ASAP7_75t_L g11937 ( 
.A(n_11184),
.Y(n_11937)
);

NAND2xp5_ASAP7_75t_L g11938 ( 
.A(n_11362),
.B(n_7225),
.Y(n_11938)
);

AND2x2_ASAP7_75t_L g11939 ( 
.A(n_11348),
.B(n_8490),
.Y(n_11939)
);

AND2x2_ASAP7_75t_L g11940 ( 
.A(n_11223),
.B(n_8494),
.Y(n_11940)
);

NAND2xp5_ASAP7_75t_L g11941 ( 
.A(n_11202),
.B(n_11459),
.Y(n_11941)
);

OR2x2_ASAP7_75t_L g11942 ( 
.A(n_11481),
.B(n_8494),
.Y(n_11942)
);

AND2x2_ASAP7_75t_L g11943 ( 
.A(n_11242),
.B(n_8499),
.Y(n_11943)
);

NOR2xp67_ASAP7_75t_L g11944 ( 
.A(n_11495),
.B(n_8901),
.Y(n_11944)
);

AND2x2_ASAP7_75t_L g11945 ( 
.A(n_11540),
.B(n_11333),
.Y(n_11945)
);

INVx1_ASAP7_75t_L g11946 ( 
.A(n_11583),
.Y(n_11946)
);

AND2x4_ASAP7_75t_L g11947 ( 
.A(n_11549),
.B(n_11498),
.Y(n_11947)
);

AND2x2_ASAP7_75t_L g11948 ( 
.A(n_11544),
.B(n_11372),
.Y(n_11948)
);

AND2x4_ASAP7_75t_L g11949 ( 
.A(n_11653),
.B(n_11092),
.Y(n_11949)
);

INVx1_ASAP7_75t_L g11950 ( 
.A(n_11583),
.Y(n_11950)
);

NOR2xp33_ASAP7_75t_L g11951 ( 
.A(n_11737),
.B(n_11179),
.Y(n_11951)
);

AND2x2_ASAP7_75t_L g11952 ( 
.A(n_11520),
.B(n_11094),
.Y(n_11952)
);

AND2x4_ASAP7_75t_L g11953 ( 
.A(n_11850),
.B(n_11107),
.Y(n_11953)
);

NAND2xp5_ASAP7_75t_L g11954 ( 
.A(n_11593),
.B(n_11551),
.Y(n_11954)
);

AND2x2_ASAP7_75t_L g11955 ( 
.A(n_11783),
.B(n_11115),
.Y(n_11955)
);

AND2x2_ASAP7_75t_L g11956 ( 
.A(n_11717),
.B(n_11135),
.Y(n_11956)
);

INVx2_ASAP7_75t_L g11957 ( 
.A(n_11527),
.Y(n_11957)
);

OAI33xp33_ASAP7_75t_L g11958 ( 
.A1(n_11521),
.A2(n_11256),
.A3(n_11236),
.B1(n_11330),
.B2(n_11247),
.B3(n_11234),
.Y(n_11958)
);

INVx2_ASAP7_75t_L g11959 ( 
.A(n_11527),
.Y(n_11959)
);

NAND2xp5_ASAP7_75t_L g11960 ( 
.A(n_11758),
.B(n_11143),
.Y(n_11960)
);

AND2x2_ASAP7_75t_L g11961 ( 
.A(n_11509),
.B(n_11147),
.Y(n_11961)
);

INVx1_ASAP7_75t_L g11962 ( 
.A(n_11757),
.Y(n_11962)
);

INVx1_ASAP7_75t_L g11963 ( 
.A(n_11570),
.Y(n_11963)
);

NAND2xp5_ASAP7_75t_L g11964 ( 
.A(n_11615),
.B(n_11149),
.Y(n_11964)
);

OR2x2_ASAP7_75t_L g11965 ( 
.A(n_11582),
.B(n_11151),
.Y(n_11965)
);

BUFx3_ASAP7_75t_L g11966 ( 
.A(n_11699),
.Y(n_11966)
);

OR2x2_ASAP7_75t_L g11967 ( 
.A(n_11569),
.B(n_11154),
.Y(n_11967)
);

AND2x2_ASAP7_75t_L g11968 ( 
.A(n_11595),
.B(n_11765),
.Y(n_11968)
);

AND2x2_ASAP7_75t_L g11969 ( 
.A(n_11577),
.B(n_11155),
.Y(n_11969)
);

AND2x2_ASAP7_75t_L g11970 ( 
.A(n_11562),
.B(n_11530),
.Y(n_11970)
);

AND2x2_ASAP7_75t_L g11971 ( 
.A(n_11662),
.B(n_11604),
.Y(n_11971)
);

INVx1_ASAP7_75t_L g11972 ( 
.A(n_11570),
.Y(n_11972)
);

INVx1_ASAP7_75t_L g11973 ( 
.A(n_11698),
.Y(n_11973)
);

AND2x2_ASAP7_75t_L g11974 ( 
.A(n_11539),
.B(n_11162),
.Y(n_11974)
);

INVx1_ASAP7_75t_SL g11975 ( 
.A(n_11515),
.Y(n_11975)
);

HB1xp67_ASAP7_75t_L g11976 ( 
.A(n_11515),
.Y(n_11976)
);

INVx1_ASAP7_75t_L g11977 ( 
.A(n_11698),
.Y(n_11977)
);

NAND2xp5_ASAP7_75t_L g11978 ( 
.A(n_11699),
.B(n_11461),
.Y(n_11978)
);

AND2x4_ASAP7_75t_L g11979 ( 
.A(n_11508),
.B(n_11332),
.Y(n_11979)
);

NAND2xp5_ASAP7_75t_L g11980 ( 
.A(n_11635),
.B(n_11472),
.Y(n_11980)
);

INVx1_ASAP7_75t_L g11981 ( 
.A(n_11613),
.Y(n_11981)
);

NOR2xp33_ASAP7_75t_L g11982 ( 
.A(n_11814),
.B(n_11089),
.Y(n_11982)
);

INVx1_ASAP7_75t_L g11983 ( 
.A(n_11613),
.Y(n_11983)
);

INVx1_ASAP7_75t_L g11984 ( 
.A(n_11686),
.Y(n_11984)
);

AND2x2_ASAP7_75t_L g11985 ( 
.A(n_11518),
.B(n_11563),
.Y(n_11985)
);

INVx1_ASAP7_75t_L g11986 ( 
.A(n_11639),
.Y(n_11986)
);

AND2x2_ASAP7_75t_L g11987 ( 
.A(n_11522),
.B(n_11499),
.Y(n_11987)
);

INVx1_ASAP7_75t_L g11988 ( 
.A(n_11681),
.Y(n_11988)
);

NAND2xp5_ASAP7_75t_L g11989 ( 
.A(n_11744),
.B(n_11496),
.Y(n_11989)
);

INVx1_ASAP7_75t_L g11990 ( 
.A(n_11681),
.Y(n_11990)
);

BUFx3_ASAP7_75t_L g11991 ( 
.A(n_11859),
.Y(n_11991)
);

INVx2_ASAP7_75t_L g11992 ( 
.A(n_11814),
.Y(n_11992)
);

INVx1_ASAP7_75t_L g11993 ( 
.A(n_11772),
.Y(n_11993)
);

INVx1_ASAP7_75t_L g11994 ( 
.A(n_11514),
.Y(n_11994)
);

AND2x2_ASAP7_75t_L g11995 ( 
.A(n_11505),
.B(n_11458),
.Y(n_11995)
);

AND2x2_ASAP7_75t_L g11996 ( 
.A(n_11621),
.B(n_11460),
.Y(n_11996)
);

INVx1_ASAP7_75t_L g11997 ( 
.A(n_11743),
.Y(n_11997)
);

NAND2xp5_ASAP7_75t_L g11998 ( 
.A(n_11787),
.B(n_11430),
.Y(n_11998)
);

AND2x2_ASAP7_75t_L g11999 ( 
.A(n_11599),
.B(n_11429),
.Y(n_11999)
);

AOI22xp33_ASAP7_75t_L g12000 ( 
.A1(n_11605),
.A2(n_11412),
.B1(n_11229),
.B2(n_11132),
.Y(n_12000)
);

NAND2xp5_ASAP7_75t_L g12001 ( 
.A(n_11668),
.B(n_11433),
.Y(n_12001)
);

AND2x4_ASAP7_75t_SL g12002 ( 
.A(n_11510),
.B(n_11494),
.Y(n_12002)
);

HB1xp67_ASAP7_75t_L g12003 ( 
.A(n_11623),
.Y(n_12003)
);

INVx2_ASAP7_75t_L g12004 ( 
.A(n_11510),
.Y(n_12004)
);

INVx1_ASAP7_75t_L g12005 ( 
.A(n_11789),
.Y(n_12005)
);

AND2x2_ASAP7_75t_L g12006 ( 
.A(n_11610),
.B(n_11503),
.Y(n_12006)
);

AND2x2_ASAP7_75t_L g12007 ( 
.A(n_11638),
.B(n_11608),
.Y(n_12007)
);

INVx1_ASAP7_75t_L g12008 ( 
.A(n_11513),
.Y(n_12008)
);

AND2x2_ASAP7_75t_L g12009 ( 
.A(n_11682),
.B(n_11503),
.Y(n_12009)
);

AND2x2_ASAP7_75t_L g12010 ( 
.A(n_11689),
.B(n_11291),
.Y(n_12010)
);

AND2x2_ASAP7_75t_L g12011 ( 
.A(n_11606),
.B(n_11320),
.Y(n_12011)
);

INVx2_ASAP7_75t_L g12012 ( 
.A(n_11534),
.Y(n_12012)
);

OR2x2_ASAP7_75t_L g12013 ( 
.A(n_11597),
.B(n_11321),
.Y(n_12013)
);

INVx1_ASAP7_75t_L g12014 ( 
.A(n_11516),
.Y(n_12014)
);

INVx1_ASAP7_75t_L g12015 ( 
.A(n_11916),
.Y(n_12015)
);

INVx1_ASAP7_75t_SL g12016 ( 
.A(n_11782),
.Y(n_12016)
);

INVx1_ASAP7_75t_L g12017 ( 
.A(n_11607),
.Y(n_12017)
);

INVx2_ASAP7_75t_L g12018 ( 
.A(n_11723),
.Y(n_12018)
);

NAND3xp33_ASAP7_75t_L g12019 ( 
.A(n_11742),
.B(n_11078),
.C(n_11190),
.Y(n_12019)
);

AND2x2_ASAP7_75t_L g12020 ( 
.A(n_11598),
.B(n_11325),
.Y(n_12020)
);

NAND2xp5_ASAP7_75t_L g12021 ( 
.A(n_11713),
.B(n_11192),
.Y(n_12021)
);

INVx2_ASAP7_75t_SL g12022 ( 
.A(n_11584),
.Y(n_12022)
);

AND2x2_ASAP7_75t_L g12023 ( 
.A(n_11630),
.B(n_11326),
.Y(n_12023)
);

INVx1_ASAP7_75t_L g12024 ( 
.A(n_11600),
.Y(n_12024)
);

INVx2_ASAP7_75t_SL g12025 ( 
.A(n_11933),
.Y(n_12025)
);

NAND2xp5_ASAP7_75t_L g12026 ( 
.A(n_11694),
.B(n_11213),
.Y(n_12026)
);

NAND2xp5_ASAP7_75t_L g12027 ( 
.A(n_11654),
.B(n_11446),
.Y(n_12027)
);

AND2x2_ASAP7_75t_L g12028 ( 
.A(n_11609),
.B(n_11447),
.Y(n_12028)
);

AND2x2_ASAP7_75t_L g12029 ( 
.A(n_11626),
.B(n_11448),
.Y(n_12029)
);

INVx3_ASAP7_75t_L g12030 ( 
.A(n_11560),
.Y(n_12030)
);

AND2x2_ASAP7_75t_L g12031 ( 
.A(n_11646),
.B(n_11452),
.Y(n_12031)
);

AND2x2_ASAP7_75t_L g12032 ( 
.A(n_11506),
.B(n_11337),
.Y(n_12032)
);

AND2x2_ASAP7_75t_L g12033 ( 
.A(n_11655),
.B(n_11342),
.Y(n_12033)
);

NOR2xp33_ASAP7_75t_L g12034 ( 
.A(n_11553),
.B(n_11492),
.Y(n_12034)
);

AND2x4_ASAP7_75t_L g12035 ( 
.A(n_11560),
.B(n_11219),
.Y(n_12035)
);

INVx1_ASAP7_75t_L g12036 ( 
.A(n_11729),
.Y(n_12036)
);

INVx1_ASAP7_75t_SL g12037 ( 
.A(n_11782),
.Y(n_12037)
);

INVx1_ASAP7_75t_L g12038 ( 
.A(n_11661),
.Y(n_12038)
);

INVx1_ASAP7_75t_L g12039 ( 
.A(n_11691),
.Y(n_12039)
);

AND2x2_ASAP7_75t_L g12040 ( 
.A(n_11754),
.B(n_11471),
.Y(n_12040)
);

INVx1_ASAP7_75t_L g12041 ( 
.A(n_11692),
.Y(n_12041)
);

INVx1_ASAP7_75t_L g12042 ( 
.A(n_11644),
.Y(n_12042)
);

AND2x2_ASAP7_75t_L g12043 ( 
.A(n_11642),
.B(n_11233),
.Y(n_12043)
);

INVx2_ASAP7_75t_L g12044 ( 
.A(n_11780),
.Y(n_12044)
);

NAND2xp5_ASAP7_75t_L g12045 ( 
.A(n_11707),
.B(n_11293),
.Y(n_12045)
);

NOR2xp33_ASAP7_75t_R g12046 ( 
.A(n_11619),
.B(n_8097),
.Y(n_12046)
);

AND2x2_ASAP7_75t_L g12047 ( 
.A(n_11622),
.B(n_11439),
.Y(n_12047)
);

INVx1_ASAP7_75t_L g12048 ( 
.A(n_11651),
.Y(n_12048)
);

INVx1_ASAP7_75t_L g12049 ( 
.A(n_11652),
.Y(n_12049)
);

INVx1_ASAP7_75t_L g12050 ( 
.A(n_11664),
.Y(n_12050)
);

INVx1_ASAP7_75t_L g12051 ( 
.A(n_11673),
.Y(n_12051)
);

INVx1_ASAP7_75t_L g12052 ( 
.A(n_11675),
.Y(n_12052)
);

OR2x2_ASAP7_75t_L g12053 ( 
.A(n_11632),
.B(n_11187),
.Y(n_12053)
);

INVx1_ASAP7_75t_L g12054 ( 
.A(n_11678),
.Y(n_12054)
);

NAND2xp5_ASAP7_75t_L g12055 ( 
.A(n_11587),
.B(n_11297),
.Y(n_12055)
);

AND2x2_ASAP7_75t_L g12056 ( 
.A(n_11624),
.B(n_11191),
.Y(n_12056)
);

NAND2xp5_ASAP7_75t_SL g12057 ( 
.A(n_11566),
.B(n_11482),
.Y(n_12057)
);

INVx2_ASAP7_75t_L g12058 ( 
.A(n_11922),
.Y(n_12058)
);

INVx1_ASAP7_75t_L g12059 ( 
.A(n_11533),
.Y(n_12059)
);

AND2x4_ASAP7_75t_L g12060 ( 
.A(n_11566),
.B(n_11301),
.Y(n_12060)
);

INVx1_ASAP7_75t_L g12061 ( 
.A(n_11643),
.Y(n_12061)
);

INVx1_ASAP7_75t_L g12062 ( 
.A(n_11710),
.Y(n_12062)
);

INVx1_ASAP7_75t_SL g12063 ( 
.A(n_11550),
.Y(n_12063)
);

OR2x2_ASAP7_75t_L g12064 ( 
.A(n_11573),
.B(n_11376),
.Y(n_12064)
);

BUFx2_ASAP7_75t_L g12065 ( 
.A(n_11538),
.Y(n_12065)
);

AND2x2_ASAP7_75t_L g12066 ( 
.A(n_11716),
.B(n_11377),
.Y(n_12066)
);

NAND2xp5_ASAP7_75t_L g12067 ( 
.A(n_11587),
.B(n_11304),
.Y(n_12067)
);

BUFx2_ASAP7_75t_L g12068 ( 
.A(n_11511),
.Y(n_12068)
);

BUFx2_ASAP7_75t_L g12069 ( 
.A(n_11519),
.Y(n_12069)
);

AND2x2_ASAP7_75t_L g12070 ( 
.A(n_11538),
.B(n_11385),
.Y(n_12070)
);

AND2x4_ASAP7_75t_L g12071 ( 
.A(n_11541),
.B(n_11310),
.Y(n_12071)
);

INVx1_ASAP7_75t_L g12072 ( 
.A(n_11701),
.Y(n_12072)
);

INVx1_ASAP7_75t_L g12073 ( 
.A(n_11526),
.Y(n_12073)
);

AND2x2_ASAP7_75t_L g12074 ( 
.A(n_11807),
.B(n_11402),
.Y(n_12074)
);

INVx1_ASAP7_75t_L g12075 ( 
.A(n_11746),
.Y(n_12075)
);

INVx1_ASAP7_75t_L g12076 ( 
.A(n_11660),
.Y(n_12076)
);

INVx3_ASAP7_75t_L g12077 ( 
.A(n_11541),
.Y(n_12077)
);

HB1xp67_ASAP7_75t_L g12078 ( 
.A(n_11578),
.Y(n_12078)
);

INVx2_ASAP7_75t_L g12079 ( 
.A(n_11712),
.Y(n_12079)
);

NOR2xp33_ASAP7_75t_L g12080 ( 
.A(n_11629),
.B(n_11556),
.Y(n_12080)
);

NAND2xp5_ASAP7_75t_L g12081 ( 
.A(n_11883),
.B(n_11314),
.Y(n_12081)
);

NAND2xp5_ASAP7_75t_L g12082 ( 
.A(n_11658),
.B(n_11315),
.Y(n_12082)
);

INVx2_ASAP7_75t_L g12083 ( 
.A(n_11712),
.Y(n_12083)
);

INVx2_ASAP7_75t_L g12084 ( 
.A(n_11901),
.Y(n_12084)
);

INVx1_ASAP7_75t_L g12085 ( 
.A(n_11834),
.Y(n_12085)
);

AND2x2_ASAP7_75t_L g12086 ( 
.A(n_11891),
.B(n_11405),
.Y(n_12086)
);

AND2x2_ASAP7_75t_L g12087 ( 
.A(n_11517),
.B(n_11410),
.Y(n_12087)
);

INVx2_ASAP7_75t_L g12088 ( 
.A(n_11816),
.Y(n_12088)
);

AND2x4_ASAP7_75t_L g12089 ( 
.A(n_11658),
.B(n_11319),
.Y(n_12089)
);

AND2x4_ASAP7_75t_L g12090 ( 
.A(n_11590),
.B(n_11411),
.Y(n_12090)
);

AND2x2_ASAP7_75t_L g12091 ( 
.A(n_11809),
.B(n_11545),
.Y(n_12091)
);

NAND2xp5_ASAP7_75t_L g12092 ( 
.A(n_11637),
.B(n_11204),
.Y(n_12092)
);

AND2x4_ASAP7_75t_L g12093 ( 
.A(n_11590),
.B(n_11419),
.Y(n_12093)
);

INVx1_ASAP7_75t_L g12094 ( 
.A(n_11841),
.Y(n_12094)
);

INVx1_ASAP7_75t_L g12095 ( 
.A(n_11685),
.Y(n_12095)
);

INVx1_ASAP7_75t_L g12096 ( 
.A(n_11900),
.Y(n_12096)
);

INVx2_ASAP7_75t_L g12097 ( 
.A(n_11820),
.Y(n_12097)
);

INVx1_ASAP7_75t_L g12098 ( 
.A(n_11620),
.Y(n_12098)
);

NAND2xp5_ASAP7_75t_SL g12099 ( 
.A(n_11634),
.B(n_11106),
.Y(n_12099)
);

INVx2_ASAP7_75t_L g12100 ( 
.A(n_11786),
.Y(n_12100)
);

INVx1_ASAP7_75t_L g12101 ( 
.A(n_11627),
.Y(n_12101)
);

INVx3_ASAP7_75t_L g12102 ( 
.A(n_11848),
.Y(n_12102)
);

NAND2xp5_ASAP7_75t_L g12103 ( 
.A(n_11637),
.B(n_11218),
.Y(n_12103)
);

INVx1_ASAP7_75t_L g12104 ( 
.A(n_11706),
.Y(n_12104)
);

NAND2xp5_ASAP7_75t_L g12105 ( 
.A(n_11680),
.B(n_8901),
.Y(n_12105)
);

INVx2_ASAP7_75t_L g12106 ( 
.A(n_11786),
.Y(n_12106)
);

NAND2xp5_ASAP7_75t_L g12107 ( 
.A(n_11680),
.B(n_8912),
.Y(n_12107)
);

NAND2x1_ASAP7_75t_L g12108 ( 
.A(n_11878),
.B(n_11881),
.Y(n_12108)
);

NAND2x1_ASAP7_75t_L g12109 ( 
.A(n_11878),
.B(n_8912),
.Y(n_12109)
);

INVx1_ASAP7_75t_L g12110 ( 
.A(n_11818),
.Y(n_12110)
);

OR2x2_ASAP7_75t_L g12111 ( 
.A(n_11592),
.B(n_8499),
.Y(n_12111)
);

INVx2_ASAP7_75t_L g12112 ( 
.A(n_11797),
.Y(n_12112)
);

HB1xp67_ASAP7_75t_L g12113 ( 
.A(n_11808),
.Y(n_12113)
);

INVx1_ASAP7_75t_L g12114 ( 
.A(n_11528),
.Y(n_12114)
);

NOR2xp67_ASAP7_75t_L g12115 ( 
.A(n_11819),
.B(n_11537),
.Y(n_12115)
);

INVx1_ASAP7_75t_L g12116 ( 
.A(n_11536),
.Y(n_12116)
);

INVx1_ASAP7_75t_L g12117 ( 
.A(n_11543),
.Y(n_12117)
);

AND2x2_ASAP7_75t_L g12118 ( 
.A(n_11865),
.B(n_8501),
.Y(n_12118)
);

NAND2x1_ASAP7_75t_L g12119 ( 
.A(n_11881),
.B(n_8912),
.Y(n_12119)
);

AND2x2_ASAP7_75t_L g12120 ( 
.A(n_11864),
.B(n_8501),
.Y(n_12120)
);

NAND2xp5_ASAP7_75t_L g12121 ( 
.A(n_11711),
.B(n_8933),
.Y(n_12121)
);

AND2x2_ASAP7_75t_L g12122 ( 
.A(n_11811),
.B(n_8502),
.Y(n_12122)
);

INVx2_ASAP7_75t_L g12123 ( 
.A(n_11797),
.Y(n_12123)
);

AND2x2_ASAP7_75t_L g12124 ( 
.A(n_11602),
.B(n_8502),
.Y(n_12124)
);

INVx1_ASAP7_75t_L g12125 ( 
.A(n_11547),
.Y(n_12125)
);

AND2x4_ASAP7_75t_SL g12126 ( 
.A(n_11848),
.B(n_6847),
.Y(n_12126)
);

INVx1_ASAP7_75t_L g12127 ( 
.A(n_11832),
.Y(n_12127)
);

OAI21xp5_ASAP7_75t_L g12128 ( 
.A1(n_11648),
.A2(n_11625),
.B(n_11714),
.Y(n_12128)
);

INVx1_ASAP7_75t_L g12129 ( 
.A(n_11833),
.Y(n_12129)
);

AND2x2_ASAP7_75t_L g12130 ( 
.A(n_11555),
.B(n_8503),
.Y(n_12130)
);

INVx2_ASAP7_75t_L g12131 ( 
.A(n_11813),
.Y(n_12131)
);

NOR2xp33_ASAP7_75t_L g12132 ( 
.A(n_11586),
.B(n_11858),
.Y(n_12132)
);

AND2x2_ASAP7_75t_L g12133 ( 
.A(n_11656),
.B(n_11853),
.Y(n_12133)
);

INVx1_ASAP7_75t_L g12134 ( 
.A(n_11867),
.Y(n_12134)
);

NAND2xp5_ASAP7_75t_L g12135 ( 
.A(n_11711),
.B(n_8933),
.Y(n_12135)
);

OR2x2_ASAP7_75t_L g12136 ( 
.A(n_11640),
.B(n_8503),
.Y(n_12136)
);

NOR3xp33_ASAP7_75t_SL g12137 ( 
.A(n_11532),
.B(n_11473),
.C(n_10256),
.Y(n_12137)
);

NAND2xp5_ASAP7_75t_SL g12138 ( 
.A(n_11748),
.B(n_8097),
.Y(n_12138)
);

AND2x2_ASAP7_75t_L g12139 ( 
.A(n_11871),
.B(n_8504),
.Y(n_12139)
);

BUFx2_ASAP7_75t_L g12140 ( 
.A(n_11875),
.Y(n_12140)
);

OR2x2_ASAP7_75t_L g12141 ( 
.A(n_11665),
.B(n_8504),
.Y(n_12141)
);

INVx1_ASAP7_75t_L g12142 ( 
.A(n_11581),
.Y(n_12142)
);

INVx1_ASAP7_75t_L g12143 ( 
.A(n_11567),
.Y(n_12143)
);

INVx1_ASAP7_75t_L g12144 ( 
.A(n_11666),
.Y(n_12144)
);

AND2x2_ASAP7_75t_L g12145 ( 
.A(n_11817),
.B(n_8509),
.Y(n_12145)
);

NAND2xp5_ASAP7_75t_L g12146 ( 
.A(n_11750),
.B(n_11759),
.Y(n_12146)
);

BUFx2_ASAP7_75t_L g12147 ( 
.A(n_11735),
.Y(n_12147)
);

INVx1_ASAP7_75t_L g12148 ( 
.A(n_11670),
.Y(n_12148)
);

AND2x2_ASAP7_75t_L g12149 ( 
.A(n_11659),
.B(n_8509),
.Y(n_12149)
);

NAND2xp5_ASAP7_75t_L g12150 ( 
.A(n_11762),
.B(n_8933),
.Y(n_12150)
);

AND2x2_ASAP7_75t_L g12151 ( 
.A(n_11839),
.B(n_8519),
.Y(n_12151)
);

OR2x2_ASAP7_75t_L g12152 ( 
.A(n_11572),
.B(n_8519),
.Y(n_12152)
);

AND2x2_ASAP7_75t_L g12153 ( 
.A(n_11831),
.B(n_8523),
.Y(n_12153)
);

AND2x2_ASAP7_75t_L g12154 ( 
.A(n_11773),
.B(n_8523),
.Y(n_12154)
);

AND2x2_ASAP7_75t_L g12155 ( 
.A(n_11542),
.B(n_8525),
.Y(n_12155)
);

AND2x2_ASAP7_75t_L g12156 ( 
.A(n_11542),
.B(n_8525),
.Y(n_12156)
);

OR2x2_ASAP7_75t_L g12157 ( 
.A(n_11585),
.B(n_8531),
.Y(n_12157)
);

AND2x2_ASAP7_75t_L g12158 ( 
.A(n_11546),
.B(n_8531),
.Y(n_12158)
);

INVx1_ASAP7_75t_L g12159 ( 
.A(n_11614),
.Y(n_12159)
);

INVxp67_ASAP7_75t_L g12160 ( 
.A(n_11851),
.Y(n_12160)
);

AND2x2_ASAP7_75t_L g12161 ( 
.A(n_11546),
.B(n_8533),
.Y(n_12161)
);

NAND2x1p5_ASAP7_75t_L g12162 ( 
.A(n_11767),
.B(n_5673),
.Y(n_12162)
);

NAND2xp5_ASAP7_75t_L g12163 ( 
.A(n_11768),
.B(n_11775),
.Y(n_12163)
);

AND2x2_ASAP7_75t_L g12164 ( 
.A(n_11745),
.B(n_8533),
.Y(n_12164)
);

INVx5_ASAP7_75t_L g12165 ( 
.A(n_11813),
.Y(n_12165)
);

AND2x2_ASAP7_75t_SL g12166 ( 
.A(n_11728),
.B(n_10270),
.Y(n_12166)
);

AND2x2_ASAP7_75t_L g12167 ( 
.A(n_11705),
.B(n_8947),
.Y(n_12167)
);

AND2x2_ASAP7_75t_L g12168 ( 
.A(n_11718),
.B(n_8947),
.Y(n_12168)
);

AND2x2_ASAP7_75t_L g12169 ( 
.A(n_11724),
.B(n_8947),
.Y(n_12169)
);

AND2x4_ASAP7_75t_SL g12170 ( 
.A(n_11930),
.B(n_6847),
.Y(n_12170)
);

INVx1_ASAP7_75t_SL g12171 ( 
.A(n_11693),
.Y(n_12171)
);

NAND2xp5_ASAP7_75t_L g12172 ( 
.A(n_11827),
.B(n_8957),
.Y(n_12172)
);

OR2x2_ASAP7_75t_L g12173 ( 
.A(n_11594),
.B(n_11588),
.Y(n_12173)
);

HB1xp67_ASAP7_75t_L g12174 ( 
.A(n_11868),
.Y(n_12174)
);

INVx3_ASAP7_75t_L g12175 ( 
.A(n_11669),
.Y(n_12175)
);

NAND2xp5_ASAP7_75t_L g12176 ( 
.A(n_11649),
.B(n_8957),
.Y(n_12176)
);

AOI22xp33_ASAP7_75t_L g12177 ( 
.A1(n_11617),
.A2(n_10305),
.B1(n_10306),
.B2(n_10302),
.Y(n_12177)
);

AND2x2_ASAP7_75t_L g12178 ( 
.A(n_11882),
.B(n_8957),
.Y(n_12178)
);

AND2x4_ASAP7_75t_L g12179 ( 
.A(n_11721),
.B(n_8963),
.Y(n_12179)
);

INVx3_ASAP7_75t_L g12180 ( 
.A(n_11790),
.Y(n_12180)
);

NOR2xp67_ASAP7_75t_L g12181 ( 
.A(n_11603),
.B(n_8963),
.Y(n_12181)
);

INVx1_ASAP7_75t_L g12182 ( 
.A(n_11616),
.Y(n_12182)
);

INVx1_ASAP7_75t_L g12183 ( 
.A(n_11683),
.Y(n_12183)
);

INVx1_ASAP7_75t_L g12184 ( 
.A(n_11684),
.Y(n_12184)
);

NAND2xp5_ASAP7_75t_L g12185 ( 
.A(n_11910),
.B(n_8963),
.Y(n_12185)
);

NOR3xp33_ASAP7_75t_SL g12186 ( 
.A(n_11579),
.B(n_10273),
.C(n_10272),
.Y(n_12186)
);

AND2x2_ASAP7_75t_L g12187 ( 
.A(n_11631),
.B(n_8965),
.Y(n_12187)
);

INVx3_ASAP7_75t_L g12188 ( 
.A(n_11866),
.Y(n_12188)
);

HB1xp67_ASAP7_75t_L g12189 ( 
.A(n_11876),
.Y(n_12189)
);

INVx2_ASAP7_75t_L g12190 ( 
.A(n_11829),
.Y(n_12190)
);

AND2x2_ASAP7_75t_L g12191 ( 
.A(n_11709),
.B(n_8965),
.Y(n_12191)
);

INVx2_ASAP7_75t_L g12192 ( 
.A(n_11740),
.Y(n_12192)
);

INVx1_ASAP7_75t_L g12193 ( 
.A(n_11557),
.Y(n_12193)
);

AND2x4_ASAP7_75t_L g12194 ( 
.A(n_11726),
.B(n_8965),
.Y(n_12194)
);

INVx1_ASAP7_75t_L g12195 ( 
.A(n_11559),
.Y(n_12195)
);

NAND2xp5_ASAP7_75t_L g12196 ( 
.A(n_11568),
.B(n_9006),
.Y(n_12196)
);

NAND2xp5_ASAP7_75t_L g12197 ( 
.A(n_11571),
.B(n_9006),
.Y(n_12197)
);

AND2x2_ASAP7_75t_L g12198 ( 
.A(n_11898),
.B(n_9006),
.Y(n_12198)
);

INVx1_ASAP7_75t_L g12199 ( 
.A(n_11561),
.Y(n_12199)
);

INVx1_ASAP7_75t_L g12200 ( 
.A(n_11564),
.Y(n_12200)
);

AND2x2_ASAP7_75t_L g12201 ( 
.A(n_11633),
.B(n_9008),
.Y(n_12201)
);

AND2x2_ASAP7_75t_L g12202 ( 
.A(n_11636),
.B(n_9008),
.Y(n_12202)
);

AOI22xp5_ASAP7_75t_L g12203 ( 
.A1(n_11730),
.A2(n_10312),
.B1(n_10318),
.B2(n_10307),
.Y(n_12203)
);

AND2x2_ASAP7_75t_L g12204 ( 
.A(n_11715),
.B(n_9008),
.Y(n_12204)
);

INVx1_ASAP7_75t_L g12205 ( 
.A(n_11611),
.Y(n_12205)
);

INVx1_ASAP7_75t_L g12206 ( 
.A(n_11612),
.Y(n_12206)
);

INVx1_ASAP7_75t_L g12207 ( 
.A(n_11688),
.Y(n_12207)
);

NAND2xp5_ASAP7_75t_L g12208 ( 
.A(n_11576),
.B(n_9011),
.Y(n_12208)
);

INVx1_ASAP7_75t_L g12209 ( 
.A(n_11722),
.Y(n_12209)
);

INVx1_ASAP7_75t_L g12210 ( 
.A(n_11741),
.Y(n_12210)
);

AND2x2_ASAP7_75t_L g12211 ( 
.A(n_11917),
.B(n_9011),
.Y(n_12211)
);

AND2x2_ASAP7_75t_L g12212 ( 
.A(n_11507),
.B(n_9011),
.Y(n_12212)
);

NAND2xp5_ASAP7_75t_L g12213 ( 
.A(n_11580),
.B(n_8797),
.Y(n_12213)
);

NAND2xp5_ASAP7_75t_L g12214 ( 
.A(n_11589),
.B(n_11601),
.Y(n_12214)
);

OR2x2_ASAP7_75t_L g12215 ( 
.A(n_11628),
.B(n_9052),
.Y(n_12215)
);

AND2x2_ASAP7_75t_L g12216 ( 
.A(n_11512),
.B(n_7230),
.Y(n_12216)
);

AND2x2_ASAP7_75t_L g12217 ( 
.A(n_11880),
.B(n_7230),
.Y(n_12217)
);

INVx1_ASAP7_75t_L g12218 ( 
.A(n_11690),
.Y(n_12218)
);

AND2x2_ASAP7_75t_L g12219 ( 
.A(n_11903),
.B(n_7230),
.Y(n_12219)
);

HB1xp67_ASAP7_75t_L g12220 ( 
.A(n_11524),
.Y(n_12220)
);

OR2x2_ASAP7_75t_L g12221 ( 
.A(n_11913),
.B(n_9052),
.Y(n_12221)
);

AND2x2_ASAP7_75t_L g12222 ( 
.A(n_11919),
.B(n_7238),
.Y(n_12222)
);

HB1xp67_ASAP7_75t_L g12223 ( 
.A(n_11535),
.Y(n_12223)
);

NAND2xp5_ASAP7_75t_L g12224 ( 
.A(n_11672),
.B(n_8806),
.Y(n_12224)
);

INVx2_ASAP7_75t_L g12225 ( 
.A(n_11761),
.Y(n_12225)
);

AND2x2_ASAP7_75t_L g12226 ( 
.A(n_11890),
.B(n_7238),
.Y(n_12226)
);

NOR2x1_ASAP7_75t_L g12227 ( 
.A(n_11618),
.B(n_10275),
.Y(n_12227)
);

INVx1_ASAP7_75t_L g12228 ( 
.A(n_11860),
.Y(n_12228)
);

INVx4_ASAP7_75t_L g12229 ( 
.A(n_11554),
.Y(n_12229)
);

AND2x2_ASAP7_75t_L g12230 ( 
.A(n_11844),
.B(n_7238),
.Y(n_12230)
);

INVx1_ASAP7_75t_L g12231 ( 
.A(n_11704),
.Y(n_12231)
);

INVx1_ASAP7_75t_L g12232 ( 
.A(n_11671),
.Y(n_12232)
);

INVx1_ASAP7_75t_L g12233 ( 
.A(n_11838),
.Y(n_12233)
);

AND2x2_ASAP7_75t_L g12234 ( 
.A(n_11703),
.B(n_7252),
.Y(n_12234)
);

AND2x2_ASAP7_75t_L g12235 ( 
.A(n_11884),
.B(n_7252),
.Y(n_12235)
);

AOI22xp5_ASAP7_75t_L g12236 ( 
.A1(n_11874),
.A2(n_10326),
.B1(n_10335),
.B2(n_10334),
.Y(n_12236)
);

INVx1_ASAP7_75t_L g12237 ( 
.A(n_11845),
.Y(n_12237)
);

INVx1_ASAP7_75t_L g12238 ( 
.A(n_11779),
.Y(n_12238)
);

AND2x2_ASAP7_75t_L g12239 ( 
.A(n_11727),
.B(n_7252),
.Y(n_12239)
);

AND2x2_ASAP7_75t_L g12240 ( 
.A(n_11802),
.B(n_9052),
.Y(n_12240)
);

OR2x2_ASAP7_75t_L g12241 ( 
.A(n_11738),
.B(n_9071),
.Y(n_12241)
);

BUFx3_ASAP7_75t_L g12242 ( 
.A(n_11931),
.Y(n_12242)
);

AND2x2_ASAP7_75t_L g12243 ( 
.A(n_11732),
.B(n_9071),
.Y(n_12243)
);

BUFx3_ASAP7_75t_L g12244 ( 
.A(n_11936),
.Y(n_12244)
);

NAND2xp5_ASAP7_75t_L g12245 ( 
.A(n_11677),
.B(n_8806),
.Y(n_12245)
);

NAND2xp5_ASAP7_75t_L g12246 ( 
.A(n_11679),
.B(n_8807),
.Y(n_12246)
);

AND2x2_ASAP7_75t_L g12247 ( 
.A(n_11733),
.B(n_9071),
.Y(n_12247)
);

OR2x2_ASAP7_75t_L g12248 ( 
.A(n_11525),
.B(n_9101),
.Y(n_12248)
);

AND2x2_ASAP7_75t_L g12249 ( 
.A(n_11753),
.B(n_9101),
.Y(n_12249)
);

INVx1_ASAP7_75t_L g12250 ( 
.A(n_11548),
.Y(n_12250)
);

AND2x4_ASAP7_75t_L g12251 ( 
.A(n_11763),
.B(n_9101),
.Y(n_12251)
);

HB1xp67_ASAP7_75t_L g12252 ( 
.A(n_11558),
.Y(n_12252)
);

INVx1_ASAP7_75t_SL g12253 ( 
.A(n_11720),
.Y(n_12253)
);

AND2x2_ASAP7_75t_L g12254 ( 
.A(n_11781),
.B(n_9085),
.Y(n_12254)
);

INVx2_ASAP7_75t_L g12255 ( 
.A(n_11894),
.Y(n_12255)
);

NOR2xp33_ASAP7_75t_L g12256 ( 
.A(n_11565),
.B(n_7647),
.Y(n_12256)
);

NOR2xp33_ASAP7_75t_SL g12257 ( 
.A(n_11731),
.B(n_7234),
.Y(n_12257)
);

INVx2_ASAP7_75t_L g12258 ( 
.A(n_11826),
.Y(n_12258)
);

AND2x2_ASAP7_75t_L g12259 ( 
.A(n_11906),
.B(n_9085),
.Y(n_12259)
);

AND2x2_ASAP7_75t_L g12260 ( 
.A(n_11869),
.B(n_9102),
.Y(n_12260)
);

OR2x2_ASAP7_75t_L g12261 ( 
.A(n_11552),
.B(n_11747),
.Y(n_12261)
);

AND2x2_ASAP7_75t_L g12262 ( 
.A(n_11828),
.B(n_9102),
.Y(n_12262)
);

OR2x2_ASAP7_75t_L g12263 ( 
.A(n_11695),
.B(n_7875),
.Y(n_12263)
);

AND2x4_ASAP7_75t_SL g12264 ( 
.A(n_11574),
.B(n_6984),
.Y(n_12264)
);

AND2x2_ASAP7_75t_L g12265 ( 
.A(n_11823),
.B(n_8824),
.Y(n_12265)
);

INVx1_ASAP7_75t_L g12266 ( 
.A(n_11687),
.Y(n_12266)
);

INVx1_ASAP7_75t_L g12267 ( 
.A(n_11696),
.Y(n_12267)
);

INVx1_ASAP7_75t_L g12268 ( 
.A(n_11697),
.Y(n_12268)
);

AND2x4_ASAP7_75t_L g12269 ( 
.A(n_11575),
.B(n_11591),
.Y(n_12269)
);

INVx2_ASAP7_75t_L g12270 ( 
.A(n_11596),
.Y(n_12270)
);

INVx4_ASAP7_75t_L g12271 ( 
.A(n_11523),
.Y(n_12271)
);

NAND2xp5_ASAP7_75t_L g12272 ( 
.A(n_11801),
.B(n_8807),
.Y(n_12272)
);

AND2x4_ASAP7_75t_L g12273 ( 
.A(n_11529),
.B(n_8824),
.Y(n_12273)
);

INVx2_ASAP7_75t_L g12274 ( 
.A(n_11756),
.Y(n_12274)
);

INVx1_ASAP7_75t_L g12275 ( 
.A(n_11700),
.Y(n_12275)
);

INVx1_ASAP7_75t_L g12276 ( 
.A(n_11702),
.Y(n_12276)
);

INVx1_ASAP7_75t_L g12277 ( 
.A(n_11821),
.Y(n_12277)
);

AND2x2_ASAP7_75t_L g12278 ( 
.A(n_11764),
.B(n_6642),
.Y(n_12278)
);

OR2x2_ASAP7_75t_L g12279 ( 
.A(n_11873),
.B(n_7910),
.Y(n_12279)
);

AND2x2_ASAP7_75t_L g12280 ( 
.A(n_11766),
.B(n_6642),
.Y(n_12280)
);

INVx1_ASAP7_75t_L g12281 ( 
.A(n_11776),
.Y(n_12281)
);

INVx2_ASAP7_75t_SL g12282 ( 
.A(n_11847),
.Y(n_12282)
);

AND2x2_ASAP7_75t_L g12283 ( 
.A(n_11770),
.B(n_8653),
.Y(n_12283)
);

INVx1_ASAP7_75t_L g12284 ( 
.A(n_11800),
.Y(n_12284)
);

AND2x4_ASAP7_75t_L g12285 ( 
.A(n_11531),
.B(n_9673),
.Y(n_12285)
);

AND2x2_ASAP7_75t_L g12286 ( 
.A(n_11771),
.B(n_8653),
.Y(n_12286)
);

NAND2xp5_ASAP7_75t_L g12287 ( 
.A(n_11812),
.B(n_8810),
.Y(n_12287)
);

NAND2xp5_ASAP7_75t_L g12288 ( 
.A(n_11862),
.B(n_8810),
.Y(n_12288)
);

INVx1_ASAP7_75t_L g12289 ( 
.A(n_11806),
.Y(n_12289)
);

OR2x2_ASAP7_75t_L g12290 ( 
.A(n_11734),
.B(n_7942),
.Y(n_12290)
);

INVx1_ASAP7_75t_L g12291 ( 
.A(n_11857),
.Y(n_12291)
);

NOR2x1_ASAP7_75t_L g12292 ( 
.A(n_11857),
.B(n_10281),
.Y(n_12292)
);

BUFx2_ASAP7_75t_L g12293 ( 
.A(n_11756),
.Y(n_12293)
);

OR2x2_ASAP7_75t_L g12294 ( 
.A(n_11674),
.B(n_7942),
.Y(n_12294)
);

OR2x2_ASAP7_75t_L g12295 ( 
.A(n_11676),
.B(n_11650),
.Y(n_12295)
);

NOR2xp33_ASAP7_75t_L g12296 ( 
.A(n_11647),
.B(n_7647),
.Y(n_12296)
);

INVx2_ASAP7_75t_L g12297 ( 
.A(n_11769),
.Y(n_12297)
);

INVx3_ASAP7_75t_L g12298 ( 
.A(n_11866),
.Y(n_12298)
);

INVx1_ASAP7_75t_L g12299 ( 
.A(n_11888),
.Y(n_12299)
);

HB1xp67_ASAP7_75t_L g12300 ( 
.A(n_11725),
.Y(n_12300)
);

NAND2xp5_ASAP7_75t_L g12301 ( 
.A(n_11657),
.B(n_8818),
.Y(n_12301)
);

NAND2xp5_ASAP7_75t_L g12302 ( 
.A(n_11663),
.B(n_8818),
.Y(n_12302)
);

INVx1_ASAP7_75t_L g12303 ( 
.A(n_11888),
.Y(n_12303)
);

INVx1_ASAP7_75t_L g12304 ( 
.A(n_11927),
.Y(n_12304)
);

AND2x4_ASAP7_75t_L g12305 ( 
.A(n_11803),
.B(n_11796),
.Y(n_12305)
);

OR2x2_ASAP7_75t_L g12306 ( 
.A(n_11842),
.B(n_7966),
.Y(n_12306)
);

INVx1_ASAP7_75t_L g12307 ( 
.A(n_11928),
.Y(n_12307)
);

INVx1_ASAP7_75t_L g12308 ( 
.A(n_11760),
.Y(n_12308)
);

INVx2_ASAP7_75t_L g12309 ( 
.A(n_11769),
.Y(n_12309)
);

OR2x2_ASAP7_75t_L g12310 ( 
.A(n_11846),
.B(n_7966),
.Y(n_12310)
);

OR2x2_ASAP7_75t_L g12311 ( 
.A(n_11896),
.B(n_7972),
.Y(n_12311)
);

INVx2_ASAP7_75t_L g12312 ( 
.A(n_11889),
.Y(n_12312)
);

NAND2xp5_ASAP7_75t_L g12313 ( 
.A(n_11852),
.B(n_8819),
.Y(n_12313)
);

INVx1_ASAP7_75t_L g12314 ( 
.A(n_11784),
.Y(n_12314)
);

OR2x6_ASAP7_75t_L g12315 ( 
.A(n_11641),
.B(n_7697),
.Y(n_12315)
);

AND2x2_ASAP7_75t_L g12316 ( 
.A(n_11792),
.B(n_6568),
.Y(n_12316)
);

AND2x2_ASAP7_75t_L g12317 ( 
.A(n_11794),
.B(n_6568),
.Y(n_12317)
);

NAND2xp5_ASAP7_75t_L g12318 ( 
.A(n_11939),
.B(n_8819),
.Y(n_12318)
);

INVx1_ASAP7_75t_L g12319 ( 
.A(n_11837),
.Y(n_12319)
);

NAND2xp5_ASAP7_75t_L g12320 ( 
.A(n_11920),
.B(n_8820),
.Y(n_12320)
);

INVx3_ASAP7_75t_SL g12321 ( 
.A(n_11645),
.Y(n_12321)
);

OR2x2_ASAP7_75t_L g12322 ( 
.A(n_11897),
.B(n_7980),
.Y(n_12322)
);

INVx1_ASAP7_75t_L g12323 ( 
.A(n_11785),
.Y(n_12323)
);

AND2x2_ASAP7_75t_L g12324 ( 
.A(n_11968),
.B(n_11870),
.Y(n_12324)
);

INVx3_ASAP7_75t_L g12325 ( 
.A(n_11966),
.Y(n_12325)
);

AND2x2_ASAP7_75t_L g12326 ( 
.A(n_11971),
.B(n_11798),
.Y(n_12326)
);

AOI22xp5_ASAP7_75t_L g12327 ( 
.A1(n_12019),
.A2(n_11719),
.B1(n_11911),
.B2(n_11736),
.Y(n_12327)
);

BUFx3_ASAP7_75t_L g12328 ( 
.A(n_12065),
.Y(n_12328)
);

INVx1_ASAP7_75t_L g12329 ( 
.A(n_12068),
.Y(n_12329)
);

OR2x2_ASAP7_75t_L g12330 ( 
.A(n_12016),
.B(n_11739),
.Y(n_12330)
);

INVx2_ASAP7_75t_L g12331 ( 
.A(n_12102),
.Y(n_12331)
);

INVx1_ASAP7_75t_L g12332 ( 
.A(n_12068),
.Y(n_12332)
);

OR2x2_ASAP7_75t_L g12333 ( 
.A(n_12037),
.B(n_11755),
.Y(n_12333)
);

AND2x2_ASAP7_75t_L g12334 ( 
.A(n_11948),
.B(n_11799),
.Y(n_12334)
);

INVx2_ASAP7_75t_L g12335 ( 
.A(n_12077),
.Y(n_12335)
);

INVx1_ASAP7_75t_L g12336 ( 
.A(n_12069),
.Y(n_12336)
);

INVx2_ASAP7_75t_L g12337 ( 
.A(n_12007),
.Y(n_12337)
);

NAND2xp5_ASAP7_75t_L g12338 ( 
.A(n_11947),
.B(n_12030),
.Y(n_12338)
);

INVx1_ASAP7_75t_L g12339 ( 
.A(n_12069),
.Y(n_12339)
);

OR2x2_ASAP7_75t_L g12340 ( 
.A(n_12063),
.B(n_11895),
.Y(n_12340)
);

INVx2_ASAP7_75t_SL g12341 ( 
.A(n_12002),
.Y(n_12341)
);

INVx1_ASAP7_75t_L g12342 ( 
.A(n_12043),
.Y(n_12342)
);

INVx1_ASAP7_75t_L g12343 ( 
.A(n_11954),
.Y(n_12343)
);

INVx1_ASAP7_75t_L g12344 ( 
.A(n_11956),
.Y(n_12344)
);

OR2x2_ASAP7_75t_L g12345 ( 
.A(n_12171),
.B(n_11788),
.Y(n_12345)
);

AND2x2_ASAP7_75t_L g12346 ( 
.A(n_11970),
.B(n_11886),
.Y(n_12346)
);

OR2x2_ASAP7_75t_L g12347 ( 
.A(n_11965),
.B(n_11791),
.Y(n_12347)
);

NOR3xp33_ASAP7_75t_L g12348 ( 
.A(n_12128),
.B(n_11941),
.C(n_11774),
.Y(n_12348)
);

INVx1_ASAP7_75t_L g12349 ( 
.A(n_12140),
.Y(n_12349)
);

INVx2_ASAP7_75t_L g12350 ( 
.A(n_11947),
.Y(n_12350)
);

NAND2xp5_ASAP7_75t_L g12351 ( 
.A(n_11975),
.B(n_11907),
.Y(n_12351)
);

AND2x2_ASAP7_75t_L g12352 ( 
.A(n_11985),
.B(n_11908),
.Y(n_12352)
);

INVxp67_ASAP7_75t_L g12353 ( 
.A(n_11976),
.Y(n_12353)
);

INVx2_ASAP7_75t_SL g12354 ( 
.A(n_11991),
.Y(n_12354)
);

INVx1_ASAP7_75t_L g12355 ( 
.A(n_12140),
.Y(n_12355)
);

NAND2xp5_ASAP7_75t_L g12356 ( 
.A(n_11999),
.B(n_12071),
.Y(n_12356)
);

INVx1_ASAP7_75t_L g12357 ( 
.A(n_12071),
.Y(n_12357)
);

INVxp67_ASAP7_75t_L g12358 ( 
.A(n_12034),
.Y(n_12358)
);

INVx2_ASAP7_75t_L g12359 ( 
.A(n_12165),
.Y(n_12359)
);

INVx4_ASAP7_75t_L g12360 ( 
.A(n_12175),
.Y(n_12360)
);

INVx1_ASAP7_75t_L g12361 ( 
.A(n_12003),
.Y(n_12361)
);

AND2x4_ASAP7_75t_L g12362 ( 
.A(n_12004),
.B(n_11667),
.Y(n_12362)
);

INVx1_ASAP7_75t_L g12363 ( 
.A(n_11969),
.Y(n_12363)
);

OAI211xp5_ASAP7_75t_SL g12364 ( 
.A1(n_12137),
.A2(n_11855),
.B(n_11938),
.C(n_11778),
.Y(n_12364)
);

AND2x2_ASAP7_75t_L g12365 ( 
.A(n_12009),
.B(n_11749),
.Y(n_12365)
);

INVx1_ASAP7_75t_SL g12366 ( 
.A(n_12091),
.Y(n_12366)
);

AND2x4_ASAP7_75t_L g12367 ( 
.A(n_12133),
.B(n_11708),
.Y(n_12367)
);

BUFx2_ASAP7_75t_L g12368 ( 
.A(n_12046),
.Y(n_12368)
);

AND2x2_ASAP7_75t_L g12369 ( 
.A(n_11995),
.B(n_11752),
.Y(n_12369)
);

INVx2_ASAP7_75t_L g12370 ( 
.A(n_12165),
.Y(n_12370)
);

HB1xp67_ASAP7_75t_L g12371 ( 
.A(n_12165),
.Y(n_12371)
);

AND2x2_ASAP7_75t_L g12372 ( 
.A(n_11996),
.B(n_11777),
.Y(n_12372)
);

OR2x2_ASAP7_75t_L g12373 ( 
.A(n_12173),
.B(n_11863),
.Y(n_12373)
);

AND2x2_ASAP7_75t_L g12374 ( 
.A(n_11961),
.B(n_11793),
.Y(n_12374)
);

INVxp67_ASAP7_75t_L g12375 ( 
.A(n_12092),
.Y(n_12375)
);

NOR3xp33_ASAP7_75t_SL g12376 ( 
.A(n_11982),
.B(n_11795),
.C(n_11822),
.Y(n_12376)
);

BUFx2_ASAP7_75t_SL g12377 ( 
.A(n_12022),
.Y(n_12377)
);

NAND2x1p5_ASAP7_75t_L g12378 ( 
.A(n_11949),
.B(n_11824),
.Y(n_12378)
);

AND2x4_ASAP7_75t_L g12379 ( 
.A(n_12090),
.B(n_12093),
.Y(n_12379)
);

INVx1_ASAP7_75t_L g12380 ( 
.A(n_12223),
.Y(n_12380)
);

INVx2_ASAP7_75t_L g12381 ( 
.A(n_12242),
.Y(n_12381)
);

AOI22xp33_ASAP7_75t_SL g12382 ( 
.A1(n_12166),
.A2(n_11902),
.B1(n_12027),
.B2(n_11950),
.Y(n_12382)
);

OR2x6_ASAP7_75t_L g12383 ( 
.A(n_12084),
.B(n_11825),
.Y(n_12383)
);

AND2x2_ASAP7_75t_L g12384 ( 
.A(n_12006),
.B(n_11815),
.Y(n_12384)
);

INVx1_ASAP7_75t_L g12385 ( 
.A(n_12252),
.Y(n_12385)
);

INVx1_ASAP7_75t_SL g12386 ( 
.A(n_12047),
.Y(n_12386)
);

NAND2xp5_ASAP7_75t_L g12387 ( 
.A(n_12025),
.B(n_12033),
.Y(n_12387)
);

INVx2_ASAP7_75t_L g12388 ( 
.A(n_12244),
.Y(n_12388)
);

INVx2_ASAP7_75t_L g12389 ( 
.A(n_12064),
.Y(n_12389)
);

AND2x2_ASAP7_75t_L g12390 ( 
.A(n_12066),
.B(n_11940),
.Y(n_12390)
);

INVx2_ASAP7_75t_L g12391 ( 
.A(n_12035),
.Y(n_12391)
);

NAND2xp5_ASAP7_75t_L g12392 ( 
.A(n_12035),
.B(n_11943),
.Y(n_12392)
);

AND2x2_ASAP7_75t_L g12393 ( 
.A(n_12028),
.B(n_11849),
.Y(n_12393)
);

AND2x2_ASAP7_75t_L g12394 ( 
.A(n_12086),
.B(n_11915),
.Y(n_12394)
);

INVx1_ASAP7_75t_L g12395 ( 
.A(n_12074),
.Y(n_12395)
);

AND2x2_ASAP7_75t_L g12396 ( 
.A(n_12023),
.B(n_11944),
.Y(n_12396)
);

AND2x2_ASAP7_75t_L g12397 ( 
.A(n_12031),
.B(n_11835),
.Y(n_12397)
);

NAND2xp5_ASAP7_75t_L g12398 ( 
.A(n_12060),
.B(n_11854),
.Y(n_12398)
);

AOI22xp33_ASAP7_75t_L g12399 ( 
.A1(n_12000),
.A2(n_11932),
.B1(n_11751),
.B2(n_11924),
.Y(n_12399)
);

AOI22xp33_ASAP7_75t_SL g12400 ( 
.A1(n_11946),
.A2(n_11918),
.B1(n_11912),
.B2(n_11942),
.Y(n_12400)
);

NAND2xp5_ASAP7_75t_L g12401 ( 
.A(n_12060),
.B(n_11854),
.Y(n_12401)
);

INVx3_ASAP7_75t_L g12402 ( 
.A(n_12090),
.Y(n_12402)
);

AND2x2_ASAP7_75t_L g12403 ( 
.A(n_12020),
.B(n_11836),
.Y(n_12403)
);

CKINVDCx5p33_ASAP7_75t_R g12404 ( 
.A(n_11951),
.Y(n_12404)
);

AND2x4_ASAP7_75t_L g12405 ( 
.A(n_12093),
.B(n_11935),
.Y(n_12405)
);

OR2x2_ASAP7_75t_L g12406 ( 
.A(n_12110),
.B(n_11804),
.Y(n_12406)
);

OAI211xp5_ASAP7_75t_L g12407 ( 
.A1(n_12015),
.A2(n_12057),
.B(n_12080),
.C(n_12078),
.Y(n_12407)
);

AND2x2_ASAP7_75t_L g12408 ( 
.A(n_11974),
.B(n_11840),
.Y(n_12408)
);

INVx1_ASAP7_75t_SL g12409 ( 
.A(n_12040),
.Y(n_12409)
);

NAND2xp5_ASAP7_75t_L g12410 ( 
.A(n_12010),
.B(n_11805),
.Y(n_12410)
);

INVx1_ASAP7_75t_L g12411 ( 
.A(n_12070),
.Y(n_12411)
);

AND2x2_ASAP7_75t_L g12412 ( 
.A(n_11952),
.B(n_11843),
.Y(n_12412)
);

AND2x2_ASAP7_75t_L g12413 ( 
.A(n_12032),
.B(n_11856),
.Y(n_12413)
);

AND2x2_ASAP7_75t_L g12414 ( 
.A(n_12056),
.B(n_11861),
.Y(n_12414)
);

NAND2xp5_ASAP7_75t_L g12415 ( 
.A(n_12089),
.B(n_11810),
.Y(n_12415)
);

AND2x4_ASAP7_75t_L g12416 ( 
.A(n_12089),
.B(n_11937),
.Y(n_12416)
);

AOI22xp33_ASAP7_75t_L g12417 ( 
.A1(n_12103),
.A2(n_8851),
.B1(n_8899),
.B2(n_9055),
.Y(n_12417)
);

OR2x2_ASAP7_75t_L g12418 ( 
.A(n_12190),
.B(n_11830),
.Y(n_12418)
);

INVx1_ASAP7_75t_L g12419 ( 
.A(n_11955),
.Y(n_12419)
);

INVx2_ASAP7_75t_L g12420 ( 
.A(n_12293),
.Y(n_12420)
);

NAND2xp5_ASAP7_75t_L g12421 ( 
.A(n_12011),
.B(n_11872),
.Y(n_12421)
);

INVx1_ASAP7_75t_L g12422 ( 
.A(n_12292),
.Y(n_12422)
);

INVx2_ASAP7_75t_L g12423 ( 
.A(n_11967),
.Y(n_12423)
);

NAND2xp5_ASAP7_75t_L g12424 ( 
.A(n_12029),
.B(n_11877),
.Y(n_12424)
);

AND2x2_ASAP7_75t_L g12425 ( 
.A(n_11945),
.B(n_12209),
.Y(n_12425)
);

NAND2x1p5_ASAP7_75t_L g12426 ( 
.A(n_11949),
.B(n_11879),
.Y(n_12426)
);

INVx1_ASAP7_75t_L g12427 ( 
.A(n_12147),
.Y(n_12427)
);

OR2x2_ASAP7_75t_L g12428 ( 
.A(n_12210),
.B(n_11885),
.Y(n_12428)
);

INVx2_ASAP7_75t_L g12429 ( 
.A(n_11953),
.Y(n_12429)
);

INVxp33_ASAP7_75t_L g12430 ( 
.A(n_11978),
.Y(n_12430)
);

INVx1_ASAP7_75t_L g12431 ( 
.A(n_12147),
.Y(n_12431)
);

NAND2xp5_ASAP7_75t_L g12432 ( 
.A(n_12253),
.B(n_11887),
.Y(n_12432)
);

NAND2xp5_ASAP7_75t_L g12433 ( 
.A(n_11953),
.B(n_11892),
.Y(n_12433)
);

AND2x2_ASAP7_75t_L g12434 ( 
.A(n_12024),
.B(n_11893),
.Y(n_12434)
);

AND2x2_ASAP7_75t_L g12435 ( 
.A(n_12058),
.B(n_11909),
.Y(n_12435)
);

OR2x2_ASAP7_75t_L g12436 ( 
.A(n_12075),
.B(n_11914),
.Y(n_12436)
);

INVx1_ASAP7_75t_L g12437 ( 
.A(n_11981),
.Y(n_12437)
);

INVx1_ASAP7_75t_L g12438 ( 
.A(n_11983),
.Y(n_12438)
);

NOR3xp33_ASAP7_75t_L g12439 ( 
.A(n_12099),
.B(n_11926),
.C(n_11925),
.Y(n_12439)
);

INVx1_ASAP7_75t_L g12440 ( 
.A(n_11973),
.Y(n_12440)
);

AND2x4_ASAP7_75t_L g12441 ( 
.A(n_12269),
.B(n_11929),
.Y(n_12441)
);

INVx2_ASAP7_75t_L g12442 ( 
.A(n_11957),
.Y(n_12442)
);

NAND2xp5_ASAP7_75t_L g12443 ( 
.A(n_12144),
.B(n_11934),
.Y(n_12443)
);

AND2x2_ASAP7_75t_L g12444 ( 
.A(n_11987),
.B(n_11899),
.Y(n_12444)
);

AOI32xp33_ASAP7_75t_L g12445 ( 
.A1(n_11963),
.A2(n_11904),
.A3(n_11905),
.B1(n_11923),
.B2(n_11921),
.Y(n_12445)
);

AOI211xp5_ASAP7_75t_L g12446 ( 
.A1(n_12115),
.A2(n_8551),
.B(n_8949),
.C(n_8943),
.Y(n_12446)
);

INVxp67_ASAP7_75t_SL g12447 ( 
.A(n_12021),
.Y(n_12447)
);

INVx1_ASAP7_75t_L g12448 ( 
.A(n_11977),
.Y(n_12448)
);

INVx1_ASAP7_75t_L g12449 ( 
.A(n_12113),
.Y(n_12449)
);

HB1xp67_ASAP7_75t_L g12450 ( 
.A(n_12291),
.Y(n_12450)
);

BUFx3_ASAP7_75t_L g12451 ( 
.A(n_12269),
.Y(n_12451)
);

NAND2xp5_ASAP7_75t_L g12452 ( 
.A(n_12148),
.B(n_8820),
.Y(n_12452)
);

NAND2xp5_ASAP7_75t_L g12453 ( 
.A(n_12062),
.B(n_8822),
.Y(n_12453)
);

INVx1_ASAP7_75t_L g12454 ( 
.A(n_12299),
.Y(n_12454)
);

AND2x4_ASAP7_75t_L g12455 ( 
.A(n_11979),
.B(n_12229),
.Y(n_12455)
);

INVx1_ASAP7_75t_L g12456 ( 
.A(n_12303),
.Y(n_12456)
);

INVx2_ASAP7_75t_L g12457 ( 
.A(n_11959),
.Y(n_12457)
);

NAND2xp5_ASAP7_75t_L g12458 ( 
.A(n_12143),
.B(n_8822),
.Y(n_12458)
);

INVx1_ASAP7_75t_L g12459 ( 
.A(n_11989),
.Y(n_12459)
);

INVx2_ASAP7_75t_L g12460 ( 
.A(n_12188),
.Y(n_12460)
);

OR2x2_ASAP7_75t_L g12461 ( 
.A(n_12026),
.B(n_9152),
.Y(n_12461)
);

NOR2xp33_ASAP7_75t_L g12462 ( 
.A(n_12271),
.B(n_8825),
.Y(n_12462)
);

NAND2xp5_ASAP7_75t_L g12463 ( 
.A(n_12017),
.B(n_8825),
.Y(n_12463)
);

INVx2_ASAP7_75t_L g12464 ( 
.A(n_12298),
.Y(n_12464)
);

BUFx3_ASAP7_75t_L g12465 ( 
.A(n_12012),
.Y(n_12465)
);

INVxp67_ASAP7_75t_SL g12466 ( 
.A(n_12045),
.Y(n_12466)
);

AND2x2_ASAP7_75t_L g12467 ( 
.A(n_12061),
.B(n_9162),
.Y(n_12467)
);

AND2x2_ASAP7_75t_L g12468 ( 
.A(n_12039),
.B(n_12041),
.Y(n_12468)
);

NAND2xp5_ASAP7_75t_SL g12469 ( 
.A(n_11979),
.B(n_9676),
.Y(n_12469)
);

AOI21xp5_ASAP7_75t_L g12470 ( 
.A1(n_12108),
.A2(n_9162),
.B(n_8743),
.Y(n_12470)
);

NOR2x1_ASAP7_75t_L g12471 ( 
.A(n_11988),
.B(n_8826),
.Y(n_12471)
);

AND2x2_ASAP7_75t_L g12472 ( 
.A(n_12076),
.B(n_9679),
.Y(n_12472)
);

AND2x2_ASAP7_75t_L g12473 ( 
.A(n_12095),
.B(n_9693),
.Y(n_12473)
);

INVx2_ASAP7_75t_L g12474 ( 
.A(n_12155),
.Y(n_12474)
);

AND2x2_ASAP7_75t_L g12475 ( 
.A(n_12142),
.B(n_12216),
.Y(n_12475)
);

AND2x2_ASAP7_75t_L g12476 ( 
.A(n_12180),
.B(n_9695),
.Y(n_12476)
);

INVx1_ASAP7_75t_L g12477 ( 
.A(n_12055),
.Y(n_12477)
);

OR2x2_ASAP7_75t_L g12478 ( 
.A(n_12001),
.B(n_8826),
.Y(n_12478)
);

AND2x2_ASAP7_75t_L g12479 ( 
.A(n_12239),
.B(n_6568),
.Y(n_12479)
);

AND2x2_ASAP7_75t_L g12480 ( 
.A(n_12234),
.B(n_12258),
.Y(n_12480)
);

AOI22xp33_ASAP7_75t_L g12481 ( 
.A1(n_11972),
.A2(n_8899),
.B1(n_9077),
.B2(n_9055),
.Y(n_12481)
);

NAND2xp5_ASAP7_75t_L g12482 ( 
.A(n_12149),
.B(n_8827),
.Y(n_12482)
);

OR2x2_ASAP7_75t_L g12483 ( 
.A(n_11962),
.B(n_8827),
.Y(n_12483)
);

AND2x2_ASAP7_75t_L g12484 ( 
.A(n_12315),
.B(n_12321),
.Y(n_12484)
);

OR2x2_ASAP7_75t_L g12485 ( 
.A(n_12067),
.B(n_8828),
.Y(n_12485)
);

INVx1_ASAP7_75t_L g12486 ( 
.A(n_12082),
.Y(n_12486)
);

OR2x2_ASAP7_75t_L g12487 ( 
.A(n_11960),
.B(n_8828),
.Y(n_12487)
);

INVx2_ASAP7_75t_L g12488 ( 
.A(n_12156),
.Y(n_12488)
);

INVx2_ASAP7_75t_L g12489 ( 
.A(n_12158),
.Y(n_12489)
);

AND2x2_ASAP7_75t_L g12490 ( 
.A(n_12315),
.B(n_6568),
.Y(n_12490)
);

INVx2_ASAP7_75t_L g12491 ( 
.A(n_12161),
.Y(n_12491)
);

AOI22xp33_ASAP7_75t_L g12492 ( 
.A1(n_11986),
.A2(n_9077),
.B1(n_8743),
.B2(n_8974),
.Y(n_12492)
);

INVx1_ASAP7_75t_L g12493 ( 
.A(n_12087),
.Y(n_12493)
);

HB1xp67_ASAP7_75t_L g12494 ( 
.A(n_12181),
.Y(n_12494)
);

AND2x2_ASAP7_75t_L g12495 ( 
.A(n_12255),
.B(n_12122),
.Y(n_12495)
);

INVx1_ASAP7_75t_L g12496 ( 
.A(n_12220),
.Y(n_12496)
);

NOR2xp33_ASAP7_75t_L g12497 ( 
.A(n_12257),
.B(n_8962),
.Y(n_12497)
);

INVx1_ASAP7_75t_L g12498 ( 
.A(n_12053),
.Y(n_12498)
);

NAND2xp5_ASAP7_75t_L g12499 ( 
.A(n_12304),
.B(n_8962),
.Y(n_12499)
);

INVx1_ASAP7_75t_L g12500 ( 
.A(n_12131),
.Y(n_12500)
);

INVx1_ASAP7_75t_L g12501 ( 
.A(n_12261),
.Y(n_12501)
);

AND2x2_ASAP7_75t_L g12502 ( 
.A(n_12120),
.B(n_12008),
.Y(n_12502)
);

NOR2xp33_ASAP7_75t_L g12503 ( 
.A(n_12038),
.B(n_8974),
.Y(n_12503)
);

AND2x2_ASAP7_75t_L g12504 ( 
.A(n_12014),
.B(n_6568),
.Y(n_12504)
);

AND2x2_ASAP7_75t_L g12505 ( 
.A(n_12073),
.B(n_6568),
.Y(n_12505)
);

HB1xp67_ASAP7_75t_L g12506 ( 
.A(n_12174),
.Y(n_12506)
);

AOI22xp33_ASAP7_75t_L g12507 ( 
.A1(n_12088),
.A2(n_9077),
.B1(n_8743),
.B2(n_8982),
.Y(n_12507)
);

AND2x2_ASAP7_75t_L g12508 ( 
.A(n_12219),
.B(n_7066),
.Y(n_12508)
);

HB1xp67_ASAP7_75t_L g12509 ( 
.A(n_12189),
.Y(n_12509)
);

INVx3_ASAP7_75t_L g12510 ( 
.A(n_12305),
.Y(n_12510)
);

NAND2xp5_ASAP7_75t_L g12511 ( 
.A(n_12307),
.B(n_8978),
.Y(n_12511)
);

NAND5xp2_ASAP7_75t_L g12512 ( 
.A(n_12132),
.B(n_12308),
.C(n_12162),
.D(n_12094),
.E(n_12085),
.Y(n_12512)
);

AND2x4_ASAP7_75t_L g12513 ( 
.A(n_12312),
.B(n_8978),
.Y(n_12513)
);

OR2x2_ASAP7_75t_L g12514 ( 
.A(n_12225),
.B(n_8982),
.Y(n_12514)
);

NOR2xp67_ASAP7_75t_L g12515 ( 
.A(n_12005),
.B(n_12079),
.Y(n_12515)
);

AND2x2_ASAP7_75t_L g12516 ( 
.A(n_12222),
.B(n_7066),
.Y(n_12516)
);

AND2x2_ASAP7_75t_SL g12517 ( 
.A(n_12295),
.B(n_6263),
.Y(n_12517)
);

NOR2xp33_ASAP7_75t_L g12518 ( 
.A(n_12160),
.B(n_8995),
.Y(n_12518)
);

NAND2xp5_ASAP7_75t_L g12519 ( 
.A(n_12124),
.B(n_8995),
.Y(n_12519)
);

AND2x2_ASAP7_75t_L g12520 ( 
.A(n_12285),
.B(n_7066),
.Y(n_12520)
);

OR2x2_ASAP7_75t_L g12521 ( 
.A(n_11998),
.B(n_8999),
.Y(n_12521)
);

AND2x2_ASAP7_75t_L g12522 ( 
.A(n_12285),
.B(n_7111),
.Y(n_12522)
);

INVx2_ASAP7_75t_SL g12523 ( 
.A(n_12126),
.Y(n_12523)
);

INVx1_ASAP7_75t_L g12524 ( 
.A(n_12111),
.Y(n_12524)
);

AND2x2_ASAP7_75t_L g12525 ( 
.A(n_12059),
.B(n_7111),
.Y(n_12525)
);

NOR2x1p5_ASAP7_75t_L g12526 ( 
.A(n_11980),
.B(n_6679),
.Y(n_12526)
);

AND2x4_ASAP7_75t_L g12527 ( 
.A(n_12305),
.B(n_12274),
.Y(n_12527)
);

INVx1_ASAP7_75t_L g12528 ( 
.A(n_12152),
.Y(n_12528)
);

INVx1_ASAP7_75t_L g12529 ( 
.A(n_12300),
.Y(n_12529)
);

INVx1_ASAP7_75t_L g12530 ( 
.A(n_12157),
.Y(n_12530)
);

AND2x2_ASAP7_75t_L g12531 ( 
.A(n_12270),
.B(n_7111),
.Y(n_12531)
);

AND2x2_ASAP7_75t_L g12532 ( 
.A(n_12231),
.B(n_7150),
.Y(n_12532)
);

INVx2_ASAP7_75t_SL g12533 ( 
.A(n_12221),
.Y(n_12533)
);

AND2x2_ASAP7_75t_L g12534 ( 
.A(n_11994),
.B(n_12036),
.Y(n_12534)
);

NOR2x1p5_ASAP7_75t_L g12535 ( 
.A(n_11964),
.B(n_6679),
.Y(n_12535)
);

NAND2xp5_ASAP7_75t_L g12536 ( 
.A(n_12281),
.B(n_8999),
.Y(n_12536)
);

INVx1_ASAP7_75t_L g12537 ( 
.A(n_12233),
.Y(n_12537)
);

AND2x2_ASAP7_75t_L g12538 ( 
.A(n_12316),
.B(n_7150),
.Y(n_12538)
);

BUFx2_ASAP7_75t_L g12539 ( 
.A(n_12179),
.Y(n_12539)
);

AND2x4_ASAP7_75t_SL g12540 ( 
.A(n_12018),
.B(n_6984),
.Y(n_12540)
);

INVx1_ASAP7_75t_L g12541 ( 
.A(n_12237),
.Y(n_12541)
);

BUFx2_ASAP7_75t_L g12542 ( 
.A(n_11990),
.Y(n_12542)
);

NOR2xp33_ASAP7_75t_L g12543 ( 
.A(n_12044),
.B(n_9001),
.Y(n_12543)
);

INVx1_ASAP7_75t_L g12544 ( 
.A(n_12013),
.Y(n_12544)
);

NAND2xp5_ASAP7_75t_L g12545 ( 
.A(n_12284),
.B(n_9001),
.Y(n_12545)
);

OR2x2_ASAP7_75t_L g12546 ( 
.A(n_12127),
.B(n_9005),
.Y(n_12546)
);

AND2x2_ASAP7_75t_L g12547 ( 
.A(n_12317),
.B(n_7150),
.Y(n_12547)
);

INVx1_ASAP7_75t_L g12548 ( 
.A(n_12129),
.Y(n_12548)
);

OR2x2_ASAP7_75t_L g12549 ( 
.A(n_12134),
.B(n_9005),
.Y(n_12549)
);

AND2x2_ASAP7_75t_L g12550 ( 
.A(n_12104),
.B(n_12167),
.Y(n_12550)
);

OAI21xp33_ASAP7_75t_L g12551 ( 
.A1(n_12146),
.A2(n_9024),
.B(n_9019),
.Y(n_12551)
);

NOR3xp33_ASAP7_75t_L g12552 ( 
.A(n_12163),
.B(n_9645),
.C(n_9591),
.Y(n_12552)
);

INVx2_ASAP7_75t_L g12553 ( 
.A(n_12151),
.Y(n_12553)
);

OAI31xp33_ASAP7_75t_SL g12554 ( 
.A1(n_12227),
.A2(n_9007),
.A3(n_9009),
.B(n_8968),
.Y(n_12554)
);

OR2x2_ASAP7_75t_L g12555 ( 
.A(n_12072),
.B(n_12228),
.Y(n_12555)
);

AND2x2_ASAP7_75t_L g12556 ( 
.A(n_12118),
.B(n_8253),
.Y(n_12556)
);

HB1xp67_ASAP7_75t_L g12557 ( 
.A(n_12083),
.Y(n_12557)
);

NAND2xp5_ASAP7_75t_L g12558 ( 
.A(n_12289),
.B(n_9019),
.Y(n_12558)
);

INVx1_ASAP7_75t_L g12559 ( 
.A(n_12320),
.Y(n_12559)
);

INVx1_ASAP7_75t_L g12560 ( 
.A(n_12288),
.Y(n_12560)
);

INVx1_ASAP7_75t_L g12561 ( 
.A(n_12313),
.Y(n_12561)
);

INVx2_ASAP7_75t_L g12562 ( 
.A(n_12241),
.Y(n_12562)
);

AND2x2_ASAP7_75t_L g12563 ( 
.A(n_12207),
.B(n_8253),
.Y(n_12563)
);

AND2x2_ASAP7_75t_L g12564 ( 
.A(n_12218),
.B(n_8253),
.Y(n_12564)
);

OR2x2_ASAP7_75t_L g12565 ( 
.A(n_12238),
.B(n_9024),
.Y(n_12565)
);

INVx1_ASAP7_75t_L g12566 ( 
.A(n_12081),
.Y(n_12566)
);

AND2x2_ASAP7_75t_L g12567 ( 
.A(n_12230),
.B(n_8253),
.Y(n_12567)
);

INVx1_ASAP7_75t_L g12568 ( 
.A(n_12224),
.Y(n_12568)
);

INVx2_ASAP7_75t_L g12569 ( 
.A(n_12109),
.Y(n_12569)
);

NAND2x1_ASAP7_75t_L g12570 ( 
.A(n_12179),
.B(n_6679),
.Y(n_12570)
);

INVx1_ASAP7_75t_L g12571 ( 
.A(n_12245),
.Y(n_12571)
);

AND2x2_ASAP7_75t_L g12572 ( 
.A(n_12154),
.B(n_8849),
.Y(n_12572)
);

AND2x2_ASAP7_75t_L g12573 ( 
.A(n_12100),
.B(n_8849),
.Y(n_12573)
);

NOR2xp33_ASAP7_75t_L g12574 ( 
.A(n_12105),
.B(n_7697),
.Y(n_12574)
);

NAND2xp5_ASAP7_75t_L g12575 ( 
.A(n_12232),
.B(n_9016),
.Y(n_12575)
);

INVx1_ASAP7_75t_L g12576 ( 
.A(n_12246),
.Y(n_12576)
);

AND2x2_ASAP7_75t_L g12577 ( 
.A(n_12106),
.B(n_8874),
.Y(n_12577)
);

INVx1_ASAP7_75t_L g12578 ( 
.A(n_11984),
.Y(n_12578)
);

INVx1_ASAP7_75t_L g12579 ( 
.A(n_12290),
.Y(n_12579)
);

AND2x4_ASAP7_75t_L g12580 ( 
.A(n_12297),
.B(n_7373),
.Y(n_12580)
);

OR2x2_ASAP7_75t_L g12581 ( 
.A(n_12098),
.B(n_7982),
.Y(n_12581)
);

OR2x2_ASAP7_75t_L g12582 ( 
.A(n_12101),
.B(n_7982),
.Y(n_12582)
);

INVx2_ASAP7_75t_L g12583 ( 
.A(n_12119),
.Y(n_12583)
);

INVx1_ASAP7_75t_SL g12584 ( 
.A(n_12243),
.Y(n_12584)
);

INVx1_ASAP7_75t_SL g12585 ( 
.A(n_12247),
.Y(n_12585)
);

AND2x2_ASAP7_75t_L g12586 ( 
.A(n_12112),
.B(n_8904),
.Y(n_12586)
);

HB1xp67_ASAP7_75t_L g12587 ( 
.A(n_12309),
.Y(n_12587)
);

AND2x2_ASAP7_75t_L g12588 ( 
.A(n_12123),
.B(n_8904),
.Y(n_12588)
);

INVx3_ASAP7_75t_SL g12589 ( 
.A(n_11992),
.Y(n_12589)
);

INVx1_ASAP7_75t_L g12590 ( 
.A(n_12136),
.Y(n_12590)
);

INVx1_ASAP7_75t_L g12591 ( 
.A(n_12141),
.Y(n_12591)
);

INVx1_ASAP7_75t_L g12592 ( 
.A(n_12318),
.Y(n_12592)
);

INVxp67_ASAP7_75t_L g12593 ( 
.A(n_12296),
.Y(n_12593)
);

NAND2xp5_ASAP7_75t_L g12594 ( 
.A(n_12153),
.B(n_9016),
.Y(n_12594)
);

NOR2xp33_ASAP7_75t_SL g12595 ( 
.A(n_11958),
.B(n_7697),
.Y(n_12595)
);

AOI22xp33_ASAP7_75t_L g12596 ( 
.A1(n_12097),
.A2(n_9012),
.B1(n_9661),
.B2(n_9660),
.Y(n_12596)
);

NAND2xp5_ASAP7_75t_L g12597 ( 
.A(n_12194),
.B(n_9016),
.Y(n_12597)
);

OR2x2_ASAP7_75t_L g12598 ( 
.A(n_12159),
.B(n_7992),
.Y(n_12598)
);

NAND2xp5_ASAP7_75t_L g12599 ( 
.A(n_12194),
.B(n_9016),
.Y(n_12599)
);

AND2x2_ASAP7_75t_L g12600 ( 
.A(n_12249),
.B(n_7992),
.Y(n_12600)
);

INVx4_ASAP7_75t_L g12601 ( 
.A(n_12114),
.Y(n_12601)
);

AND2x2_ASAP7_75t_L g12602 ( 
.A(n_12170),
.B(n_7995),
.Y(n_12602)
);

OR2x2_ASAP7_75t_L g12603 ( 
.A(n_12182),
.B(n_7995),
.Y(n_12603)
);

OR2x2_ASAP7_75t_L g12604 ( 
.A(n_12183),
.B(n_12184),
.Y(n_12604)
);

AND2x2_ASAP7_75t_L g12605 ( 
.A(n_12139),
.B(n_12282),
.Y(n_12605)
);

INVx1_ASAP7_75t_L g12606 ( 
.A(n_12164),
.Y(n_12606)
);

INVx1_ASAP7_75t_L g12607 ( 
.A(n_12263),
.Y(n_12607)
);

AND4x1_ASAP7_75t_L g12608 ( 
.A(n_12186),
.B(n_7395),
.C(n_7139),
.D(n_7119),
.Y(n_12608)
);

OR2x2_ASAP7_75t_L g12609 ( 
.A(n_12096),
.B(n_8008),
.Y(n_12609)
);

INVx2_ASAP7_75t_L g12610 ( 
.A(n_12211),
.Y(n_12610)
);

AND2x2_ASAP7_75t_L g12611 ( 
.A(n_12212),
.B(n_8008),
.Y(n_12611)
);

NAND2xp5_ASAP7_75t_L g12612 ( 
.A(n_12251),
.B(n_9016),
.Y(n_12612)
);

AND2x4_ASAP7_75t_L g12613 ( 
.A(n_12277),
.B(n_7373),
.Y(n_12613)
);

AND2x4_ASAP7_75t_L g12614 ( 
.A(n_12116),
.B(n_8968),
.Y(n_12614)
);

INVx3_ASAP7_75t_L g12615 ( 
.A(n_12251),
.Y(n_12615)
);

OAI221xp5_ASAP7_75t_L g12616 ( 
.A1(n_12177),
.A2(n_8850),
.B1(n_8809),
.B2(n_9670),
.C(n_9667),
.Y(n_12616)
);

AND2x2_ASAP7_75t_L g12617 ( 
.A(n_12168),
.B(n_12169),
.Y(n_12617)
);

INVx1_ASAP7_75t_L g12618 ( 
.A(n_12306),
.Y(n_12618)
);

INVx1_ASAP7_75t_L g12619 ( 
.A(n_12192),
.Y(n_12619)
);

INVx3_ASAP7_75t_L g12620 ( 
.A(n_12264),
.Y(n_12620)
);

AND2x2_ASAP7_75t_L g12621 ( 
.A(n_12201),
.B(n_8011),
.Y(n_12621)
);

INVx1_ASAP7_75t_L g12622 ( 
.A(n_12310),
.Y(n_12622)
);

AOI221xp5_ASAP7_75t_L g12623 ( 
.A1(n_11993),
.A2(n_9691),
.B1(n_9704),
.B2(n_9678),
.C(n_9677),
.Y(n_12623)
);

AOI22xp33_ASAP7_75t_L g12624 ( 
.A1(n_11997),
.A2(n_9012),
.B1(n_9719),
.B2(n_9713),
.Y(n_12624)
);

INVx1_ASAP7_75t_L g12625 ( 
.A(n_12130),
.Y(n_12625)
);

INVx1_ASAP7_75t_L g12626 ( 
.A(n_12272),
.Y(n_12626)
);

AND2x4_ASAP7_75t_L g12627 ( 
.A(n_12117),
.B(n_9007),
.Y(n_12627)
);

OR2x2_ASAP7_75t_L g12628 ( 
.A(n_12205),
.B(n_8011),
.Y(n_12628)
);

NAND2xp5_ASAP7_75t_SL g12629 ( 
.A(n_12198),
.B(n_5673),
.Y(n_12629)
);

NOR3xp33_ASAP7_75t_SL g12630 ( 
.A(n_12138),
.B(n_7265),
.C(n_7286),
.Y(n_12630)
);

NAND3x1_ASAP7_75t_L g12631 ( 
.A(n_12214),
.B(n_6759),
.C(n_6679),
.Y(n_12631)
);

OR2x2_ASAP7_75t_L g12632 ( 
.A(n_12206),
.B(n_12042),
.Y(n_12632)
);

NAND2xp5_ASAP7_75t_L g12633 ( 
.A(n_12314),
.B(n_9029),
.Y(n_12633)
);

AND2x2_ASAP7_75t_L g12634 ( 
.A(n_12202),
.B(n_8018),
.Y(n_12634)
);

AND2x2_ASAP7_75t_L g12635 ( 
.A(n_12187),
.B(n_8018),
.Y(n_12635)
);

INVx1_ASAP7_75t_SL g12636 ( 
.A(n_12176),
.Y(n_12636)
);

INVx2_ASAP7_75t_L g12637 ( 
.A(n_12145),
.Y(n_12637)
);

AND2x2_ASAP7_75t_L g12638 ( 
.A(n_12191),
.B(n_8023),
.Y(n_12638)
);

AND3x2_ASAP7_75t_L g12639 ( 
.A(n_12048),
.B(n_6086),
.C(n_6062),
.Y(n_12639)
);

AND2x2_ASAP7_75t_L g12640 ( 
.A(n_12204),
.B(n_8023),
.Y(n_12640)
);

NAND2xp5_ASAP7_75t_L g12641 ( 
.A(n_12319),
.B(n_9029),
.Y(n_12641)
);

OR2x2_ASAP7_75t_L g12642 ( 
.A(n_12049),
.B(n_8027),
.Y(n_12642)
);

HB1xp67_ASAP7_75t_L g12643 ( 
.A(n_12107),
.Y(n_12643)
);

INVx2_ASAP7_75t_L g12644 ( 
.A(n_12273),
.Y(n_12644)
);

NAND2xp5_ASAP7_75t_L g12645 ( 
.A(n_12323),
.B(n_9029),
.Y(n_12645)
);

INVx1_ASAP7_75t_L g12646 ( 
.A(n_12294),
.Y(n_12646)
);

INVx6_ASAP7_75t_L g12647 ( 
.A(n_12248),
.Y(n_12647)
);

NOR2xp33_ASAP7_75t_SL g12648 ( 
.A(n_12125),
.B(n_12250),
.Y(n_12648)
);

AOI31xp33_ASAP7_75t_L g12649 ( 
.A1(n_12266),
.A2(n_7286),
.A3(n_7297),
.B(n_7265),
.Y(n_12649)
);

INVx2_ASAP7_75t_L g12650 ( 
.A(n_12273),
.Y(n_12650)
);

INVx1_ASAP7_75t_L g12651 ( 
.A(n_12287),
.Y(n_12651)
);

AND2x2_ASAP7_75t_L g12652 ( 
.A(n_12217),
.B(n_8027),
.Y(n_12652)
);

AND2x2_ASAP7_75t_L g12653 ( 
.A(n_12256),
.B(n_8033),
.Y(n_12653)
);

BUFx2_ASAP7_75t_L g12654 ( 
.A(n_12240),
.Y(n_12654)
);

INVx1_ASAP7_75t_L g12655 ( 
.A(n_12301),
.Y(n_12655)
);

NAND2xp5_ASAP7_75t_L g12656 ( 
.A(n_12050),
.B(n_9029),
.Y(n_12656)
);

AND2x2_ASAP7_75t_L g12657 ( 
.A(n_12235),
.B(n_8033),
.Y(n_12657)
);

INVx1_ASAP7_75t_SL g12658 ( 
.A(n_12215),
.Y(n_12658)
);

AND2x2_ASAP7_75t_L g12659 ( 
.A(n_12226),
.B(n_8035),
.Y(n_12659)
);

OR2x2_ASAP7_75t_L g12660 ( 
.A(n_12051),
.B(n_8035),
.Y(n_12660)
);

AND2x4_ASAP7_75t_L g12661 ( 
.A(n_12052),
.B(n_9009),
.Y(n_12661)
);

INVx6_ASAP7_75t_L g12662 ( 
.A(n_12311),
.Y(n_12662)
);

INVx1_ASAP7_75t_L g12663 ( 
.A(n_12302),
.Y(n_12663)
);

AND2x2_ASAP7_75t_L g12664 ( 
.A(n_12265),
.B(n_8047),
.Y(n_12664)
);

INVx2_ASAP7_75t_L g12665 ( 
.A(n_12278),
.Y(n_12665)
);

INVx1_ASAP7_75t_L g12666 ( 
.A(n_12322),
.Y(n_12666)
);

NAND2xp5_ASAP7_75t_L g12667 ( 
.A(n_12054),
.B(n_9029),
.Y(n_12667)
);

NAND4xp25_ASAP7_75t_L g12668 ( 
.A(n_12150),
.B(n_7297),
.C(n_7401),
.D(n_7331),
.Y(n_12668)
);

AND2x4_ASAP7_75t_SL g12669 ( 
.A(n_12267),
.B(n_6984),
.Y(n_12669)
);

AOI22xp5_ASAP7_75t_L g12670 ( 
.A1(n_12364),
.A2(n_12260),
.B1(n_12254),
.B2(n_12259),
.Y(n_12670)
);

AND2x2_ASAP7_75t_L g12671 ( 
.A(n_12390),
.B(n_12193),
.Y(n_12671)
);

INVx1_ASAP7_75t_L g12672 ( 
.A(n_12451),
.Y(n_12672)
);

INVx1_ASAP7_75t_L g12673 ( 
.A(n_12510),
.Y(n_12673)
);

INVx2_ASAP7_75t_SL g12674 ( 
.A(n_12379),
.Y(n_12674)
);

INVx1_ASAP7_75t_L g12675 ( 
.A(n_12328),
.Y(n_12675)
);

INVx1_ASAP7_75t_L g12676 ( 
.A(n_12527),
.Y(n_12676)
);

OR2x2_ASAP7_75t_L g12677 ( 
.A(n_12366),
.B(n_12195),
.Y(n_12677)
);

INVx3_ASAP7_75t_L g12678 ( 
.A(n_12379),
.Y(n_12678)
);

AND2x2_ASAP7_75t_L g12679 ( 
.A(n_12324),
.B(n_12199),
.Y(n_12679)
);

INVx1_ASAP7_75t_SL g12680 ( 
.A(n_12386),
.Y(n_12680)
);

NAND2xp5_ASAP7_75t_L g12681 ( 
.A(n_12402),
.B(n_12200),
.Y(n_12681)
);

NAND2xp5_ASAP7_75t_L g12682 ( 
.A(n_12455),
.B(n_12121),
.Y(n_12682)
);

OAI322xp33_ASAP7_75t_L g12683 ( 
.A1(n_12327),
.A2(n_12172),
.A3(n_12203),
.B1(n_12268),
.B2(n_12275),
.C1(n_12276),
.C2(n_12236),
.Y(n_12683)
);

AOI22xp5_ASAP7_75t_L g12684 ( 
.A1(n_12348),
.A2(n_12262),
.B1(n_12286),
.B2(n_12283),
.Y(n_12684)
);

NAND2xp5_ASAP7_75t_L g12685 ( 
.A(n_12455),
.B(n_12135),
.Y(n_12685)
);

INVx1_ASAP7_75t_L g12686 ( 
.A(n_12527),
.Y(n_12686)
);

INVx1_ASAP7_75t_SL g12687 ( 
.A(n_12377),
.Y(n_12687)
);

INVx1_ASAP7_75t_L g12688 ( 
.A(n_12587),
.Y(n_12688)
);

INVxp67_ASAP7_75t_L g12689 ( 
.A(n_12356),
.Y(n_12689)
);

INVx1_ASAP7_75t_L g12690 ( 
.A(n_12371),
.Y(n_12690)
);

OAI22xp5_ASAP7_75t_L g12691 ( 
.A1(n_12340),
.A2(n_12185),
.B1(n_12213),
.B2(n_12279),
.Y(n_12691)
);

AND2x2_ASAP7_75t_L g12692 ( 
.A(n_12352),
.B(n_12280),
.Y(n_12692)
);

INVx1_ASAP7_75t_L g12693 ( 
.A(n_12441),
.Y(n_12693)
);

NAND2xp5_ASAP7_75t_L g12694 ( 
.A(n_12382),
.B(n_12178),
.Y(n_12694)
);

INVx1_ASAP7_75t_L g12695 ( 
.A(n_12441),
.Y(n_12695)
);

INVx1_ASAP7_75t_L g12696 ( 
.A(n_12374),
.Y(n_12696)
);

AOI33xp33_ASAP7_75t_L g12697 ( 
.A1(n_12380),
.A2(n_12197),
.A3(n_12208),
.B1(n_12196),
.B2(n_5850),
.B3(n_5721),
.Y(n_12697)
);

INVx1_ASAP7_75t_L g12698 ( 
.A(n_12495),
.Y(n_12698)
);

AOI33xp33_ASAP7_75t_L g12699 ( 
.A1(n_12385),
.A2(n_5850),
.A3(n_5721),
.B1(n_5906),
.B2(n_5757),
.B3(n_5680),
.Y(n_12699)
);

AOI22xp5_ASAP7_75t_L g12700 ( 
.A1(n_12399),
.A2(n_9110),
.B1(n_9105),
.B2(n_8850),
.Y(n_12700)
);

INVx1_ASAP7_75t_L g12701 ( 
.A(n_12372),
.Y(n_12701)
);

INVx1_ASAP7_75t_L g12702 ( 
.A(n_12412),
.Y(n_12702)
);

NAND2xp5_ASAP7_75t_L g12703 ( 
.A(n_12394),
.B(n_8047),
.Y(n_12703)
);

NAND2xp5_ASAP7_75t_R g12704 ( 
.A(n_12354),
.B(n_8259),
.Y(n_12704)
);

INVx1_ASAP7_75t_L g12705 ( 
.A(n_12393),
.Y(n_12705)
);

A2O1A1Ixp33_ASAP7_75t_L g12706 ( 
.A1(n_12554),
.A2(n_8949),
.B(n_8956),
.C(n_8943),
.Y(n_12706)
);

A2O1A1Ixp33_ASAP7_75t_L g12707 ( 
.A1(n_12422),
.A2(n_8956),
.B(n_8639),
.C(n_8641),
.Y(n_12707)
);

OR2x2_ASAP7_75t_L g12708 ( 
.A(n_12429),
.B(n_8053),
.Y(n_12708)
);

INVx1_ASAP7_75t_L g12709 ( 
.A(n_12387),
.Y(n_12709)
);

AND2x2_ASAP7_75t_L g12710 ( 
.A(n_12346),
.B(n_6679),
.Y(n_12710)
);

INVxp67_ASAP7_75t_L g12711 ( 
.A(n_12512),
.Y(n_12711)
);

INVx1_ASAP7_75t_L g12712 ( 
.A(n_12397),
.Y(n_12712)
);

AOI22xp5_ASAP7_75t_L g12713 ( 
.A1(n_12409),
.A2(n_9110),
.B1(n_9105),
.B2(n_8850),
.Y(n_12713)
);

AOI211xp5_ASAP7_75t_L g12714 ( 
.A1(n_12407),
.A2(n_6647),
.B(n_7401),
.C(n_7331),
.Y(n_12714)
);

OR2x2_ASAP7_75t_L g12715 ( 
.A(n_12337),
.B(n_8053),
.Y(n_12715)
);

OAI22xp5_ASAP7_75t_L g12716 ( 
.A1(n_12389),
.A2(n_9132),
.B1(n_9138),
.B2(n_9131),
.Y(n_12716)
);

OAI32xp33_ASAP7_75t_L g12717 ( 
.A1(n_12439),
.A2(n_8641),
.A3(n_8652),
.B1(n_8639),
.B2(n_8636),
.Y(n_12717)
);

INVx1_ASAP7_75t_L g12718 ( 
.A(n_12403),
.Y(n_12718)
);

INVx2_ASAP7_75t_L g12719 ( 
.A(n_12360),
.Y(n_12719)
);

OAI31xp33_ASAP7_75t_SL g12720 ( 
.A1(n_12447),
.A2(n_7833),
.A3(n_5757),
.B(n_5906),
.Y(n_12720)
);

INVx1_ASAP7_75t_L g12721 ( 
.A(n_12408),
.Y(n_12721)
);

INVx1_ASAP7_75t_L g12722 ( 
.A(n_12405),
.Y(n_12722)
);

INVx2_ASAP7_75t_SL g12723 ( 
.A(n_12367),
.Y(n_12723)
);

INVx1_ASAP7_75t_L g12724 ( 
.A(n_12405),
.Y(n_12724)
);

INVx1_ASAP7_75t_L g12725 ( 
.A(n_12414),
.Y(n_12725)
);

NAND2xp5_ASAP7_75t_L g12726 ( 
.A(n_12367),
.B(n_8055),
.Y(n_12726)
);

AOI22xp5_ASAP7_75t_L g12727 ( 
.A1(n_12375),
.A2(n_12616),
.B1(n_12351),
.B2(n_12467),
.Y(n_12727)
);

AND2x2_ASAP7_75t_L g12728 ( 
.A(n_12326),
.B(n_12369),
.Y(n_12728)
);

AND2x2_ASAP7_75t_L g12729 ( 
.A(n_12365),
.B(n_6759),
.Y(n_12729)
);

INVx3_ASAP7_75t_L g12730 ( 
.A(n_12416),
.Y(n_12730)
);

OAI322xp33_ASAP7_75t_L g12731 ( 
.A1(n_12648),
.A2(n_8657),
.A3(n_8636),
.B1(n_8658),
.B2(n_8661),
.C1(n_8659),
.C2(n_8652),
.Y(n_12731)
);

INVx2_ASAP7_75t_L g12732 ( 
.A(n_12378),
.Y(n_12732)
);

AOI22xp5_ASAP7_75t_L g12733 ( 
.A1(n_12644),
.A2(n_9105),
.B1(n_9110),
.B2(n_8809),
.Y(n_12733)
);

OA222x2_ASAP7_75t_L g12734 ( 
.A1(n_12383),
.A2(n_6759),
.B1(n_6904),
.B2(n_6965),
.C1(n_6906),
.C2(n_6812),
.Y(n_12734)
);

INVx1_ASAP7_75t_SL g12735 ( 
.A(n_12347),
.Y(n_12735)
);

OAI22xp5_ASAP7_75t_L g12736 ( 
.A1(n_12423),
.A2(n_9132),
.B1(n_9138),
.B2(n_9131),
.Y(n_12736)
);

NOR2xp33_ASAP7_75t_L g12737 ( 
.A(n_12358),
.B(n_7697),
.Y(n_12737)
);

OAI21xp33_ASAP7_75t_SL g12738 ( 
.A1(n_12649),
.A2(n_12338),
.B(n_12445),
.Y(n_12738)
);

INVx1_ASAP7_75t_L g12739 ( 
.A(n_12542),
.Y(n_12739)
);

NAND2xp5_ASAP7_75t_L g12740 ( 
.A(n_12416),
.B(n_8055),
.Y(n_12740)
);

INVx1_ASAP7_75t_L g12741 ( 
.A(n_12542),
.Y(n_12741)
);

INVx1_ASAP7_75t_L g12742 ( 
.A(n_12413),
.Y(n_12742)
);

OR2x2_ASAP7_75t_L g12743 ( 
.A(n_12381),
.B(n_8056),
.Y(n_12743)
);

INVx2_ASAP7_75t_SL g12744 ( 
.A(n_12647),
.Y(n_12744)
);

NAND2xp5_ASAP7_75t_L g12745 ( 
.A(n_12325),
.B(n_8056),
.Y(n_12745)
);

NAND2x1_ASAP7_75t_L g12746 ( 
.A(n_12662),
.B(n_6759),
.Y(n_12746)
);

INVx1_ASAP7_75t_L g12747 ( 
.A(n_12426),
.Y(n_12747)
);

OAI22xp33_ASAP7_75t_L g12748 ( 
.A1(n_12430),
.A2(n_9140),
.B1(n_9150),
.B2(n_9149),
.Y(n_12748)
);

INVx1_ASAP7_75t_L g12749 ( 
.A(n_12465),
.Y(n_12749)
);

AND2x4_ASAP7_75t_L g12750 ( 
.A(n_12388),
.B(n_9140),
.Y(n_12750)
);

INVx1_ASAP7_75t_L g12751 ( 
.A(n_12506),
.Y(n_12751)
);

OR2x2_ASAP7_75t_L g12752 ( 
.A(n_12350),
.B(n_8060),
.Y(n_12752)
);

NAND2xp5_ASAP7_75t_L g12753 ( 
.A(n_12391),
.B(n_8067),
.Y(n_12753)
);

OAI33xp33_ASAP7_75t_L g12754 ( 
.A1(n_12329),
.A2(n_8661),
.A3(n_8658),
.B1(n_8672),
.B2(n_8659),
.B3(n_8657),
.Y(n_12754)
);

AOI211xp5_ASAP7_75t_L g12755 ( 
.A1(n_12353),
.A2(n_7175),
.B(n_9150),
.C(n_9149),
.Y(n_12755)
);

INVxp67_ASAP7_75t_L g12756 ( 
.A(n_12539),
.Y(n_12756)
);

INVx1_ASAP7_75t_L g12757 ( 
.A(n_12509),
.Y(n_12757)
);

INVx1_ASAP7_75t_L g12758 ( 
.A(n_12427),
.Y(n_12758)
);

NAND2xp5_ASAP7_75t_L g12759 ( 
.A(n_12341),
.B(n_8067),
.Y(n_12759)
);

INVx2_ASAP7_75t_L g12760 ( 
.A(n_12662),
.Y(n_12760)
);

NAND4xp75_ASAP7_75t_L g12761 ( 
.A(n_12515),
.B(n_8809),
.C(n_8588),
.D(n_6503),
.Y(n_12761)
);

INVx1_ASAP7_75t_L g12762 ( 
.A(n_12431),
.Y(n_12762)
);

INVx1_ASAP7_75t_L g12763 ( 
.A(n_12450),
.Y(n_12763)
);

INVx2_ASAP7_75t_L g12764 ( 
.A(n_12373),
.Y(n_12764)
);

AOI22xp5_ASAP7_75t_L g12765 ( 
.A1(n_12650),
.A2(n_8672),
.B1(n_8693),
.B2(n_9012),
.Y(n_12765)
);

INVx1_ASAP7_75t_L g12766 ( 
.A(n_12480),
.Y(n_12766)
);

OAI21xp5_ASAP7_75t_SL g12767 ( 
.A1(n_12334),
.A2(n_6812),
.B(n_6759),
.Y(n_12767)
);

OR2x2_ASAP7_75t_L g12768 ( 
.A(n_12383),
.B(n_8084),
.Y(n_12768)
);

INVx1_ASAP7_75t_L g12769 ( 
.A(n_12475),
.Y(n_12769)
);

INVx2_ASAP7_75t_L g12770 ( 
.A(n_12520),
.Y(n_12770)
);

INVx1_ASAP7_75t_L g12771 ( 
.A(n_12502),
.Y(n_12771)
);

AOI22xp5_ASAP7_75t_L g12772 ( 
.A1(n_12497),
.A2(n_8693),
.B1(n_9153),
.B2(n_8588),
.Y(n_12772)
);

INVx1_ASAP7_75t_L g12773 ( 
.A(n_12332),
.Y(n_12773)
);

INVx1_ASAP7_75t_L g12774 ( 
.A(n_12336),
.Y(n_12774)
);

NOR4xp25_ASAP7_75t_L g12775 ( 
.A(n_12349),
.B(n_9153),
.C(n_8084),
.D(n_8090),
.Y(n_12775)
);

INVx1_ASAP7_75t_L g12776 ( 
.A(n_12339),
.Y(n_12776)
);

OR2x2_ASAP7_75t_L g12777 ( 
.A(n_12420),
.B(n_8088),
.Y(n_12777)
);

INVx2_ASAP7_75t_SL g12778 ( 
.A(n_12647),
.Y(n_12778)
);

AND2x4_ASAP7_75t_L g12779 ( 
.A(n_12444),
.B(n_12362),
.Y(n_12779)
);

INVxp67_ASAP7_75t_L g12780 ( 
.A(n_12654),
.Y(n_12780)
);

INVx1_ASAP7_75t_L g12781 ( 
.A(n_12345),
.Y(n_12781)
);

INVx2_ASAP7_75t_L g12782 ( 
.A(n_12522),
.Y(n_12782)
);

INVx1_ASAP7_75t_L g12783 ( 
.A(n_12557),
.Y(n_12783)
);

OAI22xp33_ASAP7_75t_L g12784 ( 
.A1(n_12487),
.A2(n_7828),
.B1(n_7697),
.B2(n_8588),
.Y(n_12784)
);

AOI21xp33_ASAP7_75t_SL g12785 ( 
.A1(n_12589),
.A2(n_7828),
.B(n_7605),
.Y(n_12785)
);

INVx1_ASAP7_75t_L g12786 ( 
.A(n_12433),
.Y(n_12786)
);

O2A1O1Ixp5_ASAP7_75t_R g12787 ( 
.A1(n_12392),
.A2(n_7277),
.B(n_6149),
.C(n_7828),
.Y(n_12787)
);

OR2x2_ASAP7_75t_L g12788 ( 
.A(n_12357),
.B(n_8088),
.Y(n_12788)
);

INVx1_ASAP7_75t_L g12789 ( 
.A(n_12344),
.Y(n_12789)
);

INVx2_ASAP7_75t_L g12790 ( 
.A(n_12484),
.Y(n_12790)
);

INVx2_ASAP7_75t_SL g12791 ( 
.A(n_12362),
.Y(n_12791)
);

NAND2xp5_ASAP7_75t_L g12792 ( 
.A(n_12342),
.B(n_8090),
.Y(n_12792)
);

INVx1_ASAP7_75t_L g12793 ( 
.A(n_12330),
.Y(n_12793)
);

BUFx2_ASAP7_75t_L g12794 ( 
.A(n_12404),
.Y(n_12794)
);

INVx2_ASAP7_75t_L g12795 ( 
.A(n_12615),
.Y(n_12795)
);

NAND2xp5_ASAP7_75t_L g12796 ( 
.A(n_12363),
.B(n_8093),
.Y(n_12796)
);

HB1xp67_ASAP7_75t_L g12797 ( 
.A(n_12398),
.Y(n_12797)
);

AND2x2_ASAP7_75t_L g12798 ( 
.A(n_12425),
.B(n_6812),
.Y(n_12798)
);

NAND2xp5_ASAP7_75t_L g12799 ( 
.A(n_12466),
.B(n_8093),
.Y(n_12799)
);

AOI22xp33_ASAP7_75t_SL g12800 ( 
.A1(n_12543),
.A2(n_7828),
.B1(n_7471),
.B2(n_7605),
.Y(n_12800)
);

INVx1_ASAP7_75t_L g12801 ( 
.A(n_12333),
.Y(n_12801)
);

OR2x6_ASAP7_75t_L g12802 ( 
.A(n_12335),
.B(n_7828),
.Y(n_12802)
);

AO22x1_ASAP7_75t_L g12803 ( 
.A1(n_12419),
.A2(n_6812),
.B1(n_6906),
.B2(n_6904),
.Y(n_12803)
);

INVxp67_ASAP7_75t_L g12804 ( 
.A(n_12401),
.Y(n_12804)
);

OR2x2_ASAP7_75t_L g12805 ( 
.A(n_12424),
.B(n_12637),
.Y(n_12805)
);

INVx1_ASAP7_75t_L g12806 ( 
.A(n_12534),
.Y(n_12806)
);

INVx1_ASAP7_75t_SL g12807 ( 
.A(n_12384),
.Y(n_12807)
);

INVx1_ASAP7_75t_L g12808 ( 
.A(n_12434),
.Y(n_12808)
);

INVx1_ASAP7_75t_L g12809 ( 
.A(n_12411),
.Y(n_12809)
);

INVx1_ASAP7_75t_L g12810 ( 
.A(n_12493),
.Y(n_12810)
);

INVx2_ASAP7_75t_L g12811 ( 
.A(n_12526),
.Y(n_12811)
);

AND2x2_ASAP7_75t_L g12812 ( 
.A(n_12605),
.B(n_12617),
.Y(n_12812)
);

NOR3xp33_ASAP7_75t_L g12813 ( 
.A(n_12432),
.B(n_6687),
.C(n_6809),
.Y(n_12813)
);

NAND2xp5_ASAP7_75t_L g12814 ( 
.A(n_12501),
.B(n_8118),
.Y(n_12814)
);

OR2x2_ASAP7_75t_L g12815 ( 
.A(n_12331),
.B(n_8118),
.Y(n_12815)
);

OR2x2_ASAP7_75t_L g12816 ( 
.A(n_12415),
.B(n_8141),
.Y(n_12816)
);

NAND2xp5_ASAP7_75t_L g12817 ( 
.A(n_12544),
.B(n_8141),
.Y(n_12817)
);

INVxp67_ASAP7_75t_SL g12818 ( 
.A(n_12421),
.Y(n_12818)
);

OAI21xp33_ASAP7_75t_L g12819 ( 
.A1(n_12595),
.A2(n_12630),
.B(n_12574),
.Y(n_12819)
);

AOI22xp5_ASAP7_75t_L g12820 ( 
.A1(n_12518),
.A2(n_5680),
.B1(n_6687),
.B2(n_6936),
.Y(n_12820)
);

OR2x2_ASAP7_75t_L g12821 ( 
.A(n_12410),
.B(n_8154),
.Y(n_12821)
);

INVx1_ASAP7_75t_L g12822 ( 
.A(n_12449),
.Y(n_12822)
);

INVx2_ASAP7_75t_SL g12823 ( 
.A(n_12535),
.Y(n_12823)
);

INVx1_ASAP7_75t_L g12824 ( 
.A(n_12555),
.Y(n_12824)
);

INVx1_ASAP7_75t_L g12825 ( 
.A(n_12531),
.Y(n_12825)
);

INVxp67_ASAP7_75t_L g12826 ( 
.A(n_12494),
.Y(n_12826)
);

AND2x2_ASAP7_75t_L g12827 ( 
.A(n_12468),
.B(n_6812),
.Y(n_12827)
);

INVx1_ASAP7_75t_L g12828 ( 
.A(n_12355),
.Y(n_12828)
);

AOI22xp5_ASAP7_75t_L g12829 ( 
.A1(n_12572),
.A2(n_6988),
.B1(n_7020),
.B2(n_6959),
.Y(n_12829)
);

AOI32xp33_ASAP7_75t_L g12830 ( 
.A1(n_12396),
.A2(n_6602),
.A3(n_6604),
.B1(n_6811),
.B2(n_6809),
.Y(n_12830)
);

OAI22xp5_ASAP7_75t_L g12831 ( 
.A1(n_12442),
.A2(n_8158),
.B1(n_8159),
.B2(n_8154),
.Y(n_12831)
);

AND2x4_ASAP7_75t_L g12832 ( 
.A(n_12553),
.B(n_8158),
.Y(n_12832)
);

OR2x6_ASAP7_75t_L g12833 ( 
.A(n_12460),
.B(n_7799),
.Y(n_12833)
);

INVx1_ASAP7_75t_L g12834 ( 
.A(n_12632),
.Y(n_12834)
);

AOI22xp5_ASAP7_75t_L g12835 ( 
.A1(n_12552),
.A2(n_7020),
.B1(n_6959),
.B2(n_6904),
.Y(n_12835)
);

INVx1_ASAP7_75t_L g12836 ( 
.A(n_12435),
.Y(n_12836)
);

INVx1_ASAP7_75t_SL g12837 ( 
.A(n_12584),
.Y(n_12837)
);

INVx2_ASAP7_75t_SL g12838 ( 
.A(n_12540),
.Y(n_12838)
);

XNOR2x2_ASAP7_75t_L g12839 ( 
.A(n_12585),
.B(n_7498),
.Y(n_12839)
);

INVx1_ASAP7_75t_L g12840 ( 
.A(n_12359),
.Y(n_12840)
);

AND3x2_ASAP7_75t_L g12841 ( 
.A(n_12368),
.B(n_8161),
.C(n_8159),
.Y(n_12841)
);

OAI32xp33_ASAP7_75t_L g12842 ( 
.A1(n_12436),
.A2(n_6965),
.A3(n_6980),
.B1(n_6906),
.B2(n_6904),
.Y(n_12842)
);

HB1xp67_ASAP7_75t_L g12843 ( 
.A(n_12370),
.Y(n_12843)
);

INVx1_ASAP7_75t_L g12844 ( 
.A(n_12513),
.Y(n_12844)
);

OAI22xp33_ASAP7_75t_L g12845 ( 
.A1(n_12519),
.A2(n_7471),
.B1(n_7605),
.B2(n_7450),
.Y(n_12845)
);

INVx1_ASAP7_75t_L g12846 ( 
.A(n_12513),
.Y(n_12846)
);

OR2x2_ASAP7_75t_SL g12847 ( 
.A(n_12457),
.B(n_7033),
.Y(n_12847)
);

AO22x1_ASAP7_75t_L g12848 ( 
.A1(n_12498),
.A2(n_6906),
.B1(n_6965),
.B2(n_6904),
.Y(n_12848)
);

NAND2xp5_ASAP7_75t_L g12849 ( 
.A(n_12606),
.B(n_8161),
.Y(n_12849)
);

NAND2xp5_ASAP7_75t_L g12850 ( 
.A(n_12625),
.B(n_8166),
.Y(n_12850)
);

AND2x2_ASAP7_75t_L g12851 ( 
.A(n_12525),
.B(n_6906),
.Y(n_12851)
);

AOI22xp5_ASAP7_75t_L g12852 ( 
.A1(n_12503),
.A2(n_7020),
.B1(n_7084),
.B2(n_6965),
.Y(n_12852)
);

INVx2_ASAP7_75t_L g12853 ( 
.A(n_12478),
.Y(n_12853)
);

INVx3_ASAP7_75t_L g12854 ( 
.A(n_12601),
.Y(n_12854)
);

INVx2_ASAP7_75t_L g12855 ( 
.A(n_12604),
.Y(n_12855)
);

AND2x4_ASAP7_75t_L g12856 ( 
.A(n_12464),
.B(n_12395),
.Y(n_12856)
);

OAI21xp5_ASAP7_75t_L g12857 ( 
.A1(n_12469),
.A2(n_7514),
.B(n_7498),
.Y(n_12857)
);

NAND2xp5_ASAP7_75t_L g12858 ( 
.A(n_12579),
.B(n_12462),
.Y(n_12858)
);

OAI22xp33_ASAP7_75t_L g12859 ( 
.A1(n_12482),
.A2(n_7471),
.B1(n_7612),
.B2(n_7450),
.Y(n_12859)
);

NAND2xp5_ASAP7_75t_L g12860 ( 
.A(n_12524),
.B(n_8166),
.Y(n_12860)
);

INVx2_ASAP7_75t_L g12861 ( 
.A(n_12514),
.Y(n_12861)
);

INVx1_ASAP7_75t_L g12862 ( 
.A(n_12471),
.Y(n_12862)
);

INVx1_ASAP7_75t_L g12863 ( 
.A(n_12418),
.Y(n_12863)
);

OAI22xp33_ASAP7_75t_SL g12864 ( 
.A1(n_12461),
.A2(n_12496),
.B1(n_12529),
.B2(n_12594),
.Y(n_12864)
);

INVx1_ASAP7_75t_L g12865 ( 
.A(n_12565),
.Y(n_12865)
);

INVx1_ASAP7_75t_L g12866 ( 
.A(n_12406),
.Y(n_12866)
);

INVx1_ASAP7_75t_L g12867 ( 
.A(n_12428),
.Y(n_12867)
);

AOI22xp5_ASAP7_75t_L g12868 ( 
.A1(n_12573),
.A2(n_7084),
.B1(n_7194),
.B2(n_6965),
.Y(n_12868)
);

OAI32xp33_ASAP7_75t_L g12869 ( 
.A1(n_12619),
.A2(n_7194),
.A3(n_7219),
.B1(n_7084),
.B2(n_6980),
.Y(n_12869)
);

INVx1_ASAP7_75t_L g12870 ( 
.A(n_12343),
.Y(n_12870)
);

INVx1_ASAP7_75t_L g12871 ( 
.A(n_12500),
.Y(n_12871)
);

OAI32xp33_ASAP7_75t_L g12872 ( 
.A1(n_12443),
.A2(n_7194),
.A3(n_7219),
.B1(n_7084),
.B2(n_6980),
.Y(n_12872)
);

INVx2_ASAP7_75t_L g12873 ( 
.A(n_12570),
.Y(n_12873)
);

INVx1_ASAP7_75t_L g12874 ( 
.A(n_12528),
.Y(n_12874)
);

INVx1_ASAP7_75t_L g12875 ( 
.A(n_12530),
.Y(n_12875)
);

INVxp67_ASAP7_75t_L g12876 ( 
.A(n_12550),
.Y(n_12876)
);

INVx1_ASAP7_75t_L g12877 ( 
.A(n_12521),
.Y(n_12877)
);

INVx2_ASAP7_75t_L g12878 ( 
.A(n_12485),
.Y(n_12878)
);

NAND4xp25_ASAP7_75t_L g12879 ( 
.A(n_12459),
.B(n_6529),
.C(n_7139),
.D(n_7119),
.Y(n_12879)
);

NAND2xp5_ASAP7_75t_L g12880 ( 
.A(n_12666),
.B(n_12590),
.Y(n_12880)
);

AOI22xp5_ASAP7_75t_L g12881 ( 
.A1(n_12577),
.A2(n_7084),
.B1(n_7194),
.B2(n_6980),
.Y(n_12881)
);

INVx2_ASAP7_75t_L g12882 ( 
.A(n_12639),
.Y(n_12882)
);

NOR2xp33_ASAP7_75t_L g12883 ( 
.A(n_12551),
.B(n_8335),
.Y(n_12883)
);

NAND2xp5_ASAP7_75t_L g12884 ( 
.A(n_12591),
.B(n_8169),
.Y(n_12884)
);

OAI32xp33_ASAP7_75t_L g12885 ( 
.A1(n_12658),
.A2(n_7219),
.A3(n_7245),
.B1(n_7194),
.B2(n_6980),
.Y(n_12885)
);

INVx2_ASAP7_75t_L g12886 ( 
.A(n_12479),
.Y(n_12886)
);

INVx2_ASAP7_75t_L g12887 ( 
.A(n_12474),
.Y(n_12887)
);

INVx1_ASAP7_75t_SL g12888 ( 
.A(n_12483),
.Y(n_12888)
);

NAND2xp33_ASAP7_75t_L g12889 ( 
.A(n_12376),
.B(n_8169),
.Y(n_12889)
);

OR2x2_ASAP7_75t_L g12890 ( 
.A(n_12488),
.B(n_12489),
.Y(n_12890)
);

INVx2_ASAP7_75t_SL g12891 ( 
.A(n_12669),
.Y(n_12891)
);

INVx1_ASAP7_75t_L g12892 ( 
.A(n_12532),
.Y(n_12892)
);

AND2x2_ASAP7_75t_L g12893 ( 
.A(n_12610),
.B(n_7219),
.Y(n_12893)
);

INVx1_ASAP7_75t_L g12894 ( 
.A(n_12546),
.Y(n_12894)
);

OAI332xp33_ASAP7_75t_L g12895 ( 
.A1(n_12636),
.A2(n_7024),
.A3(n_6462),
.B1(n_6279),
.B2(n_6435),
.B3(n_6358),
.C1(n_6436),
.C2(n_6315),
.Y(n_12895)
);

OR2x2_ASAP7_75t_L g12896 ( 
.A(n_12491),
.B(n_8170),
.Y(n_12896)
);

NAND2xp5_ASAP7_75t_L g12897 ( 
.A(n_12646),
.B(n_8173),
.Y(n_12897)
);

INVx1_ASAP7_75t_L g12898 ( 
.A(n_12549),
.Y(n_12898)
);

NOR3xp33_ASAP7_75t_L g12899 ( 
.A(n_12361),
.B(n_12541),
.C(n_12537),
.Y(n_12899)
);

INVx1_ASAP7_75t_L g12900 ( 
.A(n_12452),
.Y(n_12900)
);

INVx1_ASAP7_75t_L g12901 ( 
.A(n_12453),
.Y(n_12901)
);

NAND3xp33_ASAP7_75t_L g12902 ( 
.A(n_12437),
.B(n_7033),
.C(n_7225),
.Y(n_12902)
);

INVx1_ASAP7_75t_L g12903 ( 
.A(n_12458),
.Y(n_12903)
);

O2A1O1Ixp33_ASAP7_75t_L g12904 ( 
.A1(n_12656),
.A2(n_8177),
.B(n_8179),
.C(n_8173),
.Y(n_12904)
);

HB1xp67_ASAP7_75t_L g12905 ( 
.A(n_12607),
.Y(n_12905)
);

AND2x4_ASAP7_75t_L g12906 ( 
.A(n_12665),
.B(n_7219),
.Y(n_12906)
);

INVx2_ASAP7_75t_L g12907 ( 
.A(n_12631),
.Y(n_12907)
);

OR2x2_ASAP7_75t_L g12908 ( 
.A(n_12533),
.B(n_8177),
.Y(n_12908)
);

INVx1_ASAP7_75t_L g12909 ( 
.A(n_12536),
.Y(n_12909)
);

AND2x2_ASAP7_75t_L g12910 ( 
.A(n_12490),
.B(n_7245),
.Y(n_12910)
);

AND2x4_ASAP7_75t_L g12911 ( 
.A(n_12562),
.B(n_8179),
.Y(n_12911)
);

NAND2x1p5_ASAP7_75t_L g12912 ( 
.A(n_12548),
.B(n_6263),
.Y(n_12912)
);

OR2x2_ASAP7_75t_L g12913 ( 
.A(n_12438),
.B(n_8180),
.Y(n_12913)
);

INVxp67_ASAP7_75t_SL g12914 ( 
.A(n_12643),
.Y(n_12914)
);

INVx2_ASAP7_75t_L g12915 ( 
.A(n_12517),
.Y(n_12915)
);

INVx1_ASAP7_75t_L g12916 ( 
.A(n_12545),
.Y(n_12916)
);

OR2x2_ASAP7_75t_L g12917 ( 
.A(n_12440),
.B(n_8180),
.Y(n_12917)
);

NAND2xp5_ASAP7_75t_L g12918 ( 
.A(n_12618),
.B(n_8183),
.Y(n_12918)
);

OA21x2_ASAP7_75t_L g12919 ( 
.A1(n_12569),
.A2(n_8187),
.B(n_8183),
.Y(n_12919)
);

INVx1_ASAP7_75t_L g12920 ( 
.A(n_12558),
.Y(n_12920)
);

INVx1_ASAP7_75t_L g12921 ( 
.A(n_12667),
.Y(n_12921)
);

NAND2xp5_ASAP7_75t_L g12922 ( 
.A(n_12622),
.B(n_8187),
.Y(n_12922)
);

INVx1_ASAP7_75t_L g12923 ( 
.A(n_12633),
.Y(n_12923)
);

INVx1_ASAP7_75t_SL g12924 ( 
.A(n_12504),
.Y(n_12924)
);

INVx2_ASAP7_75t_L g12925 ( 
.A(n_12556),
.Y(n_12925)
);

AND2x2_ASAP7_75t_L g12926 ( 
.A(n_12505),
.B(n_7245),
.Y(n_12926)
);

AND2x2_ASAP7_75t_L g12927 ( 
.A(n_12476),
.B(n_7245),
.Y(n_12927)
);

INVx1_ASAP7_75t_L g12928 ( 
.A(n_12641),
.Y(n_12928)
);

INVx1_ASAP7_75t_L g12929 ( 
.A(n_12645),
.Y(n_12929)
);

INVx2_ASAP7_75t_SL g12930 ( 
.A(n_12580),
.Y(n_12930)
);

AND2x4_ASAP7_75t_L g12931 ( 
.A(n_12620),
.B(n_7245),
.Y(n_12931)
);

INVxp67_ASAP7_75t_L g12932 ( 
.A(n_12448),
.Y(n_12932)
);

OAI332xp33_ASAP7_75t_L g12933 ( 
.A1(n_12486),
.A2(n_6462),
.A3(n_6279),
.B1(n_6435),
.B2(n_6358),
.B3(n_6436),
.C1(n_6315),
.C2(n_6454),
.Y(n_12933)
);

O2A1O1Ixp33_ASAP7_75t_L g12934 ( 
.A1(n_12454),
.A2(n_8194),
.B(n_8202),
.C(n_8192),
.Y(n_12934)
);

INVxp67_ASAP7_75t_L g12935 ( 
.A(n_12477),
.Y(n_12935)
);

INVx2_ASAP7_75t_L g12936 ( 
.A(n_12609),
.Y(n_12936)
);

INVx2_ASAP7_75t_L g12937 ( 
.A(n_12538),
.Y(n_12937)
);

INVx1_ASAP7_75t_L g12938 ( 
.A(n_12463),
.Y(n_12938)
);

AOI22xp5_ASAP7_75t_L g12939 ( 
.A1(n_12586),
.A2(n_7347),
.B1(n_7285),
.B2(n_8192),
.Y(n_12939)
);

INVx2_ASAP7_75t_L g12940 ( 
.A(n_12547),
.Y(n_12940)
);

NAND2xp5_ASAP7_75t_L g12941 ( 
.A(n_12568),
.B(n_8194),
.Y(n_12941)
);

NAND4xp75_ASAP7_75t_L g12942 ( 
.A(n_12456),
.B(n_6503),
.C(n_7033),
.D(n_7023),
.Y(n_12942)
);

AND2x4_ASAP7_75t_L g12943 ( 
.A(n_12578),
.B(n_8202),
.Y(n_12943)
);

AOI21xp5_ASAP7_75t_SL g12944 ( 
.A1(n_12566),
.A2(n_7033),
.B(n_8204),
.Y(n_12944)
);

INVx1_ASAP7_75t_L g12945 ( 
.A(n_12499),
.Y(n_12945)
);

INVx1_ASAP7_75t_L g12946 ( 
.A(n_12511),
.Y(n_12946)
);

OR2x2_ASAP7_75t_L g12947 ( 
.A(n_12508),
.B(n_8204),
.Y(n_12947)
);

AND2x4_ASAP7_75t_L g12948 ( 
.A(n_12655),
.B(n_8213),
.Y(n_12948)
);

INVxp67_ASAP7_75t_SL g12949 ( 
.A(n_12583),
.Y(n_12949)
);

INVx1_ASAP7_75t_L g12950 ( 
.A(n_12611),
.Y(n_12950)
);

AOI22xp5_ASAP7_75t_L g12951 ( 
.A1(n_12588),
.A2(n_7285),
.B1(n_7347),
.B2(n_8213),
.Y(n_12951)
);

NAND3xp33_ASAP7_75t_L g12952 ( 
.A(n_12626),
.B(n_7033),
.C(n_7225),
.Y(n_12952)
);

INVx1_ASAP7_75t_L g12953 ( 
.A(n_12621),
.Y(n_12953)
);

NOR2xp33_ASAP7_75t_SL g12954 ( 
.A(n_12571),
.B(n_12576),
.Y(n_12954)
);

INVx1_ASAP7_75t_L g12955 ( 
.A(n_12634),
.Y(n_12955)
);

INVx2_ASAP7_75t_SL g12956 ( 
.A(n_12580),
.Y(n_12956)
);

INVx1_ASAP7_75t_L g12957 ( 
.A(n_12635),
.Y(n_12957)
);

AND2x2_ASAP7_75t_L g12958 ( 
.A(n_12516),
.B(n_7285),
.Y(n_12958)
);

INVx2_ASAP7_75t_L g12959 ( 
.A(n_12652),
.Y(n_12959)
);

A2O1A1Ixp33_ASAP7_75t_L g12960 ( 
.A1(n_12446),
.A2(n_6537),
.B(n_6535),
.C(n_6602),
.Y(n_12960)
);

AND2x2_ASAP7_75t_L g12961 ( 
.A(n_12563),
.B(n_7285),
.Y(n_12961)
);

NAND2xp5_ASAP7_75t_L g12962 ( 
.A(n_12779),
.B(n_12663),
.Y(n_12962)
);

OR2x2_ASAP7_75t_L g12963 ( 
.A(n_12791),
.B(n_12651),
.Y(n_12963)
);

OR2x2_ASAP7_75t_L g12964 ( 
.A(n_12723),
.B(n_12592),
.Y(n_12964)
);

INVx1_ASAP7_75t_L g12965 ( 
.A(n_12779),
.Y(n_12965)
);

AND2x4_ASAP7_75t_L g12966 ( 
.A(n_12674),
.B(n_12523),
.Y(n_12966)
);

INVx1_ASAP7_75t_L g12967 ( 
.A(n_12678),
.Y(n_12967)
);

INVx1_ASAP7_75t_L g12968 ( 
.A(n_12730),
.Y(n_12968)
);

OR2x2_ASAP7_75t_L g12969 ( 
.A(n_12807),
.B(n_12628),
.Y(n_12969)
);

INVx1_ASAP7_75t_L g12970 ( 
.A(n_12794),
.Y(n_12970)
);

INVx1_ASAP7_75t_L g12971 ( 
.A(n_12728),
.Y(n_12971)
);

INVx1_ASAP7_75t_L g12972 ( 
.A(n_12914),
.Y(n_12972)
);

AND2x2_ASAP7_75t_L g12973 ( 
.A(n_12812),
.B(n_12472),
.Y(n_12973)
);

INVx1_ASAP7_75t_L g12974 ( 
.A(n_12679),
.Y(n_12974)
);

AND2x2_ASAP7_75t_L g12975 ( 
.A(n_12687),
.B(n_12680),
.Y(n_12975)
);

INVx2_ASAP7_75t_L g12976 ( 
.A(n_12764),
.Y(n_12976)
);

INVx2_ASAP7_75t_L g12977 ( 
.A(n_12744),
.Y(n_12977)
);

INVx1_ASAP7_75t_L g12978 ( 
.A(n_12671),
.Y(n_12978)
);

NAND5xp2_ASAP7_75t_L g12979 ( 
.A(n_12684),
.B(n_12400),
.C(n_12559),
.D(n_12561),
.E(n_12560),
.Y(n_12979)
);

OR2x2_ASAP7_75t_L g12980 ( 
.A(n_12778),
.B(n_12642),
.Y(n_12980)
);

AND2x2_ASAP7_75t_L g12981 ( 
.A(n_12692),
.B(n_12473),
.Y(n_12981)
);

NAND2x1p5_ASAP7_75t_L g12982 ( 
.A(n_12837),
.B(n_12564),
.Y(n_12982)
);

INVxp67_ASAP7_75t_L g12983 ( 
.A(n_12905),
.Y(n_12983)
);

AND2x2_ASAP7_75t_L g12984 ( 
.A(n_12735),
.B(n_12593),
.Y(n_12984)
);

AND2x2_ASAP7_75t_L g12985 ( 
.A(n_12705),
.B(n_12653),
.Y(n_12985)
);

NAND2xp5_ASAP7_75t_L g12986 ( 
.A(n_12676),
.B(n_12638),
.Y(n_12986)
);

INVx1_ASAP7_75t_L g12987 ( 
.A(n_12686),
.Y(n_12987)
);

INVx2_ASAP7_75t_L g12988 ( 
.A(n_12855),
.Y(n_12988)
);

BUFx2_ASAP7_75t_L g12989 ( 
.A(n_12780),
.Y(n_12989)
);

NAND2xp5_ASAP7_75t_L g12990 ( 
.A(n_12688),
.B(n_12640),
.Y(n_12990)
);

NAND2xp5_ASAP7_75t_L g12991 ( 
.A(n_12722),
.B(n_12600),
.Y(n_12991)
);

INVxp67_ASAP7_75t_L g12992 ( 
.A(n_12954),
.Y(n_12992)
);

INVx4_ASAP7_75t_L g12993 ( 
.A(n_12856),
.Y(n_12993)
);

AND2x2_ASAP7_75t_L g12994 ( 
.A(n_12801),
.B(n_12657),
.Y(n_12994)
);

NAND2xp5_ASAP7_75t_L g12995 ( 
.A(n_12724),
.B(n_12739),
.Y(n_12995)
);

OR2x6_ASAP7_75t_L g12996 ( 
.A(n_12760),
.B(n_12575),
.Y(n_12996)
);

HB1xp67_ASAP7_75t_L g12997 ( 
.A(n_12741),
.Y(n_12997)
);

INVx1_ASAP7_75t_L g12998 ( 
.A(n_12797),
.Y(n_12998)
);

AND2x2_ASAP7_75t_L g12999 ( 
.A(n_12856),
.B(n_12567),
.Y(n_12999)
);

NAND5xp2_ASAP7_75t_L g13000 ( 
.A(n_12670),
.B(n_12624),
.C(n_12623),
.D(n_12596),
.E(n_12492),
.Y(n_13000)
);

INVx1_ASAP7_75t_L g13001 ( 
.A(n_12793),
.Y(n_13001)
);

INVx1_ASAP7_75t_SL g13002 ( 
.A(n_12677),
.Y(n_13002)
);

INVx1_ASAP7_75t_L g13003 ( 
.A(n_12843),
.Y(n_13003)
);

HB1xp67_ASAP7_75t_L g13004 ( 
.A(n_12693),
.Y(n_13004)
);

OR2x2_ASAP7_75t_L g13005 ( 
.A(n_12695),
.B(n_12660),
.Y(n_13005)
);

INVx5_ASAP7_75t_L g13006 ( 
.A(n_12854),
.Y(n_13006)
);

OR2x2_ASAP7_75t_L g13007 ( 
.A(n_12930),
.B(n_12613),
.Y(n_13007)
);

BUFx2_ASAP7_75t_L g13008 ( 
.A(n_12756),
.Y(n_13008)
);

OR2x2_ASAP7_75t_L g13009 ( 
.A(n_12956),
.B(n_12613),
.Y(n_13009)
);

NOR2x1_ASAP7_75t_L g13010 ( 
.A(n_12824),
.B(n_12581),
.Y(n_13010)
);

NAND4xp25_ASAP7_75t_L g13011 ( 
.A(n_12694),
.B(n_12629),
.C(n_12582),
.D(n_12603),
.Y(n_13011)
);

INVx1_ASAP7_75t_L g13012 ( 
.A(n_12766),
.Y(n_13012)
);

AND2x2_ASAP7_75t_L g13013 ( 
.A(n_12732),
.B(n_12659),
.Y(n_13013)
);

NOR2xp33_ASAP7_75t_R g13014 ( 
.A(n_12747),
.B(n_12598),
.Y(n_13014)
);

INVx1_ASAP7_75t_L g13015 ( 
.A(n_12698),
.Y(n_13015)
);

AOI22x1_ASAP7_75t_L g13016 ( 
.A1(n_12949),
.A2(n_12470),
.B1(n_12602),
.B2(n_12664),
.Y(n_13016)
);

INVx1_ASAP7_75t_L g13017 ( 
.A(n_12769),
.Y(n_13017)
);

INVx2_ASAP7_75t_L g13018 ( 
.A(n_12805),
.Y(n_13018)
);

OAI31xp33_ASAP7_75t_L g13019 ( 
.A1(n_12864),
.A2(n_12597),
.A3(n_12612),
.B(n_12599),
.Y(n_13019)
);

INVx1_ASAP7_75t_L g13020 ( 
.A(n_12701),
.Y(n_13020)
);

INVx1_ASAP7_75t_L g13021 ( 
.A(n_12783),
.Y(n_13021)
);

NAND2xp5_ASAP7_75t_L g13022 ( 
.A(n_12818),
.B(n_12608),
.Y(n_13022)
);

AND2x2_ASAP7_75t_L g13023 ( 
.A(n_12729),
.B(n_12661),
.Y(n_13023)
);

INVx1_ASAP7_75t_L g13024 ( 
.A(n_12771),
.Y(n_13024)
);

NAND2xp5_ASAP7_75t_L g13025 ( 
.A(n_12888),
.B(n_12661),
.Y(n_13025)
);

NOR3xp33_ASAP7_75t_SL g13026 ( 
.A(n_12738),
.B(n_12668),
.C(n_12627),
.Y(n_13026)
);

INVx1_ASAP7_75t_L g13027 ( 
.A(n_12890),
.Y(n_13027)
);

NAND3xp33_ASAP7_75t_L g13028 ( 
.A(n_12899),
.B(n_12507),
.C(n_12481),
.Y(n_13028)
);

OR2x2_ASAP7_75t_L g13029 ( 
.A(n_12808),
.B(n_12614),
.Y(n_13029)
);

NOR2x1_ASAP7_75t_L g13030 ( 
.A(n_12781),
.B(n_12614),
.Y(n_13030)
);

OR2x6_ASAP7_75t_L g13031 ( 
.A(n_12826),
.B(n_12627),
.Y(n_13031)
);

HB1xp67_ASAP7_75t_L g13032 ( 
.A(n_12876),
.Y(n_13032)
);

INVx1_ASAP7_75t_L g13033 ( 
.A(n_12681),
.Y(n_13033)
);

INVx4_ASAP7_75t_L g13034 ( 
.A(n_12719),
.Y(n_13034)
);

AOI21xp33_ASAP7_75t_L g13035 ( 
.A1(n_12862),
.A2(n_12417),
.B(n_6479),
.Y(n_13035)
);

INVx1_ASAP7_75t_L g13036 ( 
.A(n_12863),
.Y(n_13036)
);

INVx1_ASAP7_75t_L g13037 ( 
.A(n_12836),
.Y(n_13037)
);

OR2x4_ASAP7_75t_L g13038 ( 
.A(n_12806),
.B(n_6513),
.Y(n_13038)
);

INVx1_ASAP7_75t_L g13039 ( 
.A(n_12867),
.Y(n_13039)
);

AND2x2_ASAP7_75t_L g13040 ( 
.A(n_12798),
.B(n_7285),
.Y(n_13040)
);

OR2x2_ASAP7_75t_L g13041 ( 
.A(n_12696),
.B(n_8216),
.Y(n_13041)
);

INVx2_ASAP7_75t_L g13042 ( 
.A(n_12847),
.Y(n_13042)
);

NOR2xp33_ASAP7_75t_L g13043 ( 
.A(n_12689),
.B(n_8216),
.Y(n_13043)
);

INVx2_ASAP7_75t_L g13044 ( 
.A(n_12841),
.Y(n_13044)
);

AND2x2_ASAP7_75t_L g13045 ( 
.A(n_12710),
.B(n_7347),
.Y(n_13045)
);

OR2x2_ASAP7_75t_L g13046 ( 
.A(n_12702),
.B(n_8230),
.Y(n_13046)
);

INVx2_ASAP7_75t_L g13047 ( 
.A(n_12827),
.Y(n_13047)
);

INVx2_ASAP7_75t_L g13048 ( 
.A(n_12853),
.Y(n_13048)
);

INVx2_ASAP7_75t_L g13049 ( 
.A(n_12878),
.Y(n_13049)
);

INVx1_ASAP7_75t_L g13050 ( 
.A(n_12749),
.Y(n_13050)
);

INVx1_ASAP7_75t_L g13051 ( 
.A(n_12712),
.Y(n_13051)
);

AND2x2_ASAP7_75t_L g13052 ( 
.A(n_12795),
.B(n_7347),
.Y(n_13052)
);

NAND2xp5_ASAP7_75t_L g13053 ( 
.A(n_12718),
.B(n_8230),
.Y(n_13053)
);

OR2x2_ASAP7_75t_L g13054 ( 
.A(n_12721),
.B(n_8241),
.Y(n_13054)
);

AND2x2_ASAP7_75t_L g13055 ( 
.A(n_12725),
.B(n_7347),
.Y(n_13055)
);

INVx1_ASAP7_75t_L g13056 ( 
.A(n_12742),
.Y(n_13056)
);

AND2x4_ASAP7_75t_L g13057 ( 
.A(n_12887),
.B(n_8258),
.Y(n_13057)
);

INVx1_ASAP7_75t_L g13058 ( 
.A(n_12763),
.Y(n_13058)
);

OR2x2_ASAP7_75t_L g13059 ( 
.A(n_12834),
.B(n_8241),
.Y(n_13059)
);

BUFx2_ASAP7_75t_L g13060 ( 
.A(n_12802),
.Y(n_13060)
);

CKINVDCx16_ASAP7_75t_R g13061 ( 
.A(n_12675),
.Y(n_13061)
);

OR2x2_ASAP7_75t_L g13062 ( 
.A(n_12866),
.B(n_8242),
.Y(n_13062)
);

INVx1_ASAP7_75t_L g13063 ( 
.A(n_12751),
.Y(n_13063)
);

NAND2xp5_ASAP7_75t_L g13064 ( 
.A(n_12936),
.B(n_8242),
.Y(n_13064)
);

INVx1_ASAP7_75t_L g13065 ( 
.A(n_12757),
.Y(n_13065)
);

CKINVDCx16_ASAP7_75t_R g13066 ( 
.A(n_12672),
.Y(n_13066)
);

BUFx2_ASAP7_75t_L g13067 ( 
.A(n_12802),
.Y(n_13067)
);

OR2x2_ASAP7_75t_L g13068 ( 
.A(n_12770),
.B(n_8252),
.Y(n_13068)
);

NAND2xp5_ASAP7_75t_L g13069 ( 
.A(n_12865),
.B(n_8252),
.Y(n_13069)
);

OAI211xp5_ASAP7_75t_L g13070 ( 
.A1(n_12711),
.A2(n_6529),
.B(n_6266),
.C(n_6388),
.Y(n_13070)
);

NOR3xp33_ASAP7_75t_L g13071 ( 
.A(n_12683),
.B(n_6811),
.C(n_6809),
.Y(n_13071)
);

NAND2xp5_ASAP7_75t_L g13072 ( 
.A(n_12894),
.B(n_8257),
.Y(n_13072)
);

OR2x2_ASAP7_75t_L g13073 ( 
.A(n_12782),
.B(n_8257),
.Y(n_13073)
);

INVx1_ASAP7_75t_L g13074 ( 
.A(n_12880),
.Y(n_13074)
);

AND2x2_ASAP7_75t_L g13075 ( 
.A(n_12937),
.B(n_8258),
.Y(n_13075)
);

OR2x2_ASAP7_75t_L g13076 ( 
.A(n_12940),
.B(n_8267),
.Y(n_13076)
);

AND2x2_ASAP7_75t_L g13077 ( 
.A(n_12927),
.B(n_8267),
.Y(n_13077)
);

INVx2_ASAP7_75t_L g13078 ( 
.A(n_12861),
.Y(n_13078)
);

INVxp67_ASAP7_75t_L g13079 ( 
.A(n_12844),
.Y(n_13079)
);

INVx1_ASAP7_75t_L g13080 ( 
.A(n_12846),
.Y(n_13080)
);

INVxp67_ASAP7_75t_L g13081 ( 
.A(n_12898),
.Y(n_13081)
);

INVx1_ASAP7_75t_L g13082 ( 
.A(n_12673),
.Y(n_13082)
);

AOI22xp33_ASAP7_75t_L g13083 ( 
.A1(n_12839),
.A2(n_7277),
.B1(n_6535),
.B2(n_6604),
.Y(n_13083)
);

AND2x2_ASAP7_75t_L g13084 ( 
.A(n_12790),
.B(n_8270),
.Y(n_13084)
);

NAND2xp33_ASAP7_75t_SL g13085 ( 
.A(n_12871),
.B(n_6388),
.Y(n_13085)
);

INVxp67_ASAP7_75t_L g13086 ( 
.A(n_12682),
.Y(n_13086)
);

BUFx12f_ASAP7_75t_L g13087 ( 
.A(n_12838),
.Y(n_13087)
);

INVx1_ASAP7_75t_L g13088 ( 
.A(n_12726),
.Y(n_13088)
);

INVx2_ASAP7_75t_L g13089 ( 
.A(n_12919),
.Y(n_13089)
);

HB1xp67_ASAP7_75t_L g13090 ( 
.A(n_12746),
.Y(n_13090)
);

INVx1_ASAP7_75t_L g13091 ( 
.A(n_12768),
.Y(n_13091)
);

OR2x2_ASAP7_75t_L g13092 ( 
.A(n_12959),
.B(n_12874),
.Y(n_13092)
);

NAND2xp5_ASAP7_75t_L g13093 ( 
.A(n_12877),
.B(n_8270),
.Y(n_13093)
);

INVx2_ASAP7_75t_L g13094 ( 
.A(n_12919),
.Y(n_13094)
);

NAND2xp5_ASAP7_75t_L g13095 ( 
.A(n_12950),
.B(n_8271),
.Y(n_13095)
);

AOI21xp5_ASAP7_75t_L g13096 ( 
.A1(n_12889),
.A2(n_8324),
.B(n_8321),
.Y(n_13096)
);

NOR3xp33_ASAP7_75t_L g13097 ( 
.A(n_12804),
.B(n_6816),
.C(n_6811),
.Y(n_13097)
);

NAND2xp5_ASAP7_75t_L g13098 ( 
.A(n_12953),
.B(n_8271),
.Y(n_13098)
);

INVx1_ASAP7_75t_SL g13099 ( 
.A(n_12685),
.Y(n_13099)
);

INVx2_ASAP7_75t_SL g13100 ( 
.A(n_12931),
.Y(n_13100)
);

INVx2_ASAP7_75t_L g13101 ( 
.A(n_12833),
.Y(n_13101)
);

AND2x2_ASAP7_75t_L g13102 ( 
.A(n_12893),
.B(n_8272),
.Y(n_13102)
);

NAND2xp33_ASAP7_75t_R g13103 ( 
.A(n_12858),
.B(n_7225),
.Y(n_13103)
);

NAND2xp5_ASAP7_75t_L g13104 ( 
.A(n_12955),
.B(n_8272),
.Y(n_13104)
);

NOR2xp33_ASAP7_75t_L g13105 ( 
.A(n_12932),
.B(n_8273),
.Y(n_13105)
);

NAND2xp5_ASAP7_75t_L g13106 ( 
.A(n_12957),
.B(n_8273),
.Y(n_13106)
);

NAND2xp5_ASAP7_75t_L g13107 ( 
.A(n_12750),
.B(n_8274),
.Y(n_13107)
);

NAND2xp5_ASAP7_75t_L g13108 ( 
.A(n_12750),
.B(n_8274),
.Y(n_13108)
);

INVx1_ASAP7_75t_L g13109 ( 
.A(n_12875),
.Y(n_13109)
);

INVx1_ASAP7_75t_SL g13110 ( 
.A(n_12924),
.Y(n_13110)
);

INVxp67_ASAP7_75t_SL g13111 ( 
.A(n_12935),
.Y(n_13111)
);

NAND4xp25_ASAP7_75t_SL g13112 ( 
.A(n_12697),
.B(n_6979),
.C(n_7395),
.D(n_8275),
.Y(n_13112)
);

NAND2xp5_ASAP7_75t_L g13113 ( 
.A(n_12892),
.B(n_8275),
.Y(n_13113)
);

OAI22xp5_ASAP7_75t_L g13114 ( 
.A1(n_12809),
.A2(n_8303),
.B1(n_8320),
.B2(n_8278),
.Y(n_13114)
);

INVx1_ASAP7_75t_L g13115 ( 
.A(n_12703),
.Y(n_13115)
);

NAND2xp5_ASAP7_75t_L g13116 ( 
.A(n_12825),
.B(n_8276),
.Y(n_13116)
);

INVx1_ASAP7_75t_L g13117 ( 
.A(n_12690),
.Y(n_13117)
);

INVx2_ASAP7_75t_SL g13118 ( 
.A(n_12906),
.Y(n_13118)
);

INVx1_ASAP7_75t_L g13119 ( 
.A(n_12786),
.Y(n_13119)
);

NAND2xp5_ASAP7_75t_SL g13120 ( 
.A(n_12882),
.B(n_8276),
.Y(n_13120)
);

AND2x2_ASAP7_75t_L g13121 ( 
.A(n_12709),
.B(n_8278),
.Y(n_13121)
);

AND2x2_ASAP7_75t_L g13122 ( 
.A(n_12810),
.B(n_8284),
.Y(n_13122)
);

INVx1_ASAP7_75t_L g13123 ( 
.A(n_12773),
.Y(n_13123)
);

NOR2xp33_ASAP7_75t_R g13124 ( 
.A(n_12789),
.B(n_6263),
.Y(n_13124)
);

NAND2xp5_ASAP7_75t_L g13125 ( 
.A(n_12870),
.B(n_8284),
.Y(n_13125)
);

NAND2xp33_ASAP7_75t_SL g13126 ( 
.A(n_12774),
.B(n_8288),
.Y(n_13126)
);

OR2x2_ASAP7_75t_L g13127 ( 
.A(n_12840),
.B(n_8288),
.Y(n_13127)
);

NAND2xp5_ASAP7_75t_L g13128 ( 
.A(n_12900),
.B(n_8297),
.Y(n_13128)
);

AND2x2_ASAP7_75t_L g13129 ( 
.A(n_12886),
.B(n_8297),
.Y(n_13129)
);

NAND2xp5_ASAP7_75t_L g13130 ( 
.A(n_12901),
.B(n_12903),
.Y(n_13130)
);

AND2x2_ASAP7_75t_L g13131 ( 
.A(n_12851),
.B(n_8298),
.Y(n_13131)
);

NOR2xp33_ASAP7_75t_L g13132 ( 
.A(n_12754),
.B(n_8298),
.Y(n_13132)
);

AOI21xp5_ASAP7_75t_L g13133 ( 
.A1(n_12819),
.A2(n_8320),
.B(n_8317),
.Y(n_13133)
);

INVx2_ASAP7_75t_L g13134 ( 
.A(n_12833),
.Y(n_13134)
);

AND2x2_ASAP7_75t_L g13135 ( 
.A(n_12776),
.B(n_8303),
.Y(n_13135)
);

OR2x2_ASAP7_75t_L g13136 ( 
.A(n_12828),
.B(n_8308),
.Y(n_13136)
);

INVx2_ASAP7_75t_L g13137 ( 
.A(n_12761),
.Y(n_13137)
);

AND2x2_ASAP7_75t_SL g13138 ( 
.A(n_12822),
.B(n_6263),
.Y(n_13138)
);

OR2x2_ASAP7_75t_L g13139 ( 
.A(n_12758),
.B(n_8308),
.Y(n_13139)
);

INVx1_ASAP7_75t_L g13140 ( 
.A(n_12740),
.Y(n_13140)
);

OR2x2_ASAP7_75t_L g13141 ( 
.A(n_12762),
.B(n_8309),
.Y(n_13141)
);

INVx2_ASAP7_75t_L g13142 ( 
.A(n_12958),
.Y(n_13142)
);

NAND2xp5_ASAP7_75t_L g13143 ( 
.A(n_12909),
.B(n_8309),
.Y(n_13143)
);

NAND2x1_ASAP7_75t_L g13144 ( 
.A(n_12944),
.B(n_8310),
.Y(n_13144)
);

AND2x2_ASAP7_75t_L g13145 ( 
.A(n_12926),
.B(n_8310),
.Y(n_13145)
);

AOI21xp5_ASAP7_75t_L g13146 ( 
.A1(n_12691),
.A2(n_8327),
.B(n_8326),
.Y(n_13146)
);

INVx1_ASAP7_75t_L g13147 ( 
.A(n_12821),
.Y(n_13147)
);

INVx1_ASAP7_75t_L g13148 ( 
.A(n_12908),
.Y(n_13148)
);

NAND2xp5_ASAP7_75t_L g13149 ( 
.A(n_12916),
.B(n_8312),
.Y(n_13149)
);

INVx1_ASAP7_75t_L g13150 ( 
.A(n_12715),
.Y(n_13150)
);

INVx6_ASAP7_75t_L g13151 ( 
.A(n_12743),
.Y(n_13151)
);

OAI21xp5_ASAP7_75t_L g13152 ( 
.A1(n_12727),
.A2(n_6535),
.B(n_7514),
.Y(n_13152)
);

INVx1_ASAP7_75t_L g13153 ( 
.A(n_12799),
.Y(n_13153)
);

INVx1_ASAP7_75t_SL g13154 ( 
.A(n_12777),
.Y(n_13154)
);

BUFx3_ASAP7_75t_L g13155 ( 
.A(n_12920),
.Y(n_13155)
);

OR2x6_ASAP7_75t_L g13156 ( 
.A(n_12915),
.B(n_7799),
.Y(n_13156)
);

AO21x2_ASAP7_75t_L g13157 ( 
.A1(n_12938),
.A2(n_8313),
.B(n_8312),
.Y(n_13157)
);

INVxp67_ASAP7_75t_SL g13158 ( 
.A(n_12737),
.Y(n_13158)
);

BUFx3_ASAP7_75t_L g13159 ( 
.A(n_12945),
.Y(n_13159)
);

NAND2xp5_ASAP7_75t_L g13160 ( 
.A(n_12946),
.B(n_8313),
.Y(n_13160)
);

AND2x2_ASAP7_75t_L g13161 ( 
.A(n_12925),
.B(n_8317),
.Y(n_13161)
);

INVx2_ASAP7_75t_L g13162 ( 
.A(n_12947),
.Y(n_13162)
);

AND2x2_ASAP7_75t_L g13163 ( 
.A(n_12891),
.B(n_8321),
.Y(n_13163)
);

AND2x2_ASAP7_75t_L g13164 ( 
.A(n_12910),
.B(n_8324),
.Y(n_13164)
);

OR2x2_ASAP7_75t_L g13165 ( 
.A(n_12759),
.B(n_12775),
.Y(n_13165)
);

NOR2xp67_ASAP7_75t_L g13166 ( 
.A(n_12823),
.B(n_8326),
.Y(n_13166)
);

NOR2xp33_ASAP7_75t_L g13167 ( 
.A(n_12811),
.B(n_8327),
.Y(n_13167)
);

OR2x2_ASAP7_75t_L g13168 ( 
.A(n_12815),
.B(n_8330),
.Y(n_13168)
);

INVx1_ASAP7_75t_L g13169 ( 
.A(n_12816),
.Y(n_13169)
);

OR2x2_ASAP7_75t_L g13170 ( 
.A(n_12708),
.B(n_8330),
.Y(n_13170)
);

INVx1_ASAP7_75t_L g13171 ( 
.A(n_12913),
.Y(n_13171)
);

AND2x2_ASAP7_75t_L g13172 ( 
.A(n_12912),
.B(n_8331),
.Y(n_13172)
);

OR2x2_ASAP7_75t_L g13173 ( 
.A(n_12752),
.B(n_8331),
.Y(n_13173)
);

OR2x2_ASAP7_75t_L g13174 ( 
.A(n_12745),
.B(n_8335),
.Y(n_13174)
);

NAND2xp5_ASAP7_75t_L g13175 ( 
.A(n_12911),
.B(n_6462),
.Y(n_13175)
);

AND2x2_ASAP7_75t_L g13176 ( 
.A(n_12961),
.B(n_7277),
.Y(n_13176)
);

OAI211xp5_ASAP7_75t_SL g13177 ( 
.A1(n_12787),
.A2(n_7175),
.B(n_6979),
.C(n_7371),
.Y(n_13177)
);

INVx1_ASAP7_75t_L g13178 ( 
.A(n_12917),
.Y(n_13178)
);

CKINVDCx16_ASAP7_75t_R g13179 ( 
.A(n_12704),
.Y(n_13179)
);

INVx1_ASAP7_75t_SL g13180 ( 
.A(n_12814),
.Y(n_13180)
);

INVx3_ASAP7_75t_L g13181 ( 
.A(n_12911),
.Y(n_13181)
);

INVx1_ASAP7_75t_L g13182 ( 
.A(n_12896),
.Y(n_13182)
);

INVx2_ASAP7_75t_L g13183 ( 
.A(n_12873),
.Y(n_13183)
);

AND2x2_ASAP7_75t_L g13184 ( 
.A(n_12699),
.B(n_7277),
.Y(n_13184)
);

OR2x6_ASAP7_75t_L g13185 ( 
.A(n_12921),
.B(n_7864),
.Y(n_13185)
);

NAND2xp5_ASAP7_75t_L g13186 ( 
.A(n_12832),
.B(n_6462),
.Y(n_13186)
);

HB1xp67_ASAP7_75t_L g13187 ( 
.A(n_12907),
.Y(n_13187)
);

CKINVDCx5p33_ASAP7_75t_R g13188 ( 
.A(n_12929),
.Y(n_13188)
);

INVx1_ASAP7_75t_L g13189 ( 
.A(n_12788),
.Y(n_13189)
);

INVx1_ASAP7_75t_L g13190 ( 
.A(n_12817),
.Y(n_13190)
);

AND2x2_ASAP7_75t_L g13191 ( 
.A(n_12714),
.B(n_5707),
.Y(n_13191)
);

AND2x2_ASAP7_75t_L g13192 ( 
.A(n_12832),
.B(n_5707),
.Y(n_13192)
);

HB1xp67_ASAP7_75t_L g13193 ( 
.A(n_12943),
.Y(n_13193)
);

BUFx3_ASAP7_75t_L g13194 ( 
.A(n_12943),
.Y(n_13194)
);

INVx2_ASAP7_75t_SL g13195 ( 
.A(n_12753),
.Y(n_13195)
);

OAI21xp5_ASAP7_75t_SL g13196 ( 
.A1(n_12785),
.A2(n_7612),
.B(n_7450),
.Y(n_13196)
);

INVx2_ASAP7_75t_L g13197 ( 
.A(n_12948),
.Y(n_13197)
);

NAND2xp5_ASAP7_75t_L g13198 ( 
.A(n_12948),
.B(n_6462),
.Y(n_13198)
);

NAND2xp5_ASAP7_75t_L g13199 ( 
.A(n_12923),
.B(n_7225),
.Y(n_13199)
);

NAND2xp5_ASAP7_75t_L g13200 ( 
.A(n_12928),
.B(n_7244),
.Y(n_13200)
);

NOR2xp33_ASAP7_75t_R g13201 ( 
.A(n_12792),
.B(n_6263),
.Y(n_13201)
);

INVx2_ASAP7_75t_L g13202 ( 
.A(n_12942),
.Y(n_13202)
);

AND2x2_ASAP7_75t_L g13203 ( 
.A(n_12734),
.B(n_5707),
.Y(n_13203)
);

INVx1_ASAP7_75t_L g13204 ( 
.A(n_12884),
.Y(n_13204)
);

AOI221xp5_ASAP7_75t_SL g13205 ( 
.A1(n_12784),
.A2(n_7210),
.B1(n_7212),
.B2(n_7203),
.C(n_7199),
.Y(n_13205)
);

AND2x2_ASAP7_75t_L g13206 ( 
.A(n_12800),
.B(n_5718),
.Y(n_13206)
);

AOI22xp5_ASAP7_75t_L g13207 ( 
.A1(n_12713),
.A2(n_6929),
.B1(n_7341),
.B2(n_6841),
.Y(n_13207)
);

NAND2xp5_ASAP7_75t_L g13208 ( 
.A(n_12883),
.B(n_7244),
.Y(n_13208)
);

AND2x2_ASAP7_75t_L g13209 ( 
.A(n_12755),
.B(n_5718),
.Y(n_13209)
);

AND2x2_ASAP7_75t_L g13210 ( 
.A(n_12767),
.B(n_5718),
.Y(n_13210)
);

INVx2_ASAP7_75t_SL g13211 ( 
.A(n_12860),
.Y(n_13211)
);

AND2x2_ASAP7_75t_L g13212 ( 
.A(n_12720),
.B(n_5733),
.Y(n_13212)
);

INVx1_ASAP7_75t_L g13213 ( 
.A(n_12897),
.Y(n_13213)
);

INVx1_ASAP7_75t_L g13214 ( 
.A(n_12941),
.Y(n_13214)
);

NOR2x1_ASAP7_75t_L g13215 ( 
.A(n_12707),
.B(n_7244),
.Y(n_13215)
);

NOR2xp33_ASAP7_75t_R g13216 ( 
.A(n_12796),
.B(n_6984),
.Y(n_13216)
);

NAND4xp25_ASAP7_75t_L g13217 ( 
.A(n_12918),
.B(n_7386),
.C(n_7397),
.D(n_7273),
.Y(n_13217)
);

AND2x2_ASAP7_75t_L g13218 ( 
.A(n_12922),
.B(n_5733),
.Y(n_13218)
);

OR2x2_ASAP7_75t_L g13219 ( 
.A(n_12849),
.B(n_7244),
.Y(n_13219)
);

INVxp67_ASAP7_75t_L g13220 ( 
.A(n_12850),
.Y(n_13220)
);

NOR2xp33_ASAP7_75t_L g13221 ( 
.A(n_12933),
.B(n_6431),
.Y(n_13221)
);

NAND2xp33_ASAP7_75t_SL g13222 ( 
.A(n_12831),
.B(n_6578),
.Y(n_13222)
);

INVx1_ASAP7_75t_L g13223 ( 
.A(n_12904),
.Y(n_13223)
);

HB1xp67_ASAP7_75t_L g13224 ( 
.A(n_12716),
.Y(n_13224)
);

INVx1_ASAP7_75t_SL g13225 ( 
.A(n_12772),
.Y(n_13225)
);

NAND2xp5_ASAP7_75t_L g13226 ( 
.A(n_12934),
.B(n_7244),
.Y(n_13226)
);

INVx1_ASAP7_75t_L g13227 ( 
.A(n_12717),
.Y(n_13227)
);

AND2x2_ASAP7_75t_L g13228 ( 
.A(n_12857),
.B(n_5733),
.Y(n_13228)
);

OR2x2_ASAP7_75t_L g13229 ( 
.A(n_12879),
.B(n_5824),
.Y(n_13229)
);

INVx1_ASAP7_75t_L g13230 ( 
.A(n_12736),
.Y(n_13230)
);

OR2x2_ASAP7_75t_L g13231 ( 
.A(n_12902),
.B(n_5824),
.Y(n_13231)
);

OR2x2_ASAP7_75t_L g13232 ( 
.A(n_12952),
.B(n_5828),
.Y(n_13232)
);

AND2x2_ASAP7_75t_L g13233 ( 
.A(n_12706),
.B(n_5769),
.Y(n_13233)
);

NOR3xp33_ASAP7_75t_L g13234 ( 
.A(n_12748),
.B(n_6816),
.C(n_6668),
.Y(n_13234)
);

OAI211xp5_ASAP7_75t_SL g13235 ( 
.A1(n_12835),
.A2(n_7204),
.B(n_7186),
.C(n_7132),
.Y(n_13235)
);

NAND2xp5_ASAP7_75t_L g13236 ( 
.A(n_12848),
.B(n_5828),
.Y(n_13236)
);

INVx2_ASAP7_75t_SL g13237 ( 
.A(n_12803),
.Y(n_13237)
);

AND2x2_ASAP7_75t_L g13238 ( 
.A(n_12868),
.B(n_5769),
.Y(n_13238)
);

AND3x1_ASAP7_75t_L g13239 ( 
.A(n_12939),
.B(n_7203),
.C(n_7199),
.Y(n_13239)
);

INVx4_ASAP7_75t_L g13240 ( 
.A(n_12993),
.Y(n_13240)
);

NAND3xp33_ASAP7_75t_L g13241 ( 
.A(n_13019),
.B(n_12765),
.C(n_12951),
.Y(n_13241)
);

INVx1_ASAP7_75t_L g13242 ( 
.A(n_12973),
.Y(n_13242)
);

INVx1_ASAP7_75t_SL g13243 ( 
.A(n_12981),
.Y(n_13243)
);

INVxp67_ASAP7_75t_L g13244 ( 
.A(n_13004),
.Y(n_13244)
);

AND2x2_ASAP7_75t_L g13245 ( 
.A(n_12966),
.B(n_12881),
.Y(n_13245)
);

INVx1_ASAP7_75t_L g13246 ( 
.A(n_12975),
.Y(n_13246)
);

INVx1_ASAP7_75t_L g13247 ( 
.A(n_12971),
.Y(n_13247)
);

NAND2xp5_ASAP7_75t_L g13248 ( 
.A(n_13061),
.B(n_12895),
.Y(n_13248)
);

BUFx2_ASAP7_75t_L g13249 ( 
.A(n_13087),
.Y(n_13249)
);

OR2x2_ASAP7_75t_L g13250 ( 
.A(n_13066),
.B(n_12829),
.Y(n_13250)
);

INVx2_ASAP7_75t_L g13251 ( 
.A(n_13151),
.Y(n_13251)
);

INVx1_ASAP7_75t_SL g13252 ( 
.A(n_13002),
.Y(n_13252)
);

AO21x2_ASAP7_75t_L g13253 ( 
.A1(n_12965),
.A2(n_12960),
.B(n_12700),
.Y(n_13253)
);

INVx2_ASAP7_75t_L g13254 ( 
.A(n_13151),
.Y(n_13254)
);

AND2x2_ASAP7_75t_L g13255 ( 
.A(n_12966),
.B(n_12813),
.Y(n_13255)
);

HB1xp67_ASAP7_75t_L g13256 ( 
.A(n_13018),
.Y(n_13256)
);

INVx1_ASAP7_75t_SL g13257 ( 
.A(n_13099),
.Y(n_13257)
);

INVx1_ASAP7_75t_L g13258 ( 
.A(n_13008),
.Y(n_13258)
);

INVx2_ASAP7_75t_L g13259 ( 
.A(n_12969),
.Y(n_13259)
);

NOR2xp33_ASAP7_75t_L g13260 ( 
.A(n_12983),
.B(n_12731),
.Y(n_13260)
);

AND2x4_ASAP7_75t_L g13261 ( 
.A(n_13027),
.B(n_12852),
.Y(n_13261)
);

AND2x2_ASAP7_75t_L g13262 ( 
.A(n_13110),
.B(n_12820),
.Y(n_13262)
);

OR2x2_ASAP7_75t_L g13263 ( 
.A(n_12979),
.B(n_12733),
.Y(n_13263)
);

INVx1_ASAP7_75t_SL g13264 ( 
.A(n_12984),
.Y(n_13264)
);

INVx1_ASAP7_75t_SL g13265 ( 
.A(n_13007),
.Y(n_13265)
);

OAI22xp5_ASAP7_75t_L g13266 ( 
.A1(n_12998),
.A2(n_12845),
.B1(n_12859),
.B2(n_12830),
.Y(n_13266)
);

INVx3_ASAP7_75t_L g13267 ( 
.A(n_13034),
.Y(n_13267)
);

INVx1_ASAP7_75t_L g13268 ( 
.A(n_12997),
.Y(n_13268)
);

INVx1_ASAP7_75t_L g13269 ( 
.A(n_13089),
.Y(n_13269)
);

INVx1_ASAP7_75t_L g13270 ( 
.A(n_13094),
.Y(n_13270)
);

AOI22xp5_ASAP7_75t_L g13271 ( 
.A1(n_13103),
.A2(n_12872),
.B1(n_12869),
.B2(n_12885),
.Y(n_13271)
);

AND2x4_ASAP7_75t_L g13272 ( 
.A(n_13003),
.B(n_12842),
.Y(n_13272)
);

HB1xp67_ASAP7_75t_L g13273 ( 
.A(n_12976),
.Y(n_13273)
);

NAND3xp33_ASAP7_75t_L g13274 ( 
.A(n_12992),
.B(n_7205),
.C(n_6075),
.Y(n_13274)
);

CKINVDCx16_ASAP7_75t_R g13275 ( 
.A(n_13179),
.Y(n_13275)
);

HB1xp67_ASAP7_75t_L g13276 ( 
.A(n_13006),
.Y(n_13276)
);

INVx2_ASAP7_75t_L g13277 ( 
.A(n_12982),
.Y(n_13277)
);

AND2x2_ASAP7_75t_L g13278 ( 
.A(n_12988),
.B(n_5769),
.Y(n_13278)
);

INVxp67_ASAP7_75t_L g13279 ( 
.A(n_13010),
.Y(n_13279)
);

OR2x2_ASAP7_75t_L g13280 ( 
.A(n_12962),
.B(n_9111),
.Y(n_13280)
);

AOI22xp33_ASAP7_75t_L g13281 ( 
.A1(n_13000),
.A2(n_7808),
.B1(n_7855),
.B2(n_7799),
.Y(n_13281)
);

HB1xp67_ASAP7_75t_L g13282 ( 
.A(n_13006),
.Y(n_13282)
);

INVx4_ASAP7_75t_L g13283 ( 
.A(n_13006),
.Y(n_13283)
);

INVx2_ASAP7_75t_L g13284 ( 
.A(n_12980),
.Y(n_13284)
);

INVxp67_ASAP7_75t_SL g13285 ( 
.A(n_13030),
.Y(n_13285)
);

INVx1_ASAP7_75t_L g13286 ( 
.A(n_13193),
.Y(n_13286)
);

NOR2xp33_ASAP7_75t_L g13287 ( 
.A(n_13086),
.B(n_6258),
.Y(n_13287)
);

AND2x2_ASAP7_75t_L g13288 ( 
.A(n_12994),
.B(n_5772),
.Y(n_13288)
);

AND3x1_ASAP7_75t_L g13289 ( 
.A(n_13026),
.B(n_7212),
.C(n_7210),
.Y(n_13289)
);

NAND2xp5_ASAP7_75t_L g13290 ( 
.A(n_12974),
.B(n_9111),
.Y(n_13290)
);

INVx1_ASAP7_75t_L g13291 ( 
.A(n_12989),
.Y(n_13291)
);

OR2x2_ASAP7_75t_L g13292 ( 
.A(n_12978),
.B(n_9111),
.Y(n_13292)
);

AND2x4_ASAP7_75t_L g13293 ( 
.A(n_12977),
.B(n_8083),
.Y(n_13293)
);

INVx1_ASAP7_75t_SL g13294 ( 
.A(n_13009),
.Y(n_13294)
);

AND2x2_ASAP7_75t_L g13295 ( 
.A(n_12999),
.B(n_5772),
.Y(n_13295)
);

INVx1_ASAP7_75t_SL g13296 ( 
.A(n_12964),
.Y(n_13296)
);

NOR2x1_ASAP7_75t_L g13297 ( 
.A(n_13005),
.B(n_6578),
.Y(n_13297)
);

INVxp67_ASAP7_75t_L g13298 ( 
.A(n_13032),
.Y(n_13298)
);

BUFx3_ASAP7_75t_L g13299 ( 
.A(n_13048),
.Y(n_13299)
);

INVx1_ASAP7_75t_SL g13300 ( 
.A(n_13092),
.Y(n_13300)
);

INVx1_ASAP7_75t_SL g13301 ( 
.A(n_12963),
.Y(n_13301)
);

AOI221xp5_ASAP7_75t_L g13302 ( 
.A1(n_13028),
.A2(n_7227),
.B1(n_7229),
.B2(n_7226),
.C(n_7217),
.Y(n_13302)
);

NAND2x1p5_ASAP7_75t_L g13303 ( 
.A(n_13154),
.B(n_4782),
.Y(n_13303)
);

INVx1_ASAP7_75t_L g13304 ( 
.A(n_13049),
.Y(n_13304)
);

NAND2xp5_ASAP7_75t_L g13305 ( 
.A(n_13078),
.B(n_9111),
.Y(n_13305)
);

NOR2xp33_ASAP7_75t_L g13306 ( 
.A(n_12972),
.B(n_6258),
.Y(n_13306)
);

INVxp67_ASAP7_75t_L g13307 ( 
.A(n_12985),
.Y(n_13307)
);

INVx1_ASAP7_75t_L g13308 ( 
.A(n_12967),
.Y(n_13308)
);

NAND2xp5_ASAP7_75t_L g13309 ( 
.A(n_13181),
.B(n_9111),
.Y(n_13309)
);

BUFx3_ASAP7_75t_L g13310 ( 
.A(n_12968),
.Y(n_13310)
);

AND2x2_ASAP7_75t_L g13311 ( 
.A(n_13013),
.B(n_5772),
.Y(n_13311)
);

AOI222xp33_ASAP7_75t_L g13312 ( 
.A1(n_13215),
.A2(n_6530),
.B1(n_6455),
.B2(n_6547),
.C1(n_6524),
.C2(n_6488),
.Y(n_13312)
);

AOI22xp33_ASAP7_75t_L g13313 ( 
.A1(n_13042),
.A2(n_7855),
.B1(n_7864),
.B2(n_7808),
.Y(n_13313)
);

INVx2_ASAP7_75t_L g13314 ( 
.A(n_13194),
.Y(n_13314)
);

AOI222xp33_ASAP7_75t_L g13315 ( 
.A1(n_13225),
.A2(n_6530),
.B1(n_6455),
.B2(n_6547),
.C1(n_6524),
.C2(n_6488),
.Y(n_13315)
);

NAND2xp5_ASAP7_75t_L g13316 ( 
.A(n_13180),
.B(n_6454),
.Y(n_13316)
);

INVx1_ASAP7_75t_L g13317 ( 
.A(n_13165),
.Y(n_13317)
);

INVx1_ASAP7_75t_L g13318 ( 
.A(n_13111),
.Y(n_13318)
);

AND2x2_ASAP7_75t_L g13319 ( 
.A(n_13191),
.B(n_5774),
.Y(n_13319)
);

AOI22xp33_ASAP7_75t_L g13320 ( 
.A1(n_12996),
.A2(n_7855),
.B1(n_7864),
.B2(n_7808),
.Y(n_13320)
);

NAND2xp5_ASAP7_75t_L g13321 ( 
.A(n_13074),
.B(n_6454),
.Y(n_13321)
);

AND2x2_ASAP7_75t_L g13322 ( 
.A(n_13192),
.B(n_5774),
.Y(n_13322)
);

INVx1_ASAP7_75t_L g13323 ( 
.A(n_13025),
.Y(n_13323)
);

INVx1_ASAP7_75t_SL g13324 ( 
.A(n_13029),
.Y(n_13324)
);

INVx1_ASAP7_75t_L g13325 ( 
.A(n_13224),
.Y(n_13325)
);

INVx1_ASAP7_75t_L g13326 ( 
.A(n_13031),
.Y(n_13326)
);

OR2x2_ASAP7_75t_L g13327 ( 
.A(n_13011),
.B(n_12991),
.Y(n_13327)
);

HB1xp67_ASAP7_75t_L g13328 ( 
.A(n_13031),
.Y(n_13328)
);

AND2x2_ASAP7_75t_L g13329 ( 
.A(n_13052),
.B(n_5774),
.Y(n_13329)
);

OAI21x1_ASAP7_75t_L g13330 ( 
.A1(n_13016),
.A2(n_13044),
.B(n_13144),
.Y(n_13330)
);

OAI22xp5_ASAP7_75t_L g13331 ( 
.A1(n_13001),
.A2(n_7674),
.B1(n_7743),
.B2(n_7612),
.Y(n_13331)
);

AND2x2_ASAP7_75t_L g13332 ( 
.A(n_13218),
.B(n_5780),
.Y(n_13332)
);

AND2x2_ASAP7_75t_L g13333 ( 
.A(n_12970),
.B(n_5780),
.Y(n_13333)
);

INVx1_ASAP7_75t_L g13334 ( 
.A(n_12995),
.Y(n_13334)
);

INVx1_ASAP7_75t_L g13335 ( 
.A(n_12986),
.Y(n_13335)
);

INVx2_ASAP7_75t_L g13336 ( 
.A(n_13155),
.Y(n_13336)
);

NAND2xp5_ASAP7_75t_SL g13337 ( 
.A(n_13183),
.B(n_6513),
.Y(n_13337)
);

INVx1_ASAP7_75t_L g13338 ( 
.A(n_13036),
.Y(n_13338)
);

INVx1_ASAP7_75t_SL g13339 ( 
.A(n_13014),
.Y(n_13339)
);

AND2x4_ASAP7_75t_SL g13340 ( 
.A(n_13050),
.B(n_6984),
.Y(n_13340)
);

NAND2xp5_ASAP7_75t_L g13341 ( 
.A(n_13211),
.B(n_6454),
.Y(n_13341)
);

AND2x2_ASAP7_75t_L g13342 ( 
.A(n_13060),
.B(n_5780),
.Y(n_13342)
);

INVx2_ASAP7_75t_L g13343 ( 
.A(n_13159),
.Y(n_13343)
);

AND2x2_ASAP7_75t_L g13344 ( 
.A(n_13067),
.B(n_13212),
.Y(n_13344)
);

INVx2_ASAP7_75t_L g13345 ( 
.A(n_13157),
.Y(n_13345)
);

OAI21x1_ASAP7_75t_L g13346 ( 
.A1(n_13022),
.A2(n_7783),
.B(n_7720),
.Y(n_13346)
);

NOR2xp33_ASAP7_75t_L g13347 ( 
.A(n_13081),
.B(n_13079),
.Y(n_13347)
);

HB1xp67_ASAP7_75t_L g13348 ( 
.A(n_13090),
.Y(n_13348)
);

NAND3xp33_ASAP7_75t_L g13349 ( 
.A(n_13187),
.B(n_7205),
.C(n_6075),
.Y(n_13349)
);

INVxp67_ASAP7_75t_L g13350 ( 
.A(n_12990),
.Y(n_13350)
);

AND2x2_ASAP7_75t_L g13351 ( 
.A(n_13039),
.B(n_5805),
.Y(n_13351)
);

INVxp67_ASAP7_75t_L g13352 ( 
.A(n_12987),
.Y(n_13352)
);

OR2x2_ASAP7_75t_L g13353 ( 
.A(n_13162),
.B(n_6206),
.Y(n_13353)
);

INVx1_ASAP7_75t_L g13354 ( 
.A(n_13130),
.Y(n_13354)
);

INVx2_ASAP7_75t_L g13355 ( 
.A(n_13203),
.Y(n_13355)
);

INVxp67_ASAP7_75t_SL g13356 ( 
.A(n_13189),
.Y(n_13356)
);

INVx1_ASAP7_75t_SL g13357 ( 
.A(n_13023),
.Y(n_13357)
);

NOR2x1_ASAP7_75t_L g13358 ( 
.A(n_13012),
.B(n_7217),
.Y(n_13358)
);

OAI22xp5_ASAP7_75t_L g13359 ( 
.A1(n_13015),
.A2(n_7743),
.B1(n_7749),
.B2(n_7674),
.Y(n_13359)
);

INVx1_ASAP7_75t_L g13360 ( 
.A(n_13123),
.Y(n_13360)
);

AND2x2_ASAP7_75t_L g13361 ( 
.A(n_13055),
.B(n_5805),
.Y(n_13361)
);

NAND2xp5_ASAP7_75t_L g13362 ( 
.A(n_13195),
.B(n_6454),
.Y(n_13362)
);

NAND2xp5_ASAP7_75t_L g13363 ( 
.A(n_13171),
.B(n_6454),
.Y(n_13363)
);

AOI22xp33_ASAP7_75t_L g13364 ( 
.A1(n_12996),
.A2(n_8006),
.B1(n_8016),
.B2(n_7940),
.Y(n_13364)
);

OAI22xp5_ASAP7_75t_L g13365 ( 
.A1(n_13033),
.A2(n_7743),
.B1(n_7749),
.B2(n_7674),
.Y(n_13365)
);

NAND2xp5_ASAP7_75t_L g13366 ( 
.A(n_13178),
.B(n_13150),
.Y(n_13366)
);

OR2x2_ASAP7_75t_L g13367 ( 
.A(n_13037),
.B(n_6314),
.Y(n_13367)
);

INVx1_ASAP7_75t_L g13368 ( 
.A(n_13017),
.Y(n_13368)
);

NAND2xp5_ASAP7_75t_L g13369 ( 
.A(n_13182),
.B(n_6454),
.Y(n_13369)
);

NAND2xp5_ASAP7_75t_L g13370 ( 
.A(n_13147),
.B(n_6354),
.Y(n_13370)
);

NAND2xp5_ASAP7_75t_L g13371 ( 
.A(n_13169),
.B(n_6354),
.Y(n_13371)
);

INVx2_ASAP7_75t_L g13372 ( 
.A(n_13170),
.Y(n_13372)
);

AND2x2_ASAP7_75t_L g13373 ( 
.A(n_13024),
.B(n_5805),
.Y(n_13373)
);

OR2x2_ASAP7_75t_L g13374 ( 
.A(n_13109),
.B(n_6314),
.Y(n_13374)
);

INVx1_ASAP7_75t_SL g13375 ( 
.A(n_13080),
.Y(n_13375)
);

AOI22xp33_ASAP7_75t_L g13376 ( 
.A1(n_13233),
.A2(n_8006),
.B1(n_8016),
.B2(n_7940),
.Y(n_13376)
);

AND2x2_ASAP7_75t_L g13377 ( 
.A(n_13047),
.B(n_6103),
.Y(n_13377)
);

AND2x2_ASAP7_75t_L g13378 ( 
.A(n_13020),
.B(n_6103),
.Y(n_13378)
);

INVx2_ASAP7_75t_L g13379 ( 
.A(n_13173),
.Y(n_13379)
);

AND2x2_ASAP7_75t_L g13380 ( 
.A(n_13051),
.B(n_6103),
.Y(n_13380)
);

NAND2xp5_ASAP7_75t_L g13381 ( 
.A(n_13119),
.B(n_6065),
.Y(n_13381)
);

OR2x2_ASAP7_75t_L g13382 ( 
.A(n_13056),
.B(n_6370),
.Y(n_13382)
);

INVx1_ASAP7_75t_SL g13383 ( 
.A(n_13021),
.Y(n_13383)
);

AND2x2_ASAP7_75t_L g13384 ( 
.A(n_13142),
.B(n_6118),
.Y(n_13384)
);

INVx2_ASAP7_75t_L g13385 ( 
.A(n_13038),
.Y(n_13385)
);

OR2x6_ASAP7_75t_L g13386 ( 
.A(n_13117),
.B(n_8265),
.Y(n_13386)
);

INVx1_ASAP7_75t_L g13387 ( 
.A(n_13129),
.Y(n_13387)
);

NOR2xp33_ASAP7_75t_L g13388 ( 
.A(n_13221),
.B(n_7749),
.Y(n_13388)
);

INVx1_ASAP7_75t_L g13389 ( 
.A(n_13127),
.Y(n_13389)
);

INVx1_ASAP7_75t_L g13390 ( 
.A(n_13168),
.Y(n_13390)
);

NAND2xp5_ASAP7_75t_L g13391 ( 
.A(n_13197),
.B(n_6065),
.Y(n_13391)
);

INVx1_ASAP7_75t_SL g13392 ( 
.A(n_13082),
.Y(n_13392)
);

AND2x2_ASAP7_75t_L g13393 ( 
.A(n_13209),
.B(n_6118),
.Y(n_13393)
);

AOI22xp33_ASAP7_75t_L g13394 ( 
.A1(n_13234),
.A2(n_8006),
.B1(n_8016),
.B2(n_7940),
.Y(n_13394)
);

AND2x4_ASAP7_75t_L g13395 ( 
.A(n_13100),
.B(n_8083),
.Y(n_13395)
);

AOI222xp33_ASAP7_75t_L g13396 ( 
.A1(n_13083),
.A2(n_6547),
.B1(n_6488),
.B2(n_6561),
.C1(n_6530),
.C2(n_6524),
.Y(n_13396)
);

INVx1_ASAP7_75t_SL g13397 ( 
.A(n_13063),
.Y(n_13397)
);

INVx1_ASAP7_75t_L g13398 ( 
.A(n_13084),
.Y(n_13398)
);

AND2x2_ASAP7_75t_L g13399 ( 
.A(n_13065),
.B(n_6118),
.Y(n_13399)
);

INVx1_ASAP7_75t_L g13400 ( 
.A(n_13161),
.Y(n_13400)
);

AND2x2_ASAP7_75t_L g13401 ( 
.A(n_13138),
.B(n_6132),
.Y(n_13401)
);

AOI22xp33_ASAP7_75t_L g13402 ( 
.A1(n_13071),
.A2(n_8167),
.B1(n_8265),
.B2(n_8138),
.Y(n_13402)
);

INVx3_ASAP7_75t_L g13403 ( 
.A(n_13185),
.Y(n_13403)
);

INVxp67_ASAP7_75t_L g13404 ( 
.A(n_13148),
.Y(n_13404)
);

AND2x2_ASAP7_75t_L g13405 ( 
.A(n_13058),
.B(n_6132),
.Y(n_13405)
);

INVx1_ASAP7_75t_L g13406 ( 
.A(n_13121),
.Y(n_13406)
);

INVx4_ASAP7_75t_L g13407 ( 
.A(n_13188),
.Y(n_13407)
);

OR2x6_ASAP7_75t_L g13408 ( 
.A(n_13101),
.B(n_8294),
.Y(n_13408)
);

HB1xp67_ASAP7_75t_L g13409 ( 
.A(n_13166),
.Y(n_13409)
);

INVx1_ASAP7_75t_L g13410 ( 
.A(n_13107),
.Y(n_13410)
);

AOI22xp5_ASAP7_75t_L g13411 ( 
.A1(n_13132),
.A2(n_6929),
.B1(n_7341),
.B2(n_6841),
.Y(n_13411)
);

INVx1_ASAP7_75t_L g13412 ( 
.A(n_13108),
.Y(n_13412)
);

INVx2_ASAP7_75t_L g13413 ( 
.A(n_13156),
.Y(n_13413)
);

OR2x6_ASAP7_75t_L g13414 ( 
.A(n_13134),
.B(n_8294),
.Y(n_13414)
);

NAND2xp5_ASAP7_75t_L g13415 ( 
.A(n_13118),
.B(n_13115),
.Y(n_13415)
);

NOR2x1p5_ASAP7_75t_L g13416 ( 
.A(n_13158),
.B(n_13137),
.Y(n_13416)
);

OAI22xp33_ASAP7_75t_L g13417 ( 
.A1(n_13227),
.A2(n_8294),
.B1(n_8138),
.B2(n_8265),
.Y(n_13417)
);

INVxp67_ASAP7_75t_SL g13418 ( 
.A(n_13220),
.Y(n_13418)
);

OR2x2_ASAP7_75t_L g13419 ( 
.A(n_13076),
.B(n_6370),
.Y(n_13419)
);

INVx1_ASAP7_75t_SL g13420 ( 
.A(n_13085),
.Y(n_13420)
);

AND2x4_ASAP7_75t_L g13421 ( 
.A(n_13091),
.B(n_8148),
.Y(n_13421)
);

NAND2xp5_ASAP7_75t_L g13422 ( 
.A(n_13135),
.B(n_7226),
.Y(n_13422)
);

NAND2xp5_ASAP7_75t_L g13423 ( 
.A(n_13122),
.B(n_7227),
.Y(n_13423)
);

INVx1_ASAP7_75t_L g13424 ( 
.A(n_13062),
.Y(n_13424)
);

NAND2xp5_ASAP7_75t_L g13425 ( 
.A(n_13075),
.B(n_7229),
.Y(n_13425)
);

INVx1_ASAP7_75t_SL g13426 ( 
.A(n_13153),
.Y(n_13426)
);

INVx1_ASAP7_75t_L g13427 ( 
.A(n_13136),
.Y(n_13427)
);

AND2x4_ASAP7_75t_SL g13428 ( 
.A(n_13163),
.B(n_7127),
.Y(n_13428)
);

NAND2xp33_ASAP7_75t_L g13429 ( 
.A(n_13124),
.B(n_6412),
.Y(n_13429)
);

OA21x2_ASAP7_75t_L g13430 ( 
.A1(n_13120),
.A2(n_7669),
.B(n_7636),
.Y(n_13430)
);

INVx1_ASAP7_75t_L g13431 ( 
.A(n_13139),
.Y(n_13431)
);

INVx1_ASAP7_75t_L g13432 ( 
.A(n_13141),
.Y(n_13432)
);

AND2x2_ASAP7_75t_L g13433 ( 
.A(n_13228),
.B(n_6132),
.Y(n_13433)
);

AOI22xp33_ASAP7_75t_L g13434 ( 
.A1(n_13097),
.A2(n_8167),
.B1(n_8138),
.B2(n_6589),
.Y(n_13434)
);

INVx1_ASAP7_75t_L g13435 ( 
.A(n_13059),
.Y(n_13435)
);

AND2x2_ASAP7_75t_L g13436 ( 
.A(n_13206),
.B(n_6136),
.Y(n_13436)
);

INVx1_ASAP7_75t_L g13437 ( 
.A(n_13068),
.Y(n_13437)
);

NAND2xp5_ASAP7_75t_SL g13438 ( 
.A(n_13202),
.B(n_6513),
.Y(n_13438)
);

HB1xp67_ASAP7_75t_L g13439 ( 
.A(n_13237),
.Y(n_13439)
);

OAI22xp5_ASAP7_75t_L g13440 ( 
.A1(n_13207),
.A2(n_13208),
.B1(n_13190),
.B2(n_13204),
.Y(n_13440)
);

INVx1_ASAP7_75t_L g13441 ( 
.A(n_13073),
.Y(n_13441)
);

INVx1_ASAP7_75t_SL g13442 ( 
.A(n_13213),
.Y(n_13442)
);

OR2x6_ASAP7_75t_L g13443 ( 
.A(n_13214),
.B(n_8167),
.Y(n_13443)
);

INVx2_ASAP7_75t_L g13444 ( 
.A(n_13156),
.Y(n_13444)
);

AND2x2_ASAP7_75t_L g13445 ( 
.A(n_13184),
.B(n_6136),
.Y(n_13445)
);

INVx1_ASAP7_75t_SL g13446 ( 
.A(n_13230),
.Y(n_13446)
);

NAND2xp5_ASAP7_75t_L g13447 ( 
.A(n_13057),
.B(n_7231),
.Y(n_13447)
);

INVx1_ASAP7_75t_L g13448 ( 
.A(n_13057),
.Y(n_13448)
);

OR2x2_ASAP7_75t_L g13449 ( 
.A(n_13236),
.B(n_6412),
.Y(n_13449)
);

NAND2xp5_ASAP7_75t_L g13450 ( 
.A(n_13102),
.B(n_7231),
.Y(n_13450)
);

BUFx2_ASAP7_75t_L g13451 ( 
.A(n_13201),
.Y(n_13451)
);

INVx1_ASAP7_75t_L g13452 ( 
.A(n_13041),
.Y(n_13452)
);

NOR2xp33_ASAP7_75t_L g13453 ( 
.A(n_13223),
.B(n_6561),
.Y(n_13453)
);

BUFx12f_ASAP7_75t_L g13454 ( 
.A(n_13046),
.Y(n_13454)
);

AND2x2_ASAP7_75t_L g13455 ( 
.A(n_13210),
.B(n_6136),
.Y(n_13455)
);

NAND2xp5_ASAP7_75t_L g13456 ( 
.A(n_13077),
.B(n_7232),
.Y(n_13456)
);

INVx1_ASAP7_75t_L g13457 ( 
.A(n_13054),
.Y(n_13457)
);

NAND2xp5_ASAP7_75t_L g13458 ( 
.A(n_13145),
.B(n_7232),
.Y(n_13458)
);

INVx2_ASAP7_75t_L g13459 ( 
.A(n_13185),
.Y(n_13459)
);

OR2x2_ASAP7_75t_L g13460 ( 
.A(n_13064),
.B(n_6416),
.Y(n_13460)
);

NOR2xp33_ASAP7_75t_L g13461 ( 
.A(n_13140),
.B(n_6561),
.Y(n_13461)
);

INVx4_ASAP7_75t_L g13462 ( 
.A(n_13088),
.Y(n_13462)
);

OAI21xp5_ASAP7_75t_L g13463 ( 
.A1(n_13279),
.A2(n_13043),
.B(n_13105),
.Y(n_13463)
);

AOI32xp33_ASAP7_75t_L g13464 ( 
.A1(n_13300),
.A2(n_13126),
.A3(n_13167),
.B1(n_13172),
.B2(n_13093),
.Y(n_13464)
);

OAI21xp33_ASAP7_75t_L g13465 ( 
.A1(n_13243),
.A2(n_13216),
.B(n_13112),
.Y(n_13465)
);

NAND2xp5_ASAP7_75t_L g13466 ( 
.A(n_13249),
.B(n_13164),
.Y(n_13466)
);

AND2x2_ASAP7_75t_L g13467 ( 
.A(n_13275),
.B(n_13040),
.Y(n_13467)
);

AOI21xp33_ASAP7_75t_L g13468 ( 
.A1(n_13317),
.A2(n_13200),
.B(n_13199),
.Y(n_13468)
);

INVxp67_ASAP7_75t_L g13469 ( 
.A(n_13256),
.Y(n_13469)
);

OAI22xp5_ASAP7_75t_L g13470 ( 
.A1(n_13244),
.A2(n_13219),
.B1(n_13231),
.B2(n_13232),
.Y(n_13470)
);

AND2x2_ASAP7_75t_L g13471 ( 
.A(n_13242),
.B(n_13045),
.Y(n_13471)
);

AND2x2_ASAP7_75t_L g13472 ( 
.A(n_13265),
.B(n_13131),
.Y(n_13472)
);

INVx1_ASAP7_75t_L g13473 ( 
.A(n_13273),
.Y(n_13473)
);

OAI221xp5_ASAP7_75t_SL g13474 ( 
.A1(n_13257),
.A2(n_13198),
.B1(n_13186),
.B2(n_13175),
.C(n_13116),
.Y(n_13474)
);

OAI211xp5_ASAP7_75t_L g13475 ( 
.A1(n_13285),
.A2(n_13125),
.B(n_13143),
.C(n_13128),
.Y(n_13475)
);

INVx1_ASAP7_75t_SL g13476 ( 
.A(n_13252),
.Y(n_13476)
);

NAND2xp5_ASAP7_75t_SL g13477 ( 
.A(n_13277),
.B(n_13069),
.Y(n_13477)
);

A2O1A1Ixp33_ASAP7_75t_L g13478 ( 
.A1(n_13260),
.A2(n_13347),
.B(n_13298),
.C(n_13248),
.Y(n_13478)
);

INVx1_ASAP7_75t_L g13479 ( 
.A(n_13276),
.Y(n_13479)
);

OR2x2_ASAP7_75t_L g13480 ( 
.A(n_13294),
.B(n_13296),
.Y(n_13480)
);

INVx1_ASAP7_75t_SL g13481 ( 
.A(n_13301),
.Y(n_13481)
);

HB1xp67_ASAP7_75t_L g13482 ( 
.A(n_13282),
.Y(n_13482)
);

AND2x2_ASAP7_75t_L g13483 ( 
.A(n_13240),
.B(n_13299),
.Y(n_13483)
);

AOI22xp5_ASAP7_75t_L g13484 ( 
.A1(n_13344),
.A2(n_13152),
.B1(n_13235),
.B2(n_13176),
.Y(n_13484)
);

OAI21xp5_ASAP7_75t_SL g13485 ( 
.A1(n_13264),
.A2(n_13035),
.B(n_13196),
.Y(n_13485)
);

OAI21xp5_ASAP7_75t_L g13486 ( 
.A1(n_13328),
.A2(n_13160),
.B(n_13149),
.Y(n_13486)
);

INVx1_ASAP7_75t_L g13487 ( 
.A(n_13348),
.Y(n_13487)
);

NAND2xp5_ASAP7_75t_L g13488 ( 
.A(n_13324),
.B(n_13146),
.Y(n_13488)
);

OAI21xp33_ASAP7_75t_L g13489 ( 
.A1(n_13325),
.A2(n_13113),
.B(n_13053),
.Y(n_13489)
);

OAI22xp33_ASAP7_75t_L g13490 ( 
.A1(n_13263),
.A2(n_13375),
.B1(n_13250),
.B2(n_13411),
.Y(n_13490)
);

OAI21xp33_ASAP7_75t_L g13491 ( 
.A1(n_13246),
.A2(n_13098),
.B(n_13095),
.Y(n_13491)
);

INVx2_ASAP7_75t_L g13492 ( 
.A(n_13283),
.Y(n_13492)
);

AOI221xp5_ASAP7_75t_L g13493 ( 
.A1(n_13269),
.A2(n_13072),
.B1(n_13106),
.B2(n_13104),
.C(n_13226),
.Y(n_13493)
);

AO21x1_ASAP7_75t_L g13494 ( 
.A1(n_13407),
.A2(n_13133),
.B(n_13222),
.Y(n_13494)
);

AOI22xp5_ASAP7_75t_L g13495 ( 
.A1(n_13318),
.A2(n_13239),
.B1(n_13070),
.B2(n_13229),
.Y(n_13495)
);

OAI221xp5_ASAP7_75t_L g13496 ( 
.A1(n_13326),
.A2(n_13205),
.B1(n_13174),
.B2(n_13096),
.C(n_13177),
.Y(n_13496)
);

NAND2xp5_ASAP7_75t_L g13497 ( 
.A(n_13357),
.B(n_13238),
.Y(n_13497)
);

INVx1_ASAP7_75t_L g13498 ( 
.A(n_13267),
.Y(n_13498)
);

OA21x2_ASAP7_75t_L g13499 ( 
.A1(n_13330),
.A2(n_13114),
.B(n_13217),
.Y(n_13499)
);

INVx2_ASAP7_75t_L g13500 ( 
.A(n_13284),
.Y(n_13500)
);

NAND2xp5_ASAP7_75t_L g13501 ( 
.A(n_13339),
.B(n_13259),
.Y(n_13501)
);

OR2x2_ASAP7_75t_L g13502 ( 
.A(n_13251),
.B(n_13254),
.Y(n_13502)
);

NAND2xp5_ASAP7_75t_L g13503 ( 
.A(n_13356),
.B(n_6757),
.Y(n_13503)
);

AOI32xp33_ASAP7_75t_L g13504 ( 
.A1(n_13289),
.A2(n_6816),
.A3(n_6604),
.B1(n_6602),
.B2(n_6818),
.Y(n_13504)
);

INVx2_ASAP7_75t_L g13505 ( 
.A(n_13303),
.Y(n_13505)
);

AOI21xp33_ASAP7_75t_L g13506 ( 
.A1(n_13268),
.A2(n_6610),
.B(n_6589),
.Y(n_13506)
);

INVx1_ASAP7_75t_L g13507 ( 
.A(n_13409),
.Y(n_13507)
);

AOI22xp5_ASAP7_75t_L g13508 ( 
.A1(n_13253),
.A2(n_6929),
.B1(n_7341),
.B2(n_6841),
.Y(n_13508)
);

AND2x4_ASAP7_75t_L g13509 ( 
.A(n_13416),
.B(n_8148),
.Y(n_13509)
);

OR2x2_ASAP7_75t_L g13510 ( 
.A(n_13392),
.B(n_6416),
.Y(n_13510)
);

AOI22xp5_ASAP7_75t_L g13511 ( 
.A1(n_13383),
.A2(n_6929),
.B1(n_7341),
.B2(n_6841),
.Y(n_13511)
);

INVx1_ASAP7_75t_SL g13512 ( 
.A(n_13397),
.Y(n_13512)
);

OAI22xp5_ASAP7_75t_L g13513 ( 
.A1(n_13352),
.A2(n_7241),
.B1(n_7254),
.B2(n_7239),
.Y(n_13513)
);

INVx1_ASAP7_75t_L g13514 ( 
.A(n_13278),
.Y(n_13514)
);

INVx1_ASAP7_75t_L g13515 ( 
.A(n_13304),
.Y(n_13515)
);

OAI21xp5_ASAP7_75t_L g13516 ( 
.A1(n_13307),
.A2(n_6629),
.B(n_6605),
.Y(n_13516)
);

AOI21xp5_ASAP7_75t_L g13517 ( 
.A1(n_13366),
.A2(n_7204),
.B(n_7186),
.Y(n_13517)
);

AOI21xp5_ASAP7_75t_L g13518 ( 
.A1(n_13415),
.A2(n_7107),
.B(n_7086),
.Y(n_13518)
);

O2A1O1Ixp33_ASAP7_75t_SL g13519 ( 
.A1(n_13258),
.A2(n_5634),
.B(n_5675),
.C(n_5587),
.Y(n_13519)
);

INVx1_ASAP7_75t_L g13520 ( 
.A(n_13291),
.Y(n_13520)
);

NOR2xp33_ASAP7_75t_SL g13521 ( 
.A(n_13336),
.B(n_7127),
.Y(n_13521)
);

INVx1_ASAP7_75t_L g13522 ( 
.A(n_13342),
.Y(n_13522)
);

INVx1_ASAP7_75t_L g13523 ( 
.A(n_13286),
.Y(n_13523)
);

AOI22xp5_ASAP7_75t_L g13524 ( 
.A1(n_13270),
.A2(n_6929),
.B1(n_7341),
.B2(n_6841),
.Y(n_13524)
);

INVx1_ASAP7_75t_L g13525 ( 
.A(n_13310),
.Y(n_13525)
);

INVx1_ASAP7_75t_L g13526 ( 
.A(n_13351),
.Y(n_13526)
);

OAI22xp5_ASAP7_75t_L g13527 ( 
.A1(n_13334),
.A2(n_7241),
.B1(n_7254),
.B2(n_7239),
.Y(n_13527)
);

NAND2xp5_ASAP7_75t_L g13528 ( 
.A(n_13288),
.B(n_6757),
.Y(n_13528)
);

NAND2xp5_ASAP7_75t_L g13529 ( 
.A(n_13311),
.B(n_6757),
.Y(n_13529)
);

NOR2xp33_ASAP7_75t_L g13530 ( 
.A(n_13446),
.B(n_6589),
.Y(n_13530)
);

INVx2_ASAP7_75t_L g13531 ( 
.A(n_13295),
.Y(n_13531)
);

AND2x2_ASAP7_75t_L g13532 ( 
.A(n_13373),
.B(n_6850),
.Y(n_13532)
);

INVxp67_ASAP7_75t_SL g13533 ( 
.A(n_13439),
.Y(n_13533)
);

OAI21xp5_ASAP7_75t_L g13534 ( 
.A1(n_13350),
.A2(n_6629),
.B(n_6605),
.Y(n_13534)
);

O2A1O1Ixp5_ASAP7_75t_L g13535 ( 
.A1(n_13343),
.A2(n_7255),
.B(n_7266),
.C(n_7263),
.Y(n_13535)
);

NOR3xp33_ASAP7_75t_SL g13536 ( 
.A(n_13241),
.B(n_5931),
.C(n_7103),
.Y(n_13536)
);

OAI22xp33_ASAP7_75t_SL g13537 ( 
.A1(n_13355),
.A2(n_6473),
.B1(n_6692),
.B2(n_6557),
.Y(n_13537)
);

OAI22xp33_ASAP7_75t_L g13538 ( 
.A1(n_13338),
.A2(n_6513),
.B1(n_6722),
.B2(n_6720),
.Y(n_13538)
);

INVx1_ASAP7_75t_L g13539 ( 
.A(n_13327),
.Y(n_13539)
);

INVxp67_ASAP7_75t_L g13540 ( 
.A(n_13245),
.Y(n_13540)
);

INVxp67_ASAP7_75t_L g13541 ( 
.A(n_13314),
.Y(n_13541)
);

INVx1_ASAP7_75t_SL g13542 ( 
.A(n_13426),
.Y(n_13542)
);

OAI22xp33_ASAP7_75t_SL g13543 ( 
.A1(n_13280),
.A2(n_6473),
.B1(n_6692),
.B2(n_6557),
.Y(n_13543)
);

INVx2_ASAP7_75t_L g13544 ( 
.A(n_13354),
.Y(n_13544)
);

OAI21xp33_ASAP7_75t_L g13545 ( 
.A1(n_13388),
.A2(n_7263),
.B(n_7255),
.Y(n_13545)
);

OAI22xp33_ASAP7_75t_L g13546 ( 
.A1(n_13385),
.A2(n_6513),
.B1(n_6722),
.B2(n_6720),
.Y(n_13546)
);

INVx1_ASAP7_75t_L g13547 ( 
.A(n_13333),
.Y(n_13547)
);

AOI22xp5_ASAP7_75t_L g13548 ( 
.A1(n_13418),
.A2(n_7343),
.B1(n_6473),
.B2(n_6692),
.Y(n_13548)
);

O2A1O1Ixp5_ASAP7_75t_L g13549 ( 
.A1(n_13462),
.A2(n_7266),
.B(n_7281),
.C(n_7268),
.Y(n_13549)
);

INVx1_ASAP7_75t_L g13550 ( 
.A(n_13247),
.Y(n_13550)
);

INVx2_ASAP7_75t_L g13551 ( 
.A(n_13454),
.Y(n_13551)
);

BUFx2_ASAP7_75t_L g13552 ( 
.A(n_13335),
.Y(n_13552)
);

INVxp67_ASAP7_75t_L g13553 ( 
.A(n_13255),
.Y(n_13553)
);

AND2x2_ASAP7_75t_L g13554 ( 
.A(n_13319),
.B(n_13378),
.Y(n_13554)
);

INVx1_ASAP7_75t_L g13555 ( 
.A(n_13345),
.Y(n_13555)
);

NAND2xp5_ASAP7_75t_L g13556 ( 
.A(n_13442),
.B(n_6757),
.Y(n_13556)
);

AND2x2_ASAP7_75t_L g13557 ( 
.A(n_13380),
.B(n_6850),
.Y(n_13557)
);

INVx1_ASAP7_75t_L g13558 ( 
.A(n_13368),
.Y(n_13558)
);

AND2x2_ASAP7_75t_L g13559 ( 
.A(n_13377),
.B(n_6850),
.Y(n_13559)
);

INVx2_ASAP7_75t_L g13560 ( 
.A(n_13372),
.Y(n_13560)
);

INVx2_ASAP7_75t_L g13561 ( 
.A(n_13379),
.Y(n_13561)
);

NAND2xp5_ASAP7_75t_L g13562 ( 
.A(n_13406),
.B(n_6757),
.Y(n_13562)
);

INVx1_ASAP7_75t_SL g13563 ( 
.A(n_13420),
.Y(n_13563)
);

OAI22xp5_ASAP7_75t_L g13564 ( 
.A1(n_13404),
.A2(n_7281),
.B1(n_7290),
.B2(n_7268),
.Y(n_13564)
);

INVx1_ASAP7_75t_L g13565 ( 
.A(n_13323),
.Y(n_13565)
);

INVx1_ASAP7_75t_L g13566 ( 
.A(n_13308),
.Y(n_13566)
);

OAI22xp5_ASAP7_75t_L g13567 ( 
.A1(n_13271),
.A2(n_7307),
.B1(n_7328),
.B2(n_7290),
.Y(n_13567)
);

OAI22xp33_ASAP7_75t_L g13568 ( 
.A1(n_13360),
.A2(n_6720),
.B1(n_6738),
.B2(n_6722),
.Y(n_13568)
);

INVx2_ASAP7_75t_L g13569 ( 
.A(n_13443),
.Y(n_13569)
);

NAND2xp5_ASAP7_75t_L g13570 ( 
.A(n_13427),
.B(n_6757),
.Y(n_13570)
);

AOI221xp5_ASAP7_75t_L g13571 ( 
.A1(n_13440),
.A2(n_7307),
.B1(n_7328),
.B2(n_6995),
.C(n_6916),
.Y(n_13571)
);

AOI22xp33_ASAP7_75t_SL g13572 ( 
.A1(n_13262),
.A2(n_6725),
.B1(n_6735),
.B2(n_6557),
.Y(n_13572)
);

OAI21xp5_ASAP7_75t_L g13573 ( 
.A1(n_13261),
.A2(n_6629),
.B(n_6605),
.Y(n_13573)
);

OAI32xp33_ASAP7_75t_L g13574 ( 
.A1(n_13353),
.A2(n_7138),
.A3(n_7149),
.B1(n_7064),
.B2(n_7045),
.Y(n_13574)
);

NAND2xp5_ASAP7_75t_L g13575 ( 
.A(n_13431),
.B(n_6757),
.Y(n_13575)
);

INVx1_ASAP7_75t_L g13576 ( 
.A(n_13432),
.Y(n_13576)
);

INVx1_ASAP7_75t_L g13577 ( 
.A(n_13389),
.Y(n_13577)
);

AOI22xp5_ASAP7_75t_L g13578 ( 
.A1(n_13261),
.A2(n_7343),
.B1(n_6735),
.B2(n_6741),
.Y(n_13578)
);

INVx1_ASAP7_75t_L g13579 ( 
.A(n_13424),
.Y(n_13579)
);

AOI22xp33_ASAP7_75t_SL g13580 ( 
.A1(n_13413),
.A2(n_6735),
.B1(n_6741),
.B2(n_6725),
.Y(n_13580)
);

AOI21xp33_ASAP7_75t_L g13581 ( 
.A1(n_13305),
.A2(n_6626),
.B(n_6610),
.Y(n_13581)
);

NOR2xp33_ASAP7_75t_L g13582 ( 
.A(n_13403),
.B(n_6610),
.Y(n_13582)
);

NAND2xp5_ASAP7_75t_L g13583 ( 
.A(n_13435),
.B(n_13452),
.Y(n_13583)
);

AOI22xp5_ASAP7_75t_L g13584 ( 
.A1(n_13437),
.A2(n_7343),
.B1(n_6741),
.B2(n_6751),
.Y(n_13584)
);

INVx1_ASAP7_75t_L g13585 ( 
.A(n_13448),
.Y(n_13585)
);

NAND2xp5_ASAP7_75t_L g13586 ( 
.A(n_13457),
.B(n_6499),
.Y(n_13586)
);

OAI21xp33_ASAP7_75t_L g13587 ( 
.A1(n_13287),
.A2(n_13340),
.B(n_13297),
.Y(n_13587)
);

AOI22xp5_ASAP7_75t_L g13588 ( 
.A1(n_13441),
.A2(n_7343),
.B1(n_6751),
.B2(n_6754),
.Y(n_13588)
);

INVx1_ASAP7_75t_L g13589 ( 
.A(n_13399),
.Y(n_13589)
);

NAND2xp5_ASAP7_75t_L g13590 ( 
.A(n_13387),
.B(n_6499),
.Y(n_13590)
);

AOI322xp5_ASAP7_75t_L g13591 ( 
.A1(n_13316),
.A2(n_7240),
.A3(n_6499),
.B1(n_6086),
.B2(n_6062),
.C1(n_7103),
.C2(n_7172),
.Y(n_13591)
);

OAI21xp5_ASAP7_75t_L g13592 ( 
.A1(n_13337),
.A2(n_6631),
.B(n_6630),
.Y(n_13592)
);

INVx2_ASAP7_75t_SL g13593 ( 
.A(n_13272),
.Y(n_13593)
);

OAI221xp5_ASAP7_75t_L g13594 ( 
.A1(n_13429),
.A2(n_6754),
.B1(n_6871),
.B2(n_6751),
.C(n_6725),
.Y(n_13594)
);

NAND4xp25_ASAP7_75t_L g13595 ( 
.A(n_13451),
.B(n_7023),
.C(n_7104),
.D(n_6768),
.Y(n_13595)
);

INVx1_ASAP7_75t_L g13596 ( 
.A(n_13405),
.Y(n_13596)
);

INVx1_ASAP7_75t_L g13597 ( 
.A(n_13398),
.Y(n_13597)
);

NAND2xp5_ASAP7_75t_L g13598 ( 
.A(n_13400),
.B(n_6499),
.Y(n_13598)
);

NAND2xp5_ASAP7_75t_L g13599 ( 
.A(n_13384),
.B(n_6499),
.Y(n_13599)
);

OR2x2_ASAP7_75t_L g13600 ( 
.A(n_13390),
.B(n_7325),
.Y(n_13600)
);

INVx1_ASAP7_75t_L g13601 ( 
.A(n_13292),
.Y(n_13601)
);

INVx1_ASAP7_75t_L g13602 ( 
.A(n_13370),
.Y(n_13602)
);

INVx2_ASAP7_75t_L g13603 ( 
.A(n_13443),
.Y(n_13603)
);

INVx1_ASAP7_75t_L g13604 ( 
.A(n_13371),
.Y(n_13604)
);

OR2x2_ASAP7_75t_L g13605 ( 
.A(n_13367),
.B(n_7325),
.Y(n_13605)
);

OAI22xp5_ASAP7_75t_SL g13606 ( 
.A1(n_13272),
.A2(n_6025),
.B1(n_6228),
.B2(n_6018),
.Y(n_13606)
);

AOI21xp33_ASAP7_75t_SL g13607 ( 
.A1(n_13444),
.A2(n_7122),
.B(n_6871),
.Y(n_13607)
);

INVx3_ASAP7_75t_L g13608 ( 
.A(n_13382),
.Y(n_13608)
);

OAI21xp5_ASAP7_75t_SL g13609 ( 
.A1(n_13266),
.A2(n_7122),
.B(n_7064),
.Y(n_13609)
);

NAND2xp5_ASAP7_75t_L g13610 ( 
.A(n_13306),
.B(n_6499),
.Y(n_13610)
);

INVx1_ASAP7_75t_SL g13611 ( 
.A(n_13321),
.Y(n_13611)
);

NOR2xp33_ASAP7_75t_L g13612 ( 
.A(n_13459),
.B(n_6626),
.Y(n_13612)
);

A2O1A1Ixp33_ASAP7_75t_L g13613 ( 
.A1(n_13453),
.A2(n_7783),
.B(n_7720),
.C(n_6786),
.Y(n_13613)
);

AO22x1_ASAP7_75t_L g13614 ( 
.A1(n_13410),
.A2(n_6867),
.B1(n_6950),
.B2(n_6850),
.Y(n_13614)
);

O2A1O1Ixp33_ASAP7_75t_L g13615 ( 
.A1(n_13412),
.A2(n_6995),
.B(n_6916),
.C(n_5931),
.Y(n_13615)
);

AND2x2_ASAP7_75t_L g13616 ( 
.A(n_13332),
.B(n_6850),
.Y(n_13616)
);

NAND3xp33_ASAP7_75t_L g13617 ( 
.A(n_13290),
.B(n_6627),
.C(n_6626),
.Y(n_13617)
);

OAI22xp5_ASAP7_75t_SL g13618 ( 
.A1(n_13381),
.A2(n_6025),
.B1(n_6228),
.B2(n_6018),
.Y(n_13618)
);

INVx1_ASAP7_75t_L g13619 ( 
.A(n_13341),
.Y(n_13619)
);

AOI21xp5_ASAP7_75t_L g13620 ( 
.A1(n_13438),
.A2(n_7107),
.B(n_7086),
.Y(n_13620)
);

NAND2xp5_ASAP7_75t_L g13621 ( 
.A(n_13461),
.B(n_6499),
.Y(n_13621)
);

AOI21xp5_ASAP7_75t_L g13622 ( 
.A1(n_13358),
.A2(n_7148),
.B(n_7123),
.Y(n_13622)
);

AOI221xp5_ASAP7_75t_L g13623 ( 
.A1(n_13362),
.A2(n_6682),
.B1(n_6701),
.B2(n_6654),
.C(n_6627),
.Y(n_13623)
);

INVx1_ASAP7_75t_L g13624 ( 
.A(n_13309),
.Y(n_13624)
);

NOR2x1_ASAP7_75t_L g13625 ( 
.A(n_13374),
.B(n_4782),
.Y(n_13625)
);

OAI22xp5_ASAP7_75t_L g13626 ( 
.A1(n_13402),
.A2(n_7148),
.B1(n_7123),
.B2(n_7385),
.Y(n_13626)
);

AND2x2_ASAP7_75t_L g13627 ( 
.A(n_13393),
.B(n_6867),
.Y(n_13627)
);

INVx2_ASAP7_75t_L g13628 ( 
.A(n_13386),
.Y(n_13628)
);

NAND2xp5_ASAP7_75t_L g13629 ( 
.A(n_13401),
.B(n_6627),
.Y(n_13629)
);

INVx1_ASAP7_75t_L g13630 ( 
.A(n_13369),
.Y(n_13630)
);

NAND3xp33_ASAP7_75t_L g13631 ( 
.A(n_13363),
.B(n_6682),
.C(n_6654),
.Y(n_13631)
);

INVx2_ASAP7_75t_SL g13632 ( 
.A(n_13428),
.Y(n_13632)
);

OAI21xp33_ASAP7_75t_L g13633 ( 
.A1(n_13281),
.A2(n_7330),
.B(n_7322),
.Y(n_13633)
);

OAI321xp33_ASAP7_75t_L g13634 ( 
.A1(n_13417),
.A2(n_7034),
.A3(n_6871),
.B1(n_7068),
.B2(n_7012),
.C(n_6754),
.Y(n_13634)
);

INVx1_ASAP7_75t_L g13635 ( 
.A(n_13422),
.Y(n_13635)
);

INVx1_ASAP7_75t_L g13636 ( 
.A(n_13423),
.Y(n_13636)
);

INVx1_ASAP7_75t_L g13637 ( 
.A(n_13425),
.Y(n_13637)
);

OAI21xp5_ASAP7_75t_L g13638 ( 
.A1(n_13349),
.A2(n_6631),
.B(n_6630),
.Y(n_13638)
);

INVx1_ASAP7_75t_L g13639 ( 
.A(n_13447),
.Y(n_13639)
);

O2A1O1Ixp33_ASAP7_75t_L g13640 ( 
.A1(n_13391),
.A2(n_7385),
.B(n_7387),
.C(n_7073),
.Y(n_13640)
);

INVx2_ASAP7_75t_SL g13641 ( 
.A(n_13460),
.Y(n_13641)
);

INVx1_ASAP7_75t_L g13642 ( 
.A(n_13419),
.Y(n_13642)
);

NOR2xp33_ASAP7_75t_L g13643 ( 
.A(n_13449),
.B(n_6654),
.Y(n_13643)
);

INVx1_ASAP7_75t_SL g13644 ( 
.A(n_13445),
.Y(n_13644)
);

O2A1O1Ixp33_ASAP7_75t_L g13645 ( 
.A1(n_13450),
.A2(n_7387),
.B(n_7073),
.C(n_7282),
.Y(n_13645)
);

OAI22x1_ASAP7_75t_L g13646 ( 
.A1(n_13274),
.A2(n_6477),
.B1(n_6490),
.B2(n_6478),
.Y(n_13646)
);

INVx1_ASAP7_75t_L g13647 ( 
.A(n_13456),
.Y(n_13647)
);

INVx2_ASAP7_75t_L g13648 ( 
.A(n_13386),
.Y(n_13648)
);

INVx2_ASAP7_75t_L g13649 ( 
.A(n_13480),
.Y(n_13649)
);

NOR4xp25_ASAP7_75t_L g13650 ( 
.A(n_13476),
.B(n_13302),
.C(n_13458),
.D(n_13434),
.Y(n_13650)
);

INVx2_ASAP7_75t_L g13651 ( 
.A(n_13502),
.Y(n_13651)
);

OAI22xp33_ASAP7_75t_L g13652 ( 
.A1(n_13484),
.A2(n_13414),
.B1(n_13408),
.B2(n_13430),
.Y(n_13652)
);

AND2x2_ASAP7_75t_L g13653 ( 
.A(n_13533),
.B(n_13361),
.Y(n_13653)
);

OAI211xp5_ASAP7_75t_SL g13654 ( 
.A1(n_13469),
.A2(n_13312),
.B(n_13396),
.C(n_13376),
.Y(n_13654)
);

NAND2xp5_ASAP7_75t_L g13655 ( 
.A(n_13593),
.B(n_13329),
.Y(n_13655)
);

HB1xp67_ASAP7_75t_L g13656 ( 
.A(n_13500),
.Y(n_13656)
);

OA21x2_ASAP7_75t_L g13657 ( 
.A1(n_13501),
.A2(n_13346),
.B(n_13293),
.Y(n_13657)
);

AND2x2_ASAP7_75t_SL g13658 ( 
.A(n_13552),
.B(n_13436),
.Y(n_13658)
);

AOI221xp5_ASAP7_75t_L g13659 ( 
.A1(n_13468),
.A2(n_13395),
.B1(n_13331),
.B2(n_13421),
.C(n_13359),
.Y(n_13659)
);

INVx1_ASAP7_75t_L g13660 ( 
.A(n_13483),
.Y(n_13660)
);

INVx1_ASAP7_75t_SL g13661 ( 
.A(n_13481),
.Y(n_13661)
);

NOR2xp33_ASAP7_75t_L g13662 ( 
.A(n_13482),
.B(n_13408),
.Y(n_13662)
);

AOI21xp33_ASAP7_75t_SL g13663 ( 
.A1(n_13487),
.A2(n_13414),
.B(n_13365),
.Y(n_13663)
);

OAI21xp5_ASAP7_75t_L g13664 ( 
.A1(n_13553),
.A2(n_13313),
.B(n_13320),
.Y(n_13664)
);

INVx1_ASAP7_75t_L g13665 ( 
.A(n_13472),
.Y(n_13665)
);

OAI21xp33_ASAP7_75t_L g13666 ( 
.A1(n_13542),
.A2(n_13364),
.B(n_13433),
.Y(n_13666)
);

AOI322xp5_ASAP7_75t_L g13667 ( 
.A1(n_13644),
.A2(n_13455),
.A3(n_13394),
.B1(n_13322),
.B2(n_13421),
.C1(n_13430),
.C2(n_13315),
.Y(n_13667)
);

INVx1_ASAP7_75t_L g13668 ( 
.A(n_13473),
.Y(n_13668)
);

INVx1_ASAP7_75t_L g13669 ( 
.A(n_13560),
.Y(n_13669)
);

NAND2xp5_ASAP7_75t_L g13670 ( 
.A(n_13512),
.B(n_6682),
.Y(n_13670)
);

HB1xp67_ASAP7_75t_L g13671 ( 
.A(n_13540),
.Y(n_13671)
);

OAI21xp5_ASAP7_75t_SL g13672 ( 
.A1(n_13467),
.A2(n_7122),
.B(n_7064),
.Y(n_13672)
);

INVx2_ASAP7_75t_SL g13673 ( 
.A(n_13561),
.Y(n_13673)
);

INVx2_ASAP7_75t_SL g13674 ( 
.A(n_13471),
.Y(n_13674)
);

AOI22xp5_ASAP7_75t_L g13675 ( 
.A1(n_13470),
.A2(n_7034),
.B1(n_7068),
.B2(n_7012),
.Y(n_13675)
);

INVx1_ASAP7_75t_L g13676 ( 
.A(n_13488),
.Y(n_13676)
);

INVx1_ASAP7_75t_L g13677 ( 
.A(n_13525),
.Y(n_13677)
);

INVx1_ASAP7_75t_SL g13678 ( 
.A(n_13563),
.Y(n_13678)
);

NOR2xp33_ASAP7_75t_L g13679 ( 
.A(n_13608),
.B(n_6701),
.Y(n_13679)
);

A2O1A1Ixp33_ASAP7_75t_L g13680 ( 
.A1(n_13478),
.A2(n_8226),
.B(n_8279),
.C(n_8212),
.Y(n_13680)
);

AOI222xp33_ASAP7_75t_L g13681 ( 
.A1(n_13555),
.A2(n_6721),
.B1(n_6713),
.B2(n_6733),
.C1(n_6732),
.C2(n_6701),
.Y(n_13681)
);

INVxp67_ASAP7_75t_L g13682 ( 
.A(n_13466),
.Y(n_13682)
);

INVxp33_ASAP7_75t_L g13683 ( 
.A(n_13497),
.Y(n_13683)
);

INVx1_ASAP7_75t_L g13684 ( 
.A(n_13583),
.Y(n_13684)
);

NAND2xp5_ASAP7_75t_L g13685 ( 
.A(n_13541),
.B(n_6713),
.Y(n_13685)
);

OAI22xp33_ASAP7_75t_L g13686 ( 
.A1(n_13507),
.A2(n_6722),
.B1(n_6738),
.B2(n_6720),
.Y(n_13686)
);

NAND2xp5_ASAP7_75t_L g13687 ( 
.A(n_13608),
.B(n_6713),
.Y(n_13687)
);

AOI32xp33_ASAP7_75t_L g13688 ( 
.A1(n_13490),
.A2(n_6818),
.A3(n_6873),
.B1(n_6872),
.B2(n_8212),
.Y(n_13688)
);

INVx1_ASAP7_75t_L g13689 ( 
.A(n_13565),
.Y(n_13689)
);

INVx1_ASAP7_75t_L g13690 ( 
.A(n_13515),
.Y(n_13690)
);

AOI311xp33_ASAP7_75t_L g13691 ( 
.A1(n_13496),
.A2(n_5593),
.A3(n_5617),
.B(n_5564),
.C(n_5551),
.Y(n_13691)
);

INVx1_ASAP7_75t_L g13692 ( 
.A(n_13554),
.Y(n_13692)
);

NAND2xp5_ASAP7_75t_L g13693 ( 
.A(n_13464),
.B(n_13539),
.Y(n_13693)
);

INVx1_ASAP7_75t_L g13694 ( 
.A(n_13544),
.Y(n_13694)
);

AOI22xp5_ASAP7_75t_L g13695 ( 
.A1(n_13523),
.A2(n_7034),
.B1(n_7068),
.B2(n_7012),
.Y(n_13695)
);

INVx1_ASAP7_75t_L g13696 ( 
.A(n_13550),
.Y(n_13696)
);

AOI21xp5_ASAP7_75t_L g13697 ( 
.A1(n_13477),
.A2(n_7330),
.B(n_7322),
.Y(n_13697)
);

NOR2x1_ASAP7_75t_L g13698 ( 
.A(n_13475),
.B(n_4782),
.Y(n_13698)
);

INVx1_ASAP7_75t_L g13699 ( 
.A(n_13551),
.Y(n_13699)
);

INVx1_ASAP7_75t_L g13700 ( 
.A(n_13566),
.Y(n_13700)
);

INVx1_ASAP7_75t_L g13701 ( 
.A(n_13479),
.Y(n_13701)
);

OAI222xp33_ASAP7_75t_L g13702 ( 
.A1(n_13625),
.A2(n_7128),
.B1(n_7165),
.B2(n_7105),
.C1(n_7122),
.C2(n_7343),
.Y(n_13702)
);

INVx1_ASAP7_75t_SL g13703 ( 
.A(n_13576),
.Y(n_13703)
);

AOI21xp5_ASAP7_75t_L g13704 ( 
.A1(n_13485),
.A2(n_7361),
.B(n_7352),
.Y(n_13704)
);

NAND2xp5_ASAP7_75t_L g13705 ( 
.A(n_13522),
.B(n_6721),
.Y(n_13705)
);

NAND2xp5_ASAP7_75t_L g13706 ( 
.A(n_13530),
.B(n_6721),
.Y(n_13706)
);

OAI22xp5_ASAP7_75t_L g13707 ( 
.A1(n_13520),
.A2(n_5564),
.B1(n_5593),
.B2(n_5551),
.Y(n_13707)
);

OAI211xp5_ASAP7_75t_L g13708 ( 
.A1(n_13489),
.A2(n_5584),
.B(n_5697),
.C(n_5634),
.Y(n_13708)
);

INVx1_ASAP7_75t_L g13709 ( 
.A(n_13577),
.Y(n_13709)
);

INVxp33_ASAP7_75t_L g13710 ( 
.A(n_13531),
.Y(n_13710)
);

OAI221xp5_ASAP7_75t_L g13711 ( 
.A1(n_13609),
.A2(n_7105),
.B1(n_7165),
.B2(n_7128),
.C(n_7064),
.Y(n_13711)
);

INVx1_ASAP7_75t_L g13712 ( 
.A(n_13579),
.Y(n_13712)
);

AOI21xp33_ASAP7_75t_L g13713 ( 
.A1(n_13611),
.A2(n_13505),
.B(n_13630),
.Y(n_13713)
);

NAND2xp5_ASAP7_75t_L g13714 ( 
.A(n_13641),
.B(n_6732),
.Y(n_13714)
);

INVx1_ASAP7_75t_L g13715 ( 
.A(n_13600),
.Y(n_13715)
);

INVx1_ASAP7_75t_L g13716 ( 
.A(n_13558),
.Y(n_13716)
);

AOI221xp5_ASAP7_75t_L g13717 ( 
.A1(n_13474),
.A2(n_6734),
.B1(n_6748),
.B2(n_6733),
.C(n_6732),
.Y(n_13717)
);

INVx2_ASAP7_75t_L g13718 ( 
.A(n_13509),
.Y(n_13718)
);

INVx1_ASAP7_75t_L g13719 ( 
.A(n_13585),
.Y(n_13719)
);

OAI22xp5_ASAP7_75t_L g13720 ( 
.A1(n_13495),
.A2(n_5617),
.B1(n_5633),
.B2(n_5621),
.Y(n_13720)
);

AOI221xp5_ASAP7_75t_L g13721 ( 
.A1(n_13493),
.A2(n_6748),
.B1(n_6749),
.B2(n_6734),
.C(n_6733),
.Y(n_13721)
);

INVxp67_ASAP7_75t_SL g13722 ( 
.A(n_13494),
.Y(n_13722)
);

INVx1_ASAP7_75t_SL g13723 ( 
.A(n_13498),
.Y(n_13723)
);

HB1xp67_ASAP7_75t_L g13724 ( 
.A(n_13499),
.Y(n_13724)
);

AOI211xp5_ASAP7_75t_L g13725 ( 
.A1(n_13486),
.A2(n_7386),
.B(n_7397),
.C(n_7273),
.Y(n_13725)
);

OAI22xp5_ASAP7_75t_L g13726 ( 
.A1(n_13547),
.A2(n_5621),
.B1(n_5644),
.B2(n_5633),
.Y(n_13726)
);

NAND2xp33_ASAP7_75t_SL g13727 ( 
.A(n_13492),
.B(n_5587),
.Y(n_13727)
);

AOI22xp5_ASAP7_75t_L g13728 ( 
.A1(n_13597),
.A2(n_7128),
.B1(n_7165),
.B2(n_7105),
.Y(n_13728)
);

INVxp67_ASAP7_75t_SL g13729 ( 
.A(n_13526),
.Y(n_13729)
);

NAND2x1p5_ASAP7_75t_L g13730 ( 
.A(n_13642),
.B(n_4835),
.Y(n_13730)
);

NAND2xp33_ASAP7_75t_L g13731 ( 
.A(n_13491),
.B(n_5675),
.Y(n_13731)
);

OAI21xp5_ASAP7_75t_L g13732 ( 
.A1(n_13463),
.A2(n_6631),
.B(n_6630),
.Y(n_13732)
);

INVx1_ASAP7_75t_L g13733 ( 
.A(n_13510),
.Y(n_13733)
);

INVx1_ASAP7_75t_L g13734 ( 
.A(n_13514),
.Y(n_13734)
);

INVx1_ASAP7_75t_L g13735 ( 
.A(n_13589),
.Y(n_13735)
);

BUFx2_ASAP7_75t_L g13736 ( 
.A(n_13499),
.Y(n_13736)
);

INVx1_ASAP7_75t_L g13737 ( 
.A(n_13596),
.Y(n_13737)
);

INVx1_ASAP7_75t_L g13738 ( 
.A(n_13586),
.Y(n_13738)
);

INVx1_ASAP7_75t_L g13739 ( 
.A(n_13602),
.Y(n_13739)
);

INVx1_ASAP7_75t_L g13740 ( 
.A(n_13604),
.Y(n_13740)
);

AOI21xp33_ASAP7_75t_SL g13741 ( 
.A1(n_13628),
.A2(n_7361),
.B(n_7352),
.Y(n_13741)
);

HB1xp67_ASAP7_75t_L g13742 ( 
.A(n_13648),
.Y(n_13742)
);

INVx1_ASAP7_75t_L g13743 ( 
.A(n_13590),
.Y(n_13743)
);

AOI32xp33_ASAP7_75t_L g13744 ( 
.A1(n_13521),
.A2(n_6818),
.A3(n_6873),
.B1(n_6872),
.B2(n_8226),
.Y(n_13744)
);

INVx1_ASAP7_75t_L g13745 ( 
.A(n_13598),
.Y(n_13745)
);

OAI21xp5_ASAP7_75t_SL g13746 ( 
.A1(n_13465),
.A2(n_7138),
.B(n_7045),
.Y(n_13746)
);

OAI22xp5_ASAP7_75t_L g13747 ( 
.A1(n_13605),
.A2(n_5644),
.B1(n_5795),
.B2(n_5655),
.Y(n_13747)
);

INVx1_ASAP7_75t_L g13748 ( 
.A(n_13503),
.Y(n_13748)
);

INVx1_ASAP7_75t_SL g13749 ( 
.A(n_13635),
.Y(n_13749)
);

CKINVDCx14_ASAP7_75t_R g13750 ( 
.A(n_13647),
.Y(n_13750)
);

OAI32xp33_ASAP7_75t_L g13751 ( 
.A1(n_13556),
.A2(n_6490),
.A3(n_6614),
.B1(n_6478),
.B2(n_6477),
.Y(n_13751)
);

AOI322xp5_ASAP7_75t_L g13752 ( 
.A1(n_13570),
.A2(n_7172),
.A3(n_6556),
.B1(n_6948),
.B2(n_7056),
.C1(n_7088),
.C2(n_6937),
.Y(n_13752)
);

INVxp67_ASAP7_75t_SL g13753 ( 
.A(n_13569),
.Y(n_13753)
);

OAI222xp33_ASAP7_75t_L g13754 ( 
.A1(n_13603),
.A2(n_7314),
.B1(n_7138),
.B2(n_7377),
.C1(n_7149),
.C2(n_7045),
.Y(n_13754)
);

AOI221xp5_ASAP7_75t_L g13755 ( 
.A1(n_13639),
.A2(n_6749),
.B1(n_6775),
.B2(n_6748),
.C(n_6734),
.Y(n_13755)
);

INVx2_ASAP7_75t_L g13756 ( 
.A(n_13509),
.Y(n_13756)
);

INVx2_ASAP7_75t_L g13757 ( 
.A(n_13636),
.Y(n_13757)
);

AND2x2_ASAP7_75t_L g13758 ( 
.A(n_13532),
.B(n_6867),
.Y(n_13758)
);

AOI22xp33_ASAP7_75t_L g13759 ( 
.A1(n_13619),
.A2(n_6749),
.B1(n_6778),
.B2(n_6775),
.Y(n_13759)
);

AND2x2_ASAP7_75t_L g13760 ( 
.A(n_13557),
.B(n_13559),
.Y(n_13760)
);

INVx1_ASAP7_75t_L g13761 ( 
.A(n_13621),
.Y(n_13761)
);

INVx2_ASAP7_75t_L g13762 ( 
.A(n_13637),
.Y(n_13762)
);

AND2x2_ASAP7_75t_L g13763 ( 
.A(n_13616),
.B(n_13511),
.Y(n_13763)
);

INVx1_ASAP7_75t_L g13764 ( 
.A(n_13610),
.Y(n_13764)
);

INVx1_ASAP7_75t_L g13765 ( 
.A(n_13575),
.Y(n_13765)
);

NAND2xp5_ASAP7_75t_L g13766 ( 
.A(n_13643),
.B(n_6775),
.Y(n_13766)
);

NOR2x1_ASAP7_75t_SL g13767 ( 
.A(n_13632),
.B(n_6401),
.Y(n_13767)
);

OAI22xp5_ASAP7_75t_L g13768 ( 
.A1(n_13548),
.A2(n_5655),
.B1(n_5803),
.B2(n_5795),
.Y(n_13768)
);

OAI32xp33_ASAP7_75t_L g13769 ( 
.A1(n_13562),
.A2(n_6490),
.A3(n_6614),
.B1(n_6478),
.B2(n_6477),
.Y(n_13769)
);

NAND2xp5_ASAP7_75t_L g13770 ( 
.A(n_13582),
.B(n_6778),
.Y(n_13770)
);

AOI21xp5_ASAP7_75t_L g13771 ( 
.A1(n_13587),
.A2(n_7375),
.B(n_7363),
.Y(n_13771)
);

AOI21xp5_ASAP7_75t_L g13772 ( 
.A1(n_13601),
.A2(n_7375),
.B(n_7363),
.Y(n_13772)
);

INVx2_ASAP7_75t_L g13773 ( 
.A(n_13599),
.Y(n_13773)
);

INVxp67_ASAP7_75t_SL g13774 ( 
.A(n_13624),
.Y(n_13774)
);

BUFx3_ASAP7_75t_L g13775 ( 
.A(n_13612),
.Y(n_13775)
);

INVx1_ASAP7_75t_L g13776 ( 
.A(n_13519),
.Y(n_13776)
);

NAND3xp33_ASAP7_75t_L g13777 ( 
.A(n_13536),
.B(n_6781),
.C(n_6778),
.Y(n_13777)
);

NAND2xp5_ASAP7_75t_L g13778 ( 
.A(n_13518),
.B(n_13543),
.Y(n_13778)
);

NAND2xp5_ASAP7_75t_L g13779 ( 
.A(n_13537),
.B(n_6781),
.Y(n_13779)
);

A2O1A1Ixp33_ASAP7_75t_L g13780 ( 
.A1(n_13528),
.A2(n_13529),
.B(n_13506),
.C(n_13629),
.Y(n_13780)
);

INVx2_ASAP7_75t_L g13781 ( 
.A(n_13549),
.Y(n_13781)
);

OAI21xp5_ASAP7_75t_L g13782 ( 
.A1(n_13567),
.A2(n_8279),
.B(n_6730),
.Y(n_13782)
);

INVx1_ASAP7_75t_L g13783 ( 
.A(n_13631),
.Y(n_13783)
);

INVx1_ASAP7_75t_L g13784 ( 
.A(n_13617),
.Y(n_13784)
);

NAND3xp33_ASAP7_75t_L g13785 ( 
.A(n_13591),
.B(n_6821),
.C(n_6781),
.Y(n_13785)
);

INVx1_ASAP7_75t_L g13786 ( 
.A(n_13606),
.Y(n_13786)
);

NOR2xp33_ASAP7_75t_L g13787 ( 
.A(n_13581),
.B(n_6821),
.Y(n_13787)
);

INVx1_ASAP7_75t_L g13788 ( 
.A(n_13535),
.Y(n_13788)
);

OAI32xp33_ASAP7_75t_L g13789 ( 
.A1(n_13594),
.A2(n_6490),
.A3(n_6614),
.B1(n_6478),
.B2(n_6477),
.Y(n_13789)
);

NAND2xp5_ASAP7_75t_L g13790 ( 
.A(n_13627),
.B(n_6821),
.Y(n_13790)
);

NAND2xp5_ASAP7_75t_L g13791 ( 
.A(n_13517),
.B(n_6856),
.Y(n_13791)
);

AOI221xp5_ASAP7_75t_L g13792 ( 
.A1(n_13538),
.A2(n_6889),
.B1(n_6908),
.B2(n_6864),
.C(n_6856),
.Y(n_13792)
);

AOI22xp33_ASAP7_75t_L g13793 ( 
.A1(n_13638),
.A2(n_6856),
.B1(n_6889),
.B2(n_6864),
.Y(n_13793)
);

INVx2_ASAP7_75t_L g13794 ( 
.A(n_13646),
.Y(n_13794)
);

AOI21xp5_ASAP7_75t_L g13795 ( 
.A1(n_13568),
.A2(n_7669),
.B(n_7636),
.Y(n_13795)
);

OR2x2_ASAP7_75t_L g13796 ( 
.A(n_13524),
.B(n_5697),
.Y(n_13796)
);

AOI21xp33_ASAP7_75t_L g13797 ( 
.A1(n_13546),
.A2(n_6889),
.B(n_6864),
.Y(n_13797)
);

NAND2xp5_ASAP7_75t_L g13798 ( 
.A(n_13545),
.B(n_6908),
.Y(n_13798)
);

OAI22xp5_ASAP7_75t_L g13799 ( 
.A1(n_13584),
.A2(n_5803),
.B1(n_5726),
.B2(n_5793),
.Y(n_13799)
);

NAND2xp5_ASAP7_75t_L g13800 ( 
.A(n_13508),
.B(n_6908),
.Y(n_13800)
);

NAND3xp33_ASAP7_75t_L g13801 ( 
.A(n_13504),
.B(n_6952),
.C(n_6910),
.Y(n_13801)
);

AOI221xp5_ASAP7_75t_L g13802 ( 
.A1(n_13607),
.A2(n_6961),
.B1(n_6969),
.B2(n_6952),
.C(n_6910),
.Y(n_13802)
);

OAI211xp5_ASAP7_75t_L g13803 ( 
.A1(n_13588),
.A2(n_13578),
.B(n_13572),
.C(n_13580),
.Y(n_13803)
);

AOI21xp33_ASAP7_75t_SL g13804 ( 
.A1(n_13618),
.A2(n_7138),
.B(n_7045),
.Y(n_13804)
);

INVx1_ASAP7_75t_L g13805 ( 
.A(n_13640),
.Y(n_13805)
);

NOR2xp33_ASAP7_75t_L g13806 ( 
.A(n_13622),
.B(n_6910),
.Y(n_13806)
);

AOI21xp33_ASAP7_75t_L g13807 ( 
.A1(n_13573),
.A2(n_6961),
.B(n_6952),
.Y(n_13807)
);

AOI22xp33_ASAP7_75t_L g13808 ( 
.A1(n_13623),
.A2(n_6961),
.B1(n_6975),
.B2(n_6969),
.Y(n_13808)
);

A2O1A1Ixp33_ASAP7_75t_L g13809 ( 
.A1(n_13534),
.A2(n_6788),
.B(n_6793),
.C(n_6785),
.Y(n_13809)
);

OAI22xp5_ASAP7_75t_L g13810 ( 
.A1(n_13613),
.A2(n_5726),
.B1(n_5793),
.B2(n_5755),
.Y(n_13810)
);

OAI32xp33_ASAP7_75t_L g13811 ( 
.A1(n_13626),
.A2(n_6747),
.A3(n_6711),
.B1(n_6614),
.B2(n_7149),
.Y(n_13811)
);

INVx1_ASAP7_75t_L g13812 ( 
.A(n_13527),
.Y(n_13812)
);

XOR2x2_ASAP7_75t_L g13813 ( 
.A(n_13614),
.B(n_6143),
.Y(n_13813)
);

OAI22xp5_ASAP7_75t_L g13814 ( 
.A1(n_13620),
.A2(n_5755),
.B1(n_6228),
.B2(n_6025),
.Y(n_13814)
);

INVx1_ASAP7_75t_L g13815 ( 
.A(n_13513),
.Y(n_13815)
);

NOR2xp33_ASAP7_75t_L g13816 ( 
.A(n_13683),
.B(n_13633),
.Y(n_13816)
);

NAND2x1p5_ASAP7_75t_L g13817 ( 
.A(n_13678),
.B(n_13634),
.Y(n_13817)
);

AOI221xp5_ASAP7_75t_L g13818 ( 
.A1(n_13736),
.A2(n_13516),
.B1(n_13645),
.B2(n_13592),
.C(n_13574),
.Y(n_13818)
);

AOI22xp33_ASAP7_75t_L g13819 ( 
.A1(n_13773),
.A2(n_13595),
.B1(n_13571),
.B2(n_13564),
.Y(n_13819)
);

CKINVDCx5p33_ASAP7_75t_R g13820 ( 
.A(n_13651),
.Y(n_13820)
);

INVx1_ASAP7_75t_L g13821 ( 
.A(n_13656),
.Y(n_13821)
);

HB1xp67_ASAP7_75t_L g13822 ( 
.A(n_13724),
.Y(n_13822)
);

INVx1_ASAP7_75t_L g13823 ( 
.A(n_13671),
.Y(n_13823)
);

NAND2xp5_ASAP7_75t_L g13824 ( 
.A(n_13658),
.B(n_13615),
.Y(n_13824)
);

INVx1_ASAP7_75t_SL g13825 ( 
.A(n_13661),
.Y(n_13825)
);

INVx3_ASAP7_75t_L g13826 ( 
.A(n_13649),
.Y(n_13826)
);

NAND2xp33_ASAP7_75t_SL g13827 ( 
.A(n_13674),
.B(n_6720),
.Y(n_13827)
);

INVx1_ASAP7_75t_L g13828 ( 
.A(n_13653),
.Y(n_13828)
);

INVx1_ASAP7_75t_L g13829 ( 
.A(n_13673),
.Y(n_13829)
);

INVx1_ASAP7_75t_SL g13830 ( 
.A(n_13703),
.Y(n_13830)
);

INVx1_ASAP7_75t_L g13831 ( 
.A(n_13692),
.Y(n_13831)
);

CKINVDCx16_ASAP7_75t_R g13832 ( 
.A(n_13750),
.Y(n_13832)
);

NAND2xp5_ASAP7_75t_L g13833 ( 
.A(n_13722),
.B(n_13662),
.Y(n_13833)
);

AOI22xp5_ASAP7_75t_L g13834 ( 
.A1(n_13694),
.A2(n_6722),
.B1(n_6738),
.B2(n_6720),
.Y(n_13834)
);

INVx1_ASAP7_75t_SL g13835 ( 
.A(n_13723),
.Y(n_13835)
);

AND2x2_ASAP7_75t_L g13836 ( 
.A(n_13729),
.B(n_6867),
.Y(n_13836)
);

INVx1_ASAP7_75t_L g13837 ( 
.A(n_13742),
.Y(n_13837)
);

AND2x2_ASAP7_75t_L g13838 ( 
.A(n_13665),
.B(n_13710),
.Y(n_13838)
);

NAND2xp5_ASAP7_75t_L g13839 ( 
.A(n_13699),
.B(n_6969),
.Y(n_13839)
);

INVx1_ASAP7_75t_SL g13840 ( 
.A(n_13655),
.Y(n_13840)
);

INVx1_ASAP7_75t_L g13841 ( 
.A(n_13669),
.Y(n_13841)
);

INVx1_ASAP7_75t_L g13842 ( 
.A(n_13657),
.Y(n_13842)
);

AND2x2_ASAP7_75t_L g13843 ( 
.A(n_13660),
.B(n_6867),
.Y(n_13843)
);

NOR2xp33_ASAP7_75t_SL g13844 ( 
.A(n_13684),
.B(n_4842),
.Y(n_13844)
);

AND2x2_ASAP7_75t_L g13845 ( 
.A(n_13760),
.B(n_13715),
.Y(n_13845)
);

NAND2xp5_ASAP7_75t_L g13846 ( 
.A(n_13774),
.B(n_6975),
.Y(n_13846)
);

AND2x2_ASAP7_75t_L g13847 ( 
.A(n_13719),
.B(n_13698),
.Y(n_13847)
);

NAND2xp5_ASAP7_75t_L g13848 ( 
.A(n_13749),
.B(n_6975),
.Y(n_13848)
);

OR2x2_ASAP7_75t_L g13849 ( 
.A(n_13730),
.B(n_7283),
.Y(n_13849)
);

HB1xp67_ASAP7_75t_L g13850 ( 
.A(n_13657),
.Y(n_13850)
);

AOI221x1_ASAP7_75t_SL g13851 ( 
.A1(n_13652),
.A2(n_7136),
.B1(n_7104),
.B2(n_6768),
.C(n_6966),
.Y(n_13851)
);

AND2x2_ASAP7_75t_L g13852 ( 
.A(n_13682),
.B(n_6950),
.Y(n_13852)
);

INVx1_ASAP7_75t_L g13853 ( 
.A(n_13753),
.Y(n_13853)
);

INVx1_ASAP7_75t_SL g13854 ( 
.A(n_13709),
.Y(n_13854)
);

INVx1_ASAP7_75t_L g13855 ( 
.A(n_13712),
.Y(n_13855)
);

INVx1_ASAP7_75t_L g13856 ( 
.A(n_13690),
.Y(n_13856)
);

AND2x2_ASAP7_75t_L g13857 ( 
.A(n_13668),
.B(n_6950),
.Y(n_13857)
);

NOR2xp33_ASAP7_75t_L g13858 ( 
.A(n_13654),
.B(n_7081),
.Y(n_13858)
);

AND2x2_ASAP7_75t_L g13859 ( 
.A(n_13701),
.B(n_6950),
.Y(n_13859)
);

AND2x2_ASAP7_75t_L g13860 ( 
.A(n_13758),
.B(n_6950),
.Y(n_13860)
);

INVxp67_ASAP7_75t_L g13861 ( 
.A(n_13775),
.Y(n_13861)
);

INVx1_ASAP7_75t_L g13862 ( 
.A(n_13689),
.Y(n_13862)
);

INVx2_ASAP7_75t_L g13863 ( 
.A(n_13757),
.Y(n_13863)
);

NAND2xp5_ASAP7_75t_L g13864 ( 
.A(n_13667),
.B(n_6982),
.Y(n_13864)
);

INVx1_ASAP7_75t_L g13865 ( 
.A(n_13696),
.Y(n_13865)
);

INVx1_ASAP7_75t_SL g13866 ( 
.A(n_13693),
.Y(n_13866)
);

INVx1_ASAP7_75t_SL g13867 ( 
.A(n_13700),
.Y(n_13867)
);

NAND2xp5_ASAP7_75t_L g13868 ( 
.A(n_13781),
.B(n_6982),
.Y(n_13868)
);

OR2x2_ASAP7_75t_L g13869 ( 
.A(n_13716),
.B(n_13650),
.Y(n_13869)
);

INVx1_ASAP7_75t_L g13870 ( 
.A(n_13734),
.Y(n_13870)
);

INVxp67_ASAP7_75t_L g13871 ( 
.A(n_13776),
.Y(n_13871)
);

NOR2xp33_ASAP7_75t_L g13872 ( 
.A(n_13713),
.B(n_7144),
.Y(n_13872)
);

INVx1_ASAP7_75t_L g13873 ( 
.A(n_13735),
.Y(n_13873)
);

INVx1_ASAP7_75t_L g13874 ( 
.A(n_13737),
.Y(n_13874)
);

HB1xp67_ASAP7_75t_L g13875 ( 
.A(n_13762),
.Y(n_13875)
);

AOI22xp33_ASAP7_75t_SL g13876 ( 
.A1(n_13676),
.A2(n_6722),
.B1(n_6738),
.B2(n_6720),
.Y(n_13876)
);

INVx1_ASAP7_75t_L g13877 ( 
.A(n_13677),
.Y(n_13877)
);

NAND2xp33_ASAP7_75t_L g13878 ( 
.A(n_13666),
.B(n_6722),
.Y(n_13878)
);

INVx1_ASAP7_75t_L g13879 ( 
.A(n_13739),
.Y(n_13879)
);

INVx1_ASAP7_75t_L g13880 ( 
.A(n_13740),
.Y(n_13880)
);

NOR2xp33_ASAP7_75t_L g13881 ( 
.A(n_13718),
.B(n_7090),
.Y(n_13881)
);

NAND2xp5_ASAP7_75t_L g13882 ( 
.A(n_13788),
.B(n_6982),
.Y(n_13882)
);

NAND2xp5_ASAP7_75t_L g13883 ( 
.A(n_13679),
.B(n_6990),
.Y(n_13883)
);

INVx1_ASAP7_75t_L g13884 ( 
.A(n_13687),
.Y(n_13884)
);

NAND2xp5_ASAP7_75t_L g13885 ( 
.A(n_13756),
.B(n_6990),
.Y(n_13885)
);

INVx2_ASAP7_75t_L g13886 ( 
.A(n_13767),
.Y(n_13886)
);

AND2x2_ASAP7_75t_L g13887 ( 
.A(n_13763),
.B(n_6966),
.Y(n_13887)
);

NOR2xp33_ASAP7_75t_L g13888 ( 
.A(n_13733),
.B(n_7151),
.Y(n_13888)
);

INVx2_ASAP7_75t_L g13889 ( 
.A(n_13794),
.Y(n_13889)
);

AND2x2_ASAP7_75t_L g13890 ( 
.A(n_13691),
.B(n_13664),
.Y(n_13890)
);

NAND2xp5_ASAP7_75t_L g13891 ( 
.A(n_13784),
.B(n_6990),
.Y(n_13891)
);

INVx2_ASAP7_75t_L g13892 ( 
.A(n_13685),
.Y(n_13892)
);

INVx1_ASAP7_75t_L g13893 ( 
.A(n_13670),
.Y(n_13893)
);

INVx2_ASAP7_75t_L g13894 ( 
.A(n_13714),
.Y(n_13894)
);

AND2x2_ASAP7_75t_L g13895 ( 
.A(n_13786),
.B(n_6966),
.Y(n_13895)
);

INVx2_ASAP7_75t_L g13896 ( 
.A(n_13743),
.Y(n_13896)
);

OR2x2_ASAP7_75t_L g13897 ( 
.A(n_13778),
.B(n_7283),
.Y(n_13897)
);

NAND2x1p5_ASAP7_75t_L g13898 ( 
.A(n_13745),
.B(n_4842),
.Y(n_13898)
);

NAND2xp5_ASAP7_75t_L g13899 ( 
.A(n_13783),
.B(n_6994),
.Y(n_13899)
);

NAND2x1_ASAP7_75t_L g13900 ( 
.A(n_13812),
.B(n_7228),
.Y(n_13900)
);

NOR2xp33_ASAP7_75t_L g13901 ( 
.A(n_13738),
.B(n_7187),
.Y(n_13901)
);

INVx1_ASAP7_75t_L g13902 ( 
.A(n_13705),
.Y(n_13902)
);

NAND2xp5_ASAP7_75t_L g13903 ( 
.A(n_13764),
.B(n_6994),
.Y(n_13903)
);

AND2x2_ASAP7_75t_L g13904 ( 
.A(n_13805),
.B(n_13663),
.Y(n_13904)
);

AND2x2_ASAP7_75t_L g13905 ( 
.A(n_13813),
.B(n_6966),
.Y(n_13905)
);

INVx2_ASAP7_75t_L g13906 ( 
.A(n_13815),
.Y(n_13906)
);

NAND2xp5_ASAP7_75t_L g13907 ( 
.A(n_13761),
.B(n_6994),
.Y(n_13907)
);

NAND3xp33_ASAP7_75t_L g13908 ( 
.A(n_13748),
.B(n_7048),
.C(n_7040),
.Y(n_13908)
);

AND2x4_ASAP7_75t_SL g13909 ( 
.A(n_13765),
.B(n_7127),
.Y(n_13909)
);

HB1xp67_ASAP7_75t_L g13910 ( 
.A(n_13659),
.Y(n_13910)
);

OR2x2_ASAP7_75t_L g13911 ( 
.A(n_13790),
.B(n_7283),
.Y(n_13911)
);

NAND2xp5_ASAP7_75t_L g13912 ( 
.A(n_13806),
.B(n_13780),
.Y(n_13912)
);

INVx1_ASAP7_75t_L g13913 ( 
.A(n_13731),
.Y(n_13913)
);

INVx1_ASAP7_75t_L g13914 ( 
.A(n_13727),
.Y(n_13914)
);

NOR2xp33_ASAP7_75t_L g13915 ( 
.A(n_13791),
.B(n_7118),
.Y(n_13915)
);

INVx1_ASAP7_75t_L g13916 ( 
.A(n_13706),
.Y(n_13916)
);

HB1xp67_ASAP7_75t_L g13917 ( 
.A(n_13720),
.Y(n_13917)
);

NAND2xp5_ASAP7_75t_L g13918 ( 
.A(n_13766),
.B(n_7040),
.Y(n_13918)
);

INVx1_ASAP7_75t_SL g13919 ( 
.A(n_13796),
.Y(n_13919)
);

NOR3xp33_ASAP7_75t_L g13920 ( 
.A(n_13803),
.B(n_4842),
.C(n_6668),
.Y(n_13920)
);

NAND2xp5_ASAP7_75t_L g13921 ( 
.A(n_13770),
.B(n_7040),
.Y(n_13921)
);

BUFx2_ASAP7_75t_L g13922 ( 
.A(n_13779),
.Y(n_13922)
);

NAND2xp33_ASAP7_75t_L g13923 ( 
.A(n_13680),
.B(n_13688),
.Y(n_13923)
);

INVx1_ASAP7_75t_L g13924 ( 
.A(n_13800),
.Y(n_13924)
);

INVx2_ASAP7_75t_SL g13925 ( 
.A(n_13798),
.Y(n_13925)
);

INVx1_ASAP7_75t_L g13926 ( 
.A(n_13785),
.Y(n_13926)
);

AND2x2_ASAP7_75t_L g13927 ( 
.A(n_13741),
.B(n_6966),
.Y(n_13927)
);

NOR2xp33_ASAP7_75t_SL g13928 ( 
.A(n_13702),
.B(n_7127),
.Y(n_13928)
);

AND2x2_ASAP7_75t_L g13929 ( 
.A(n_13697),
.B(n_7032),
.Y(n_13929)
);

OAI22xp5_ASAP7_75t_L g13930 ( 
.A1(n_13695),
.A2(n_13728),
.B1(n_13809),
.B2(n_13810),
.Y(n_13930)
);

AND2x2_ASAP7_75t_L g13931 ( 
.A(n_13772),
.B(n_7032),
.Y(n_13931)
);

INVx1_ASAP7_75t_L g13932 ( 
.A(n_13787),
.Y(n_13932)
);

INVxp67_ASAP7_75t_SL g13933 ( 
.A(n_13686),
.Y(n_13933)
);

NAND2xp5_ASAP7_75t_L g13934 ( 
.A(n_13704),
.B(n_13777),
.Y(n_13934)
);

INVx1_ASAP7_75t_L g13935 ( 
.A(n_13708),
.Y(n_13935)
);

INVx2_ASAP7_75t_L g13936 ( 
.A(n_13801),
.Y(n_13936)
);

AOI22xp33_ASAP7_75t_L g13937 ( 
.A1(n_13807),
.A2(n_7048),
.B1(n_7081),
.B2(n_7074),
.Y(n_13937)
);

INVx1_ASAP7_75t_SL g13938 ( 
.A(n_13771),
.Y(n_13938)
);

NAND2xp5_ASAP7_75t_L g13939 ( 
.A(n_13768),
.B(n_7048),
.Y(n_13939)
);

INVx1_ASAP7_75t_SL g13940 ( 
.A(n_13675),
.Y(n_13940)
);

INVx1_ASAP7_75t_SL g13941 ( 
.A(n_13799),
.Y(n_13941)
);

NAND2xp5_ASAP7_75t_L g13942 ( 
.A(n_13746),
.B(n_7074),
.Y(n_13942)
);

OAI22xp5_ASAP7_75t_L g13943 ( 
.A1(n_13795),
.A2(n_6228),
.B1(n_6428),
.B2(n_6025),
.Y(n_13943)
);

AND2x2_ASAP7_75t_SL g13944 ( 
.A(n_13759),
.B(n_6738),
.Y(n_13944)
);

NOR2xp33_ASAP7_75t_L g13945 ( 
.A(n_13751),
.B(n_7256),
.Y(n_13945)
);

OR2x2_ASAP7_75t_L g13946 ( 
.A(n_13814),
.B(n_7283),
.Y(n_13946)
);

INVx2_ASAP7_75t_L g13947 ( 
.A(n_13726),
.Y(n_13947)
);

OR2x2_ASAP7_75t_L g13948 ( 
.A(n_13747),
.B(n_7283),
.Y(n_13948)
);

NOR2xp33_ASAP7_75t_L g13949 ( 
.A(n_13769),
.B(n_7256),
.Y(n_13949)
);

INVxp67_ASAP7_75t_L g13950 ( 
.A(n_13804),
.Y(n_13950)
);

NOR2xp33_ASAP7_75t_L g13951 ( 
.A(n_13732),
.B(n_7256),
.Y(n_13951)
);

OAI221xp5_ASAP7_75t_L g13952 ( 
.A1(n_13782),
.A2(n_7149),
.B1(n_7377),
.B2(n_7314),
.C(n_6747),
.Y(n_13952)
);

INVx2_ASAP7_75t_L g13953 ( 
.A(n_13707),
.Y(n_13953)
);

NOR3xp33_ASAP7_75t_L g13954 ( 
.A(n_13672),
.B(n_6668),
.C(n_6853),
.Y(n_13954)
);

NAND2xp5_ASAP7_75t_L g13955 ( 
.A(n_13717),
.B(n_13681),
.Y(n_13955)
);

NOR2xp33_ASAP7_75t_L g13956 ( 
.A(n_13797),
.B(n_7090),
.Y(n_13956)
);

AND2x2_ASAP7_75t_L g13957 ( 
.A(n_13725),
.B(n_13752),
.Y(n_13957)
);

AOI22xp33_ASAP7_75t_L g13958 ( 
.A1(n_13721),
.A2(n_7399),
.B1(n_7081),
.B2(n_7090),
.Y(n_13958)
);

AOI221x1_ASAP7_75t_SL g13959 ( 
.A1(n_13744),
.A2(n_7136),
.B1(n_7050),
.B2(n_7094),
.C(n_7047),
.Y(n_13959)
);

OR2x2_ASAP7_75t_L g13960 ( 
.A(n_13793),
.B(n_13711),
.Y(n_13960)
);

NAND2x1_ASAP7_75t_L g13961 ( 
.A(n_13808),
.B(n_7228),
.Y(n_13961)
);

NAND2xp5_ASAP7_75t_L g13962 ( 
.A(n_13755),
.B(n_7074),
.Y(n_13962)
);

NAND2xp33_ASAP7_75t_L g13963 ( 
.A(n_13789),
.B(n_6738),
.Y(n_13963)
);

INVxp67_ASAP7_75t_L g13964 ( 
.A(n_13802),
.Y(n_13964)
);

INVx1_ASAP7_75t_L g13965 ( 
.A(n_13811),
.Y(n_13965)
);

INVx1_ASAP7_75t_L g13966 ( 
.A(n_13792),
.Y(n_13966)
);

AND2x2_ASAP7_75t_L g13967 ( 
.A(n_13754),
.B(n_7032),
.Y(n_13967)
);

INVx1_ASAP7_75t_L g13968 ( 
.A(n_13656),
.Y(n_13968)
);

INVx1_ASAP7_75t_SL g13969 ( 
.A(n_13678),
.Y(n_13969)
);

OAI221xp5_ASAP7_75t_L g13970 ( 
.A1(n_13736),
.A2(n_7314),
.B1(n_7377),
.B2(n_6747),
.C(n_6711),
.Y(n_13970)
);

INVx2_ASAP7_75t_L g13971 ( 
.A(n_13651),
.Y(n_13971)
);

INVx1_ASAP7_75t_SL g13972 ( 
.A(n_13678),
.Y(n_13972)
);

NAND2xp33_ASAP7_75t_L g13973 ( 
.A(n_13678),
.B(n_6738),
.Y(n_13973)
);

NAND2xp5_ASAP7_75t_L g13974 ( 
.A(n_13736),
.B(n_7101),
.Y(n_13974)
);

NAND2xp5_ASAP7_75t_L g13975 ( 
.A(n_13736),
.B(n_7101),
.Y(n_13975)
);

NAND2xp5_ASAP7_75t_L g13976 ( 
.A(n_13736),
.B(n_7101),
.Y(n_13976)
);

OAI21xp5_ASAP7_75t_L g13977 ( 
.A1(n_13683),
.A2(n_6793),
.B(n_6788),
.Y(n_13977)
);

NAND2xp33_ASAP7_75t_L g13978 ( 
.A(n_13678),
.B(n_6814),
.Y(n_13978)
);

AND2x2_ASAP7_75t_L g13979 ( 
.A(n_13658),
.B(n_7032),
.Y(n_13979)
);

INVx2_ASAP7_75t_SL g13980 ( 
.A(n_13651),
.Y(n_13980)
);

NAND2xp5_ASAP7_75t_L g13981 ( 
.A(n_13736),
.B(n_7118),
.Y(n_13981)
);

INVx1_ASAP7_75t_L g13982 ( 
.A(n_13736),
.Y(n_13982)
);

OR2x2_ASAP7_75t_L g13983 ( 
.A(n_13832),
.B(n_6556),
.Y(n_13983)
);

HB1xp67_ASAP7_75t_L g13984 ( 
.A(n_13850),
.Y(n_13984)
);

AND2x2_ASAP7_75t_L g13985 ( 
.A(n_13825),
.B(n_7032),
.Y(n_13985)
);

NAND2xp5_ASAP7_75t_L g13986 ( 
.A(n_13822),
.B(n_7118),
.Y(n_13986)
);

INVxp67_ASAP7_75t_L g13987 ( 
.A(n_13875),
.Y(n_13987)
);

NAND2xp5_ASAP7_75t_L g13988 ( 
.A(n_13826),
.B(n_7121),
.Y(n_13988)
);

CKINVDCx5p33_ASAP7_75t_R g13989 ( 
.A(n_13820),
.Y(n_13989)
);

INVx1_ASAP7_75t_L g13990 ( 
.A(n_13845),
.Y(n_13990)
);

OR2x2_ASAP7_75t_L g13991 ( 
.A(n_13969),
.B(n_6556),
.Y(n_13991)
);

INVx1_ASAP7_75t_L g13992 ( 
.A(n_13837),
.Y(n_13992)
);

NOR3xp33_ASAP7_75t_SL g13993 ( 
.A(n_13833),
.B(n_13842),
.C(n_13982),
.Y(n_13993)
);

AND2x2_ASAP7_75t_L g13994 ( 
.A(n_13972),
.B(n_7108),
.Y(n_13994)
);

INVxp67_ASAP7_75t_L g13995 ( 
.A(n_13853),
.Y(n_13995)
);

OAI22xp5_ASAP7_75t_L g13996 ( 
.A1(n_13835),
.A2(n_6228),
.B1(n_6428),
.B2(n_6025),
.Y(n_13996)
);

AND2x2_ASAP7_75t_L g13997 ( 
.A(n_13826),
.B(n_13830),
.Y(n_13997)
);

NAND3xp33_ASAP7_75t_L g13998 ( 
.A(n_13982),
.B(n_7140),
.C(n_7121),
.Y(n_13998)
);

INVx1_ASAP7_75t_L g13999 ( 
.A(n_13869),
.Y(n_13999)
);

INVx2_ASAP7_75t_L g14000 ( 
.A(n_13980),
.Y(n_14000)
);

NAND2xp5_ASAP7_75t_L g14001 ( 
.A(n_13866),
.B(n_7121),
.Y(n_14001)
);

NAND2xp5_ASAP7_75t_L g14002 ( 
.A(n_13840),
.B(n_7140),
.Y(n_14002)
);

NAND3xp33_ASAP7_75t_L g14003 ( 
.A(n_13823),
.B(n_7144),
.C(n_7140),
.Y(n_14003)
);

AND2x2_ASAP7_75t_L g14004 ( 
.A(n_13979),
.B(n_7108),
.Y(n_14004)
);

INVx1_ASAP7_75t_SL g14005 ( 
.A(n_13854),
.Y(n_14005)
);

NAND3xp33_ASAP7_75t_SL g14006 ( 
.A(n_13867),
.B(n_7151),
.C(n_7144),
.Y(n_14006)
);

OAI21xp33_ASAP7_75t_L g14007 ( 
.A1(n_13828),
.A2(n_7050),
.B(n_7047),
.Y(n_14007)
);

NAND2x1p5_ASAP7_75t_L g14008 ( 
.A(n_13821),
.B(n_6814),
.Y(n_14008)
);

NAND2xp5_ASAP7_75t_L g14009 ( 
.A(n_13968),
.B(n_7151),
.Y(n_14009)
);

INVx1_ASAP7_75t_L g14010 ( 
.A(n_13838),
.Y(n_14010)
);

NOR2x1_ASAP7_75t_L g14011 ( 
.A(n_13831),
.B(n_6158),
.Y(n_14011)
);

NAND2xp5_ASAP7_75t_L g14012 ( 
.A(n_13971),
.B(n_7171),
.Y(n_14012)
);

AND2x2_ASAP7_75t_L g14013 ( 
.A(n_13836),
.B(n_7365),
.Y(n_14013)
);

OA21x2_ASAP7_75t_SL g14014 ( 
.A1(n_13827),
.A2(n_7050),
.B(n_7047),
.Y(n_14014)
);

INVx1_ASAP7_75t_L g14015 ( 
.A(n_13863),
.Y(n_14015)
);

AND2x2_ASAP7_75t_L g14016 ( 
.A(n_13887),
.B(n_7365),
.Y(n_14016)
);

OR2x2_ASAP7_75t_L g14017 ( 
.A(n_13889),
.B(n_13817),
.Y(n_14017)
);

NAND2xp5_ASAP7_75t_L g14018 ( 
.A(n_13904),
.B(n_7171),
.Y(n_14018)
);

INVxp67_ASAP7_75t_L g14019 ( 
.A(n_13910),
.Y(n_14019)
);

AND2x2_ASAP7_75t_L g14020 ( 
.A(n_13857),
.B(n_7365),
.Y(n_14020)
);

NOR3xp33_ASAP7_75t_SL g14021 ( 
.A(n_13912),
.B(n_6366),
.C(n_6243),
.Y(n_14021)
);

INVx1_ASAP7_75t_L g14022 ( 
.A(n_13847),
.Y(n_14022)
);

INVx1_ASAP7_75t_L g14023 ( 
.A(n_13879),
.Y(n_14023)
);

OR2x2_ASAP7_75t_L g14024 ( 
.A(n_13871),
.B(n_6556),
.Y(n_14024)
);

INVx1_ASAP7_75t_L g14025 ( 
.A(n_13880),
.Y(n_14025)
);

AND2x2_ASAP7_75t_L g14026 ( 
.A(n_13859),
.B(n_7365),
.Y(n_14026)
);

INVx1_ASAP7_75t_L g14027 ( 
.A(n_13870),
.Y(n_14027)
);

NAND2xp5_ASAP7_75t_L g14028 ( 
.A(n_13886),
.B(n_7171),
.Y(n_14028)
);

HB1xp67_ASAP7_75t_L g14029 ( 
.A(n_13861),
.Y(n_14029)
);

INVx1_ASAP7_75t_L g14030 ( 
.A(n_13873),
.Y(n_14030)
);

NAND3xp33_ASAP7_75t_L g14031 ( 
.A(n_13841),
.B(n_7187),
.C(n_7185),
.Y(n_14031)
);

XNOR2xp5_ASAP7_75t_L g14032 ( 
.A(n_13890),
.B(n_6143),
.Y(n_14032)
);

INVx1_ASAP7_75t_L g14033 ( 
.A(n_13874),
.Y(n_14033)
);

INVx1_ASAP7_75t_L g14034 ( 
.A(n_13877),
.Y(n_14034)
);

XOR2xp5_ASAP7_75t_L g14035 ( 
.A(n_13829),
.B(n_6896),
.Y(n_14035)
);

OAI21xp5_ASAP7_75t_L g14036 ( 
.A1(n_13855),
.A2(n_6761),
.B(n_7887),
.Y(n_14036)
);

NOR3xp33_ASAP7_75t_L g14037 ( 
.A(n_13856),
.B(n_6869),
.C(n_6853),
.Y(n_14037)
);

INVx1_ASAP7_75t_SL g14038 ( 
.A(n_13862),
.Y(n_14038)
);

BUFx2_ASAP7_75t_L g14039 ( 
.A(n_13906),
.Y(n_14039)
);

AND2x2_ASAP7_75t_L g14040 ( 
.A(n_13860),
.B(n_7047),
.Y(n_14040)
);

INVx1_ASAP7_75t_L g14041 ( 
.A(n_13865),
.Y(n_14041)
);

INVx1_ASAP7_75t_L g14042 ( 
.A(n_13824),
.Y(n_14042)
);

AND2x4_ASAP7_75t_SL g14043 ( 
.A(n_13852),
.B(n_13895),
.Y(n_14043)
);

CKINVDCx8_ASAP7_75t_R g14044 ( 
.A(n_13922),
.Y(n_14044)
);

AND2x2_ASAP7_75t_L g14045 ( 
.A(n_13927),
.B(n_7047),
.Y(n_14045)
);

NOR2xp33_ASAP7_75t_L g14046 ( 
.A(n_13919),
.B(n_7185),
.Y(n_14046)
);

NAND2xp5_ASAP7_75t_L g14047 ( 
.A(n_13858),
.B(n_7187),
.Y(n_14047)
);

AOI221xp5_ASAP7_75t_L g14048 ( 
.A1(n_13950),
.A2(n_7233),
.B1(n_7247),
.B2(n_7200),
.C(n_7185),
.Y(n_14048)
);

INVx1_ASAP7_75t_L g14049 ( 
.A(n_13974),
.Y(n_14049)
);

O2A1O1Ixp33_ASAP7_75t_L g14050 ( 
.A1(n_13914),
.A2(n_7282),
.B(n_7248),
.C(n_6747),
.Y(n_14050)
);

INVx1_ASAP7_75t_L g14051 ( 
.A(n_13975),
.Y(n_14051)
);

INVx1_ASAP7_75t_L g14052 ( 
.A(n_13976),
.Y(n_14052)
);

BUFx3_ASAP7_75t_L g14053 ( 
.A(n_13896),
.Y(n_14053)
);

NAND2xp5_ASAP7_75t_L g14054 ( 
.A(n_13892),
.B(n_7247),
.Y(n_14054)
);

NAND2xp5_ASAP7_75t_L g14055 ( 
.A(n_13894),
.B(n_7247),
.Y(n_14055)
);

INVx1_ASAP7_75t_L g14056 ( 
.A(n_13981),
.Y(n_14056)
);

CKINVDCx5p33_ASAP7_75t_R g14057 ( 
.A(n_13816),
.Y(n_14057)
);

INVx2_ASAP7_75t_L g14058 ( 
.A(n_13898),
.Y(n_14058)
);

BUFx2_ASAP7_75t_L g14059 ( 
.A(n_13933),
.Y(n_14059)
);

INVx1_ASAP7_75t_L g14060 ( 
.A(n_13846),
.Y(n_14060)
);

AOI211xp5_ASAP7_75t_L g14061 ( 
.A1(n_13935),
.A2(n_6814),
.B(n_7038),
.C(n_6919),
.Y(n_14061)
);

INVx1_ASAP7_75t_SL g14062 ( 
.A(n_13938),
.Y(n_14062)
);

OR2x2_ASAP7_75t_L g14063 ( 
.A(n_13864),
.B(n_6556),
.Y(n_14063)
);

INVx1_ASAP7_75t_L g14064 ( 
.A(n_13848),
.Y(n_14064)
);

NOR2xp33_ASAP7_75t_L g14065 ( 
.A(n_13926),
.B(n_7200),
.Y(n_14065)
);

AND2x2_ASAP7_75t_L g14066 ( 
.A(n_13967),
.B(n_7050),
.Y(n_14066)
);

INVx1_ASAP7_75t_L g14067 ( 
.A(n_13843),
.Y(n_14067)
);

HB1xp67_ASAP7_75t_L g14068 ( 
.A(n_13917),
.Y(n_14068)
);

AOI21xp5_ASAP7_75t_L g14069 ( 
.A1(n_13923),
.A2(n_7898),
.B(n_7887),
.Y(n_14069)
);

INVx1_ASAP7_75t_SL g14070 ( 
.A(n_13940),
.Y(n_14070)
);

AND2x2_ASAP7_75t_L g14071 ( 
.A(n_13931),
.B(n_7050),
.Y(n_14071)
);

INVx1_ASAP7_75t_L g14072 ( 
.A(n_13839),
.Y(n_14072)
);

AND2x2_ASAP7_75t_L g14073 ( 
.A(n_13929),
.B(n_7177),
.Y(n_14073)
);

OAI31xp33_ASAP7_75t_L g14074 ( 
.A1(n_13872),
.A2(n_7314),
.A3(n_7377),
.B(n_6711),
.Y(n_14074)
);

INVx1_ASAP7_75t_L g14075 ( 
.A(n_13868),
.Y(n_14075)
);

NOR2xp33_ASAP7_75t_L g14076 ( 
.A(n_13844),
.B(n_7200),
.Y(n_14076)
);

AND2x2_ASAP7_75t_L g14077 ( 
.A(n_13909),
.B(n_7177),
.Y(n_14077)
);

INVx1_ASAP7_75t_L g14078 ( 
.A(n_13882),
.Y(n_14078)
);

INVx2_ASAP7_75t_L g14079 ( 
.A(n_13944),
.Y(n_14079)
);

NOR2xp33_ASAP7_75t_L g14080 ( 
.A(n_13897),
.B(n_7233),
.Y(n_14080)
);

INVx1_ASAP7_75t_L g14081 ( 
.A(n_13888),
.Y(n_14081)
);

AND2x2_ASAP7_75t_L g14082 ( 
.A(n_13905),
.B(n_13913),
.Y(n_14082)
);

NOR3xp33_ASAP7_75t_SL g14083 ( 
.A(n_13893),
.B(n_6366),
.C(n_6243),
.Y(n_14083)
);

OR2x2_ASAP7_75t_L g14084 ( 
.A(n_13934),
.B(n_6556),
.Y(n_14084)
);

OR2x2_ASAP7_75t_L g14085 ( 
.A(n_13925),
.B(n_6556),
.Y(n_14085)
);

INVx1_ASAP7_75t_L g14086 ( 
.A(n_13902),
.Y(n_14086)
);

XNOR2xp5_ASAP7_75t_L g14087 ( 
.A(n_13818),
.B(n_7112),
.Y(n_14087)
);

INVx2_ASAP7_75t_L g14088 ( 
.A(n_13849),
.Y(n_14088)
);

INVx1_ASAP7_75t_L g14089 ( 
.A(n_13891),
.Y(n_14089)
);

INVx1_ASAP7_75t_L g14090 ( 
.A(n_13899),
.Y(n_14090)
);

HB1xp67_ASAP7_75t_L g14091 ( 
.A(n_13884),
.Y(n_14091)
);

AND2x2_ASAP7_75t_L g14092 ( 
.A(n_13965),
.B(n_7108),
.Y(n_14092)
);

INVx1_ASAP7_75t_L g14093 ( 
.A(n_13903),
.Y(n_14093)
);

AOI21xp5_ASAP7_75t_L g14094 ( 
.A1(n_13955),
.A2(n_7906),
.B(n_7898),
.Y(n_14094)
);

HB1xp67_ASAP7_75t_L g14095 ( 
.A(n_13924),
.Y(n_14095)
);

NAND2xp5_ASAP7_75t_L g14096 ( 
.A(n_13915),
.B(n_7233),
.Y(n_14096)
);

NAND2xp5_ASAP7_75t_L g14097 ( 
.A(n_13916),
.B(n_7259),
.Y(n_14097)
);

INVx1_ASAP7_75t_L g14098 ( 
.A(n_13907),
.Y(n_14098)
);

INVx1_ASAP7_75t_L g14099 ( 
.A(n_13885),
.Y(n_14099)
);

OAI221xp5_ASAP7_75t_L g14100 ( 
.A1(n_13920),
.A2(n_6711),
.B1(n_6814),
.B2(n_7038),
.C(n_6919),
.Y(n_14100)
);

INVxp67_ASAP7_75t_L g14101 ( 
.A(n_13932),
.Y(n_14101)
);

INVx2_ASAP7_75t_L g14102 ( 
.A(n_13911),
.Y(n_14102)
);

INVx1_ASAP7_75t_SL g14103 ( 
.A(n_13941),
.Y(n_14103)
);

XNOR2x2_ASAP7_75t_L g14104 ( 
.A(n_13966),
.B(n_6872),
.Y(n_14104)
);

INVx1_ASAP7_75t_L g14105 ( 
.A(n_13901),
.Y(n_14105)
);

NOR2xp33_ASAP7_75t_L g14106 ( 
.A(n_13936),
.B(n_7259),
.Y(n_14106)
);

INVxp67_ASAP7_75t_SL g14107 ( 
.A(n_13953),
.Y(n_14107)
);

XOR2xp5_ASAP7_75t_L g14108 ( 
.A(n_13957),
.B(n_6896),
.Y(n_14108)
);

INVx1_ASAP7_75t_L g14109 ( 
.A(n_13881),
.Y(n_14109)
);

INVx1_ASAP7_75t_L g14110 ( 
.A(n_13878),
.Y(n_14110)
);

INVx1_ASAP7_75t_L g14111 ( 
.A(n_13947),
.Y(n_14111)
);

INVx1_ASAP7_75t_L g14112 ( 
.A(n_13973),
.Y(n_14112)
);

INVx1_ASAP7_75t_L g14113 ( 
.A(n_13978),
.Y(n_14113)
);

INVx1_ASAP7_75t_L g14114 ( 
.A(n_13960),
.Y(n_14114)
);

NAND2xp5_ASAP7_75t_L g14115 ( 
.A(n_13964),
.B(n_7259),
.Y(n_14115)
);

AOI32xp33_ASAP7_75t_L g14116 ( 
.A1(n_13819),
.A2(n_6873),
.A3(n_6893),
.B1(n_7906),
.B2(n_6755),
.Y(n_14116)
);

NOR2xp33_ASAP7_75t_L g14117 ( 
.A(n_13930),
.B(n_7262),
.Y(n_14117)
);

NAND2xp5_ASAP7_75t_SL g14118 ( 
.A(n_13876),
.B(n_6814),
.Y(n_14118)
);

INVx3_ASAP7_75t_L g14119 ( 
.A(n_13900),
.Y(n_14119)
);

AND2x2_ASAP7_75t_L g14120 ( 
.A(n_13928),
.B(n_7094),
.Y(n_14120)
);

NOR2x1_ASAP7_75t_L g14121 ( 
.A(n_14053),
.B(n_13963),
.Y(n_14121)
);

NAND2xp5_ASAP7_75t_SL g14122 ( 
.A(n_13999),
.B(n_13834),
.Y(n_14122)
);

OAI21x1_ASAP7_75t_SL g14123 ( 
.A1(n_14000),
.A2(n_13942),
.B(n_13946),
.Y(n_14123)
);

AOI21xp33_ASAP7_75t_SL g14124 ( 
.A1(n_14019),
.A2(n_13949),
.B(n_13945),
.Y(n_14124)
);

OAI21x1_ASAP7_75t_SL g14125 ( 
.A1(n_13990),
.A2(n_13883),
.B(n_13939),
.Y(n_14125)
);

AOI211xp5_ASAP7_75t_L g14126 ( 
.A1(n_13984),
.A2(n_13951),
.B(n_13948),
.C(n_13956),
.Y(n_14126)
);

NOR2x1_ASAP7_75t_L g14127 ( 
.A(n_14017),
.B(n_13908),
.Y(n_14127)
);

AOI22xp5_ASAP7_75t_L g14128 ( 
.A1(n_14005),
.A2(n_13954),
.B1(n_13977),
.B2(n_13921),
.Y(n_14128)
);

AOI22xp5_ASAP7_75t_L g14129 ( 
.A1(n_13989),
.A2(n_13918),
.B1(n_13962),
.B2(n_13943),
.Y(n_14129)
);

AOI22xp5_ASAP7_75t_L g14130 ( 
.A1(n_13997),
.A2(n_13952),
.B1(n_13961),
.B2(n_13970),
.Y(n_14130)
);

NOR3xp33_ASAP7_75t_L g14131 ( 
.A(n_13987),
.B(n_13851),
.C(n_13959),
.Y(n_14131)
);

AND2x2_ASAP7_75t_L g14132 ( 
.A(n_14059),
.B(n_13958),
.Y(n_14132)
);

AOI22xp5_ASAP7_75t_L g14133 ( 
.A1(n_14114),
.A2(n_13937),
.B1(n_6919),
.B2(n_7038),
.Y(n_14133)
);

NOR3xp33_ASAP7_75t_L g14134 ( 
.A(n_14010),
.B(n_6869),
.C(n_6853),
.Y(n_14134)
);

AND2x2_ASAP7_75t_L g14135 ( 
.A(n_14068),
.B(n_14029),
.Y(n_14135)
);

NAND2xp5_ASAP7_75t_L g14136 ( 
.A(n_14039),
.B(n_7262),
.Y(n_14136)
);

NOR2xp33_ASAP7_75t_L g14137 ( 
.A(n_14044),
.B(n_7262),
.Y(n_14137)
);

OAI21xp5_ASAP7_75t_L g14138 ( 
.A1(n_13993),
.A2(n_6761),
.B(n_6788),
.Y(n_14138)
);

NOR3x1_ASAP7_75t_L g14139 ( 
.A(n_14022),
.B(n_8017),
.C(n_7913),
.Y(n_14139)
);

NOR2xp33_ASAP7_75t_L g14140 ( 
.A(n_14070),
.B(n_7267),
.Y(n_14140)
);

NOR2x1_ASAP7_75t_L g14141 ( 
.A(n_13992),
.B(n_6814),
.Y(n_14141)
);

AOI22xp5_ASAP7_75t_L g14142 ( 
.A1(n_14038),
.A2(n_6919),
.B1(n_7038),
.B2(n_6814),
.Y(n_14142)
);

NOR2x1_ASAP7_75t_L g14143 ( 
.A(n_14015),
.B(n_6919),
.Y(n_14143)
);

INVx1_ASAP7_75t_L g14144 ( 
.A(n_14095),
.Y(n_14144)
);

AOI22xp5_ASAP7_75t_L g14145 ( 
.A1(n_14042),
.A2(n_7038),
.B1(n_7052),
.B2(n_6919),
.Y(n_14145)
);

AOI211x1_ASAP7_75t_L g14146 ( 
.A1(n_13986),
.A2(n_7320),
.B(n_5868),
.C(n_5873),
.Y(n_14146)
);

NAND2xp5_ASAP7_75t_L g14147 ( 
.A(n_14103),
.B(n_14062),
.Y(n_14147)
);

XOR2xp5_ASAP7_75t_SL g14148 ( 
.A(n_14082),
.B(n_7209),
.Y(n_14148)
);

OA22x2_ASAP7_75t_L g14149 ( 
.A1(n_14057),
.A2(n_7248),
.B1(n_8314),
.B2(n_8017),
.Y(n_14149)
);

AO22x2_ASAP7_75t_L g14150 ( 
.A1(n_14107),
.A2(n_7292),
.B1(n_7300),
.B2(n_7267),
.Y(n_14150)
);

INVx1_ASAP7_75t_L g14151 ( 
.A(n_14091),
.Y(n_14151)
);

AOI22xp5_ASAP7_75t_L g14152 ( 
.A1(n_13995),
.A2(n_7038),
.B1(n_7052),
.B2(n_6919),
.Y(n_14152)
);

XOR2x2_ASAP7_75t_L g14153 ( 
.A(n_14111),
.B(n_5550),
.Y(n_14153)
);

NOR3xp33_ASAP7_75t_L g14154 ( 
.A(n_14023),
.B(n_6869),
.C(n_6685),
.Y(n_14154)
);

NOR2xp33_ASAP7_75t_L g14155 ( 
.A(n_14025),
.B(n_7267),
.Y(n_14155)
);

NAND4xp75_ASAP7_75t_L g14156 ( 
.A(n_14027),
.B(n_14033),
.C(n_14034),
.D(n_14030),
.Y(n_14156)
);

OAI211xp5_ASAP7_75t_SL g14157 ( 
.A1(n_14101),
.A2(n_5841),
.B(n_5832),
.C(n_6386),
.Y(n_14157)
);

NOR4xp25_ASAP7_75t_L g14158 ( 
.A(n_14041),
.B(n_5832),
.C(n_5841),
.D(n_5866),
.Y(n_14158)
);

AOI21xp5_ASAP7_75t_L g14159 ( 
.A1(n_14058),
.A2(n_6240),
.B(n_6226),
.Y(n_14159)
);

AO22x2_ASAP7_75t_L g14160 ( 
.A1(n_14119),
.A2(n_7292),
.B1(n_7300),
.B2(n_7276),
.Y(n_14160)
);

AOI21xp5_ASAP7_75t_L g14161 ( 
.A1(n_14067),
.A2(n_6240),
.B(n_6226),
.Y(n_14161)
);

NOR2x1_ASAP7_75t_L g14162 ( 
.A(n_14119),
.B(n_7038),
.Y(n_14162)
);

NOR2x1_ASAP7_75t_L g14163 ( 
.A(n_14086),
.B(n_7052),
.Y(n_14163)
);

NAND4xp25_ASAP7_75t_L g14164 ( 
.A(n_14018),
.B(n_6948),
.C(n_7056),
.D(n_6937),
.Y(n_14164)
);

NOR3xp33_ASAP7_75t_L g14165 ( 
.A(n_14078),
.B(n_6685),
.C(n_6893),
.Y(n_14165)
);

INVx1_ASAP7_75t_L g14166 ( 
.A(n_14104),
.Y(n_14166)
);

NAND4xp25_ASAP7_75t_L g14167 ( 
.A(n_14001),
.B(n_7109),
.C(n_7088),
.D(n_7112),
.Y(n_14167)
);

NOR3xp33_ASAP7_75t_L g14168 ( 
.A(n_14052),
.B(n_6685),
.C(n_6893),
.Y(n_14168)
);

INVx2_ASAP7_75t_SL g14169 ( 
.A(n_14043),
.Y(n_14169)
);

NAND2xp5_ASAP7_75t_L g14170 ( 
.A(n_14066),
.B(n_7276),
.Y(n_14170)
);

INVx1_ASAP7_75t_L g14171 ( 
.A(n_13985),
.Y(n_14171)
);

OAI222xp33_ASAP7_75t_L g14172 ( 
.A1(n_13983),
.A2(n_6888),
.B1(n_6844),
.B2(n_6941),
.C1(n_6860),
.C2(n_6771),
.Y(n_14172)
);

NOR3x1_ASAP7_75t_L g14173 ( 
.A(n_14112),
.B(n_8052),
.C(n_7913),
.Y(n_14173)
);

NAND3xp33_ASAP7_75t_L g14174 ( 
.A(n_14052),
.B(n_7292),
.C(n_7276),
.Y(n_14174)
);

INVx2_ASAP7_75t_SL g14175 ( 
.A(n_14008),
.Y(n_14175)
);

AND2x2_ASAP7_75t_L g14176 ( 
.A(n_13994),
.B(n_6497),
.Y(n_14176)
);

OAI211xp5_ASAP7_75t_SL g14177 ( 
.A1(n_14049),
.A2(n_5584),
.B(n_6207),
.C(n_6200),
.Y(n_14177)
);

AOI21xp5_ASAP7_75t_L g14178 ( 
.A1(n_14113),
.A2(n_6265),
.B(n_6253),
.Y(n_14178)
);

NOR3x1_ASAP7_75t_L g14179 ( 
.A(n_14110),
.B(n_8052),
.C(n_8293),
.Y(n_14179)
);

INVx1_ASAP7_75t_L g14180 ( 
.A(n_14108),
.Y(n_14180)
);

INVx2_ASAP7_75t_L g14181 ( 
.A(n_14084),
.Y(n_14181)
);

OAI22xp33_ASAP7_75t_L g14182 ( 
.A1(n_14079),
.A2(n_7052),
.B1(n_6228),
.B2(n_6428),
.Y(n_14182)
);

NOR2x1_ASAP7_75t_L g14183 ( 
.A(n_14105),
.B(n_7052),
.Y(n_14183)
);

AOI21xp5_ASAP7_75t_L g14184 ( 
.A1(n_14088),
.A2(n_6265),
.B(n_6253),
.Y(n_14184)
);

NOR3xp33_ASAP7_75t_L g14185 ( 
.A(n_14075),
.B(n_14056),
.C(n_14051),
.Y(n_14185)
);

NOR2x1p5_ASAP7_75t_L g14186 ( 
.A(n_14064),
.B(n_7052),
.Y(n_14186)
);

AOI21xp5_ASAP7_75t_L g14187 ( 
.A1(n_14028),
.A2(n_6290),
.B(n_6269),
.Y(n_14187)
);

AOI211xp5_ASAP7_75t_SL g14188 ( 
.A1(n_14081),
.A2(n_6163),
.B(n_6166),
.C(n_6357),
.Y(n_14188)
);

NAND2xp5_ASAP7_75t_L g14189 ( 
.A(n_14092),
.B(n_7300),
.Y(n_14189)
);

OA22x2_ASAP7_75t_L g14190 ( 
.A1(n_14032),
.A2(n_8314),
.B1(n_8293),
.B2(n_5873),
.Y(n_14190)
);

OAI211xp5_ASAP7_75t_SL g14191 ( 
.A1(n_14109),
.A2(n_5584),
.B(n_6217),
.C(n_6200),
.Y(n_14191)
);

NAND2xp5_ASAP7_75t_L g14192 ( 
.A(n_14102),
.B(n_14046),
.Y(n_14192)
);

AOI22xp33_ASAP7_75t_L g14193 ( 
.A1(n_14089),
.A2(n_7304),
.B1(n_7327),
.B2(n_7311),
.Y(n_14193)
);

AND2x2_ASAP7_75t_SL g14194 ( 
.A(n_14099),
.B(n_7052),
.Y(n_14194)
);

INVx1_ASAP7_75t_L g14195 ( 
.A(n_13988),
.Y(n_14195)
);

NOR3x1_ASAP7_75t_L g14196 ( 
.A(n_14060),
.B(n_6819),
.C(n_6849),
.Y(n_14196)
);

AOI22xp5_ASAP7_75t_L g14197 ( 
.A1(n_14087),
.A2(n_7094),
.B1(n_7145),
.B2(n_7108),
.Y(n_14197)
);

AO22x2_ASAP7_75t_L g14198 ( 
.A1(n_14090),
.A2(n_7311),
.B1(n_7356),
.B2(n_7327),
.Y(n_14198)
);

AOI21xp5_ASAP7_75t_L g14199 ( 
.A1(n_14009),
.A2(n_6290),
.B(n_6269),
.Y(n_14199)
);

OAI222xp33_ASAP7_75t_L g14200 ( 
.A1(n_14002),
.A2(n_6771),
.B1(n_6860),
.B2(n_6941),
.C1(n_6888),
.C2(n_6844),
.Y(n_14200)
);

AOI31xp33_ASAP7_75t_L g14201 ( 
.A1(n_14093),
.A2(n_6888),
.A3(n_6941),
.B(n_6860),
.Y(n_14201)
);

NAND2xp5_ASAP7_75t_L g14202 ( 
.A(n_14072),
.B(n_7304),
.Y(n_14202)
);

XNOR2xp5_ASAP7_75t_L g14203 ( 
.A(n_14035),
.B(n_7109),
.Y(n_14203)
);

OAI211xp5_ASAP7_75t_SL g14204 ( 
.A1(n_14098),
.A2(n_6217),
.B(n_6224),
.C(n_6306),
.Y(n_14204)
);

NOR3xp33_ASAP7_75t_L g14205 ( 
.A(n_14012),
.B(n_6224),
.C(n_6761),
.Y(n_14205)
);

INVx1_ASAP7_75t_L g14206 ( 
.A(n_14054),
.Y(n_14206)
);

NAND2xp5_ASAP7_75t_L g14207 ( 
.A(n_14080),
.B(n_7304),
.Y(n_14207)
);

OAI22xp5_ASAP7_75t_L g14208 ( 
.A1(n_14100),
.A2(n_6025),
.B1(n_6428),
.B2(n_5868),
.Y(n_14208)
);

NAND2xp5_ASAP7_75t_L g14209 ( 
.A(n_14065),
.B(n_7311),
.Y(n_14209)
);

INVx2_ASAP7_75t_L g14210 ( 
.A(n_14120),
.Y(n_14210)
);

NOR2xp67_ASAP7_75t_L g14211 ( 
.A(n_14117),
.B(n_7094),
.Y(n_14211)
);

NOR2xp67_ASAP7_75t_L g14212 ( 
.A(n_13996),
.B(n_7094),
.Y(n_14212)
);

AO22x1_ASAP7_75t_L g14213 ( 
.A1(n_14011),
.A2(n_7108),
.B1(n_7177),
.B2(n_7145),
.Y(n_14213)
);

INVx1_ASAP7_75t_L g14214 ( 
.A(n_14055),
.Y(n_14214)
);

AOI21xp5_ASAP7_75t_L g14215 ( 
.A1(n_14094),
.A2(n_6316),
.B(n_6306),
.Y(n_14215)
);

INVx1_ASAP7_75t_L g14216 ( 
.A(n_14115),
.Y(n_14216)
);

OAI21xp5_ASAP7_75t_L g14217 ( 
.A1(n_14106),
.A2(n_6793),
.B(n_7327),
.Y(n_14217)
);

AO22x2_ASAP7_75t_L g14218 ( 
.A1(n_14097),
.A2(n_7358),
.B1(n_7366),
.B2(n_7356),
.Y(n_14218)
);

AOI21xp5_ASAP7_75t_L g14219 ( 
.A1(n_14069),
.A2(n_6318),
.B(n_6316),
.Y(n_14219)
);

OAI21x1_ASAP7_75t_SL g14220 ( 
.A1(n_14047),
.A2(n_14063),
.B(n_14096),
.Y(n_14220)
);

AOI211x1_ASAP7_75t_L g14221 ( 
.A1(n_14006),
.A2(n_7320),
.B(n_6149),
.C(n_6343),
.Y(n_14221)
);

NAND4xp25_ASAP7_75t_L g14222 ( 
.A(n_14014),
.B(n_7333),
.C(n_7370),
.D(n_7345),
.Y(n_14222)
);

OAI222xp33_ASAP7_75t_L g14223 ( 
.A1(n_14118),
.A2(n_6771),
.B1(n_6860),
.B2(n_6941),
.C1(n_6888),
.C2(n_6844),
.Y(n_14223)
);

INVx1_ASAP7_75t_SL g14224 ( 
.A(n_14071),
.Y(n_14224)
);

NOR3x1_ASAP7_75t_L g14225 ( 
.A(n_14003),
.B(n_6819),
.C(n_6849),
.Y(n_14225)
);

INVx2_ASAP7_75t_L g14226 ( 
.A(n_14004),
.Y(n_14226)
);

OAI211xp5_ASAP7_75t_SL g14227 ( 
.A1(n_14061),
.A2(n_6343),
.B(n_6350),
.C(n_6318),
.Y(n_14227)
);

AOI21xp5_ASAP7_75t_L g14228 ( 
.A1(n_14076),
.A2(n_6360),
.B(n_6350),
.Y(n_14228)
);

INVxp67_ASAP7_75t_SL g14229 ( 
.A(n_14073),
.Y(n_14229)
);

INVx1_ASAP7_75t_L g14230 ( 
.A(n_14045),
.Y(n_14230)
);

NOR2x1_ASAP7_75t_L g14231 ( 
.A(n_13998),
.B(n_7145),
.Y(n_14231)
);

AOI22xp5_ASAP7_75t_L g14232 ( 
.A1(n_14013),
.A2(n_7145),
.B1(n_7246),
.B2(n_7177),
.Y(n_14232)
);

AOI21xp5_ASAP7_75t_L g14233 ( 
.A1(n_14020),
.A2(n_6369),
.B(n_6360),
.Y(n_14233)
);

NAND2xp5_ASAP7_75t_L g14234 ( 
.A(n_14026),
.B(n_7356),
.Y(n_14234)
);

OA21x2_ASAP7_75t_L g14235 ( 
.A1(n_14007),
.A2(n_6723),
.B(n_6714),
.Y(n_14235)
);

AOI211xp5_ASAP7_75t_L g14236 ( 
.A1(n_14077),
.A2(n_5787),
.B(n_6800),
.C(n_6755),
.Y(n_14236)
);

INVxp33_ASAP7_75t_L g14237 ( 
.A(n_14016),
.Y(n_14237)
);

NAND2xp5_ASAP7_75t_L g14238 ( 
.A(n_14040),
.B(n_7358),
.Y(n_14238)
);

AOI21xp5_ASAP7_75t_L g14239 ( 
.A1(n_14036),
.A2(n_6371),
.B(n_6369),
.Y(n_14239)
);

NAND2xp5_ASAP7_75t_L g14240 ( 
.A(n_14031),
.B(n_7358),
.Y(n_14240)
);

NOR2x1p5_ASAP7_75t_L g14241 ( 
.A(n_13991),
.B(n_5834),
.Y(n_14241)
);

AOI22xp5_ASAP7_75t_L g14242 ( 
.A1(n_14135),
.A2(n_14037),
.B1(n_14024),
.B2(n_14021),
.Y(n_14242)
);

O2A1O1Ixp33_ASAP7_75t_L g14243 ( 
.A1(n_14144),
.A2(n_14085),
.B(n_14083),
.C(n_14050),
.Y(n_14243)
);

OAI21xp5_ASAP7_75t_L g14244 ( 
.A1(n_14151),
.A2(n_14048),
.B(n_14074),
.Y(n_14244)
);

OA22x2_ASAP7_75t_L g14245 ( 
.A1(n_14169),
.A2(n_14116),
.B1(n_7177),
.B2(n_7246),
.Y(n_14245)
);

INVxp67_ASAP7_75t_L g14246 ( 
.A(n_14147),
.Y(n_14246)
);

NOR2xp33_ASAP7_75t_L g14247 ( 
.A(n_14237),
.B(n_7399),
.Y(n_14247)
);

NAND2xp5_ASAP7_75t_L g14248 ( 
.A(n_14229),
.B(n_14166),
.Y(n_14248)
);

INVxp67_ASAP7_75t_L g14249 ( 
.A(n_14156),
.Y(n_14249)
);

BUFx12f_ASAP7_75t_L g14250 ( 
.A(n_14132),
.Y(n_14250)
);

OAI22xp5_ASAP7_75t_L g14251 ( 
.A1(n_14128),
.A2(n_6428),
.B1(n_7399),
.B2(n_7366),
.Y(n_14251)
);

XNOR2xp5_ASAP7_75t_L g14252 ( 
.A(n_14224),
.B(n_6497),
.Y(n_14252)
);

NAND2xp5_ASAP7_75t_L g14253 ( 
.A(n_14175),
.B(n_7366),
.Y(n_14253)
);

NOR2x1_ASAP7_75t_L g14254 ( 
.A(n_14127),
.B(n_14121),
.Y(n_14254)
);

AOI21xp5_ASAP7_75t_L g14255 ( 
.A1(n_14122),
.A2(n_6387),
.B(n_6371),
.Y(n_14255)
);

NAND2xp5_ASAP7_75t_L g14256 ( 
.A(n_14181),
.B(n_7283),
.Y(n_14256)
);

NOR2x1_ASAP7_75t_SL g14257 ( 
.A(n_14230),
.B(n_6401),
.Y(n_14257)
);

AOI32xp33_ASAP7_75t_L g14258 ( 
.A1(n_14131),
.A2(n_6755),
.A3(n_6723),
.B1(n_6714),
.B2(n_7145),
.Y(n_14258)
);

INVx2_ASAP7_75t_SL g14259 ( 
.A(n_14143),
.Y(n_14259)
);

AOI211xp5_ASAP7_75t_L g14260 ( 
.A1(n_14124),
.A2(n_5787),
.B(n_6800),
.C(n_6730),
.Y(n_14260)
);

AOI21xp33_ASAP7_75t_L g14261 ( 
.A1(n_14192),
.A2(n_7355),
.B(n_7349),
.Y(n_14261)
);

NAND2xp33_ASAP7_75t_L g14262 ( 
.A(n_14171),
.B(n_6771),
.Y(n_14262)
);

OAI332xp33_ASAP7_75t_L g14263 ( 
.A1(n_14180),
.A2(n_5630),
.A3(n_5657),
.B1(n_5576),
.B2(n_6373),
.B3(n_6390),
.C1(n_6384),
.C2(n_6313),
.Y(n_14263)
);

AND2x2_ASAP7_75t_L g14264 ( 
.A(n_14176),
.B(n_6497),
.Y(n_14264)
);

XNOR2x1_ASAP7_75t_L g14265 ( 
.A(n_14226),
.B(n_6617),
.Y(n_14265)
);

NAND2x1_ASAP7_75t_L g14266 ( 
.A(n_14163),
.B(n_6428),
.Y(n_14266)
);

AOI211xp5_ASAP7_75t_L g14267 ( 
.A1(n_14126),
.A2(n_6800),
.B(n_6730),
.C(n_6723),
.Y(n_14267)
);

AOI21xp5_ASAP7_75t_L g14268 ( 
.A1(n_14210),
.A2(n_6391),
.B(n_6387),
.Y(n_14268)
);

CKINVDCx5p33_ASAP7_75t_R g14269 ( 
.A(n_14216),
.Y(n_14269)
);

AOI221xp5_ASAP7_75t_L g14270 ( 
.A1(n_14137),
.A2(n_6391),
.B1(n_6438),
.B2(n_6402),
.C(n_5887),
.Y(n_14270)
);

O2A1O1Ixp5_ASAP7_75t_L g14271 ( 
.A1(n_14195),
.A2(n_7294),
.B(n_7301),
.C(n_7246),
.Y(n_14271)
);

NAND2xp5_ASAP7_75t_L g14272 ( 
.A(n_14185),
.B(n_7283),
.Y(n_14272)
);

AOI21xp33_ASAP7_75t_L g14273 ( 
.A1(n_14220),
.A2(n_7355),
.B(n_7349),
.Y(n_14273)
);

AOI322xp5_ASAP7_75t_L g14274 ( 
.A1(n_14140),
.A2(n_7181),
.A3(n_7333),
.B1(n_7370),
.B2(n_7374),
.C1(n_7345),
.C2(n_5576),
.Y(n_14274)
);

INVx1_ASAP7_75t_L g14275 ( 
.A(n_14141),
.Y(n_14275)
);

AOI221xp5_ASAP7_75t_L g14276 ( 
.A1(n_14123),
.A2(n_6438),
.B1(n_6402),
.B2(n_5887),
.C(n_5898),
.Y(n_14276)
);

AOI22xp5_ASAP7_75t_L g14277 ( 
.A1(n_14162),
.A2(n_7127),
.B1(n_7294),
.B2(n_7246),
.Y(n_14277)
);

AND2x2_ASAP7_75t_L g14278 ( 
.A(n_14211),
.B(n_6497),
.Y(n_14278)
);

AOI22xp5_ASAP7_75t_L g14279 ( 
.A1(n_14129),
.A2(n_14183),
.B1(n_14241),
.B2(n_14194),
.Y(n_14279)
);

AO221x1_ASAP7_75t_L g14280 ( 
.A1(n_14125),
.A2(n_6166),
.B1(n_6163),
.B2(n_5909),
.C(n_5902),
.Y(n_14280)
);

AOI221xp5_ASAP7_75t_L g14281 ( 
.A1(n_14206),
.A2(n_5898),
.B1(n_5901),
.B2(n_5881),
.C(n_5877),
.Y(n_14281)
);

AOI221xp5_ASAP7_75t_L g14282 ( 
.A1(n_14214),
.A2(n_5901),
.B1(n_5923),
.B2(n_5881),
.C(n_5877),
.Y(n_14282)
);

OAI211xp5_ASAP7_75t_L g14283 ( 
.A1(n_14130),
.A2(n_5902),
.B(n_5909),
.C(n_5900),
.Y(n_14283)
);

OAI22xp33_ASAP7_75t_L g14284 ( 
.A1(n_14133),
.A2(n_5834),
.B1(n_5855),
.B2(n_5852),
.Y(n_14284)
);

INVx1_ASAP7_75t_L g14285 ( 
.A(n_14136),
.Y(n_14285)
);

OAI21xp33_ASAP7_75t_L g14286 ( 
.A1(n_14153),
.A2(n_7294),
.B(n_7246),
.Y(n_14286)
);

INVx1_ASAP7_75t_L g14287 ( 
.A(n_14202),
.Y(n_14287)
);

AOI21xp5_ASAP7_75t_L g14288 ( 
.A1(n_14155),
.A2(n_6784),
.B(n_6765),
.Y(n_14288)
);

NOR2x1_ASAP7_75t_L g14289 ( 
.A(n_14186),
.B(n_6497),
.Y(n_14289)
);

AOI21xp33_ASAP7_75t_L g14290 ( 
.A1(n_14189),
.A2(n_7368),
.B(n_7355),
.Y(n_14290)
);

AOI22x1_ASAP7_75t_L g14291 ( 
.A1(n_14138),
.A2(n_6401),
.B1(n_5852),
.B2(n_5855),
.Y(n_14291)
);

NOR2xp33_ASAP7_75t_R g14292 ( 
.A(n_14170),
.B(n_6181),
.Y(n_14292)
);

OAI221xp5_ASAP7_75t_L g14293 ( 
.A1(n_14217),
.A2(n_6844),
.B1(n_5657),
.B2(n_5630),
.C(n_5576),
.Y(n_14293)
);

INVx1_ASAP7_75t_L g14294 ( 
.A(n_14207),
.Y(n_14294)
);

AO221x1_ASAP7_75t_L g14295 ( 
.A1(n_14182),
.A2(n_5909),
.B1(n_5902),
.B2(n_5900),
.C(n_5565),
.Y(n_14295)
);

NAND2xp5_ASAP7_75t_L g14296 ( 
.A(n_14209),
.B(n_7337),
.Y(n_14296)
);

AOI221xp5_ASAP7_75t_L g14297 ( 
.A1(n_14158),
.A2(n_5923),
.B1(n_5944),
.B2(n_5943),
.C(n_5929),
.Y(n_14297)
);

O2A1O1Ixp33_ASAP7_75t_L g14298 ( 
.A1(n_14234),
.A2(n_5630),
.B(n_5657),
.C(n_5715),
.Y(n_14298)
);

NAND5xp2_ASAP7_75t_L g14299 ( 
.A(n_14238),
.B(n_7181),
.C(n_5550),
.D(n_7374),
.E(n_6267),
.Y(n_14299)
);

O2A1O1Ixp33_ASAP7_75t_L g14300 ( 
.A1(n_14240),
.A2(n_14177),
.B(n_14191),
.C(n_14208),
.Y(n_14300)
);

INVx1_ASAP7_75t_L g14301 ( 
.A(n_14203),
.Y(n_14301)
);

INVx1_ASAP7_75t_L g14302 ( 
.A(n_14231),
.Y(n_14302)
);

OAI22xp5_ASAP7_75t_L g14303 ( 
.A1(n_14142),
.A2(n_6209),
.B1(n_6220),
.B2(n_6034),
.Y(n_14303)
);

AOI22xp5_ASAP7_75t_L g14304 ( 
.A1(n_14212),
.A2(n_7301),
.B1(n_7319),
.B2(n_7294),
.Y(n_14304)
);

OAI22xp33_ASAP7_75t_L g14305 ( 
.A1(n_14145),
.A2(n_5834),
.B1(n_5855),
.B2(n_5852),
.Y(n_14305)
);

OAI321xp33_ASAP7_75t_L g14306 ( 
.A1(n_14174),
.A2(n_5849),
.A3(n_5797),
.B1(n_5889),
.B2(n_5817),
.C(n_5715),
.Y(n_14306)
);

AOI21xp33_ASAP7_75t_L g14307 ( 
.A1(n_14190),
.A2(n_7368),
.B(n_7355),
.Y(n_14307)
);

NAND2xp5_ASAP7_75t_L g14308 ( 
.A(n_14221),
.B(n_7337),
.Y(n_14308)
);

AO21x1_ASAP7_75t_L g14309 ( 
.A1(n_14161),
.A2(n_7301),
.B(n_7294),
.Y(n_14309)
);

AO22x1_ASAP7_75t_L g14310 ( 
.A1(n_14139),
.A2(n_7301),
.B1(n_7364),
.B2(n_7319),
.Y(n_14310)
);

AOI221xp5_ASAP7_75t_L g14311 ( 
.A1(n_14213),
.A2(n_5944),
.B1(n_5945),
.B2(n_5943),
.C(n_5929),
.Y(n_14311)
);

AOI22xp5_ASAP7_75t_L g14312 ( 
.A1(n_14235),
.A2(n_7319),
.B1(n_7364),
.B2(n_7301),
.Y(n_14312)
);

INVx1_ASAP7_75t_L g14313 ( 
.A(n_14218),
.Y(n_14313)
);

INVx1_ASAP7_75t_SL g14314 ( 
.A(n_14184),
.Y(n_14314)
);

INVx1_ASAP7_75t_L g14315 ( 
.A(n_14218),
.Y(n_14315)
);

INVx1_ASAP7_75t_L g14316 ( 
.A(n_14150),
.Y(n_14316)
);

INVx2_ASAP7_75t_L g14317 ( 
.A(n_14150),
.Y(n_14317)
);

NOR2xp33_ASAP7_75t_SL g14318 ( 
.A(n_14222),
.B(n_6540),
.Y(n_14318)
);

A2O1A1Ixp33_ASAP7_75t_L g14319 ( 
.A1(n_14215),
.A2(n_14219),
.B(n_14239),
.C(n_14178),
.Y(n_14319)
);

OAI21xp5_ASAP7_75t_L g14320 ( 
.A1(n_14205),
.A2(n_6784),
.B(n_6765),
.Y(n_14320)
);

AND3x4_ASAP7_75t_L g14321 ( 
.A(n_14165),
.B(n_6831),
.C(n_6628),
.Y(n_14321)
);

AOI221x1_ASAP7_75t_L g14322 ( 
.A1(n_14227),
.A2(n_7319),
.B1(n_7365),
.B2(n_7364),
.C(n_6385),
.Y(n_14322)
);

AOI21xp5_ASAP7_75t_L g14323 ( 
.A1(n_14148),
.A2(n_6784),
.B(n_6765),
.Y(n_14323)
);

AOI21xp5_ASAP7_75t_L g14324 ( 
.A1(n_14159),
.A2(n_6795),
.B(n_6714),
.Y(n_14324)
);

AOI22xp5_ASAP7_75t_L g14325 ( 
.A1(n_14235),
.A2(n_7364),
.B1(n_7319),
.B2(n_6365),
.Y(n_14325)
);

INVx1_ASAP7_75t_L g14326 ( 
.A(n_14198),
.Y(n_14326)
);

NOR2xp33_ASAP7_75t_L g14327 ( 
.A(n_14204),
.B(n_7117),
.Y(n_14327)
);

INVx1_ASAP7_75t_L g14328 ( 
.A(n_14198),
.Y(n_14328)
);

INVx2_ASAP7_75t_L g14329 ( 
.A(n_14160),
.Y(n_14329)
);

NAND2xp5_ASAP7_75t_SL g14330 ( 
.A(n_14152),
.B(n_6831),
.Y(n_14330)
);

INVx1_ASAP7_75t_L g14331 ( 
.A(n_14160),
.Y(n_14331)
);

NAND4xp75_ASAP7_75t_L g14332 ( 
.A(n_14225),
.B(n_5797),
.C(n_5817),
.D(n_5715),
.Y(n_14332)
);

AOI322xp5_ASAP7_75t_L g14333 ( 
.A1(n_14154),
.A2(n_6335),
.A3(n_5849),
.B1(n_5889),
.B2(n_5797),
.C1(n_5921),
.C2(n_5915),
.Y(n_14333)
);

INVx1_ASAP7_75t_L g14334 ( 
.A(n_14146),
.Y(n_14334)
);

AO22x2_ASAP7_75t_L g14335 ( 
.A1(n_14187),
.A2(n_6385),
.B1(n_6357),
.B2(n_5963),
.Y(n_14335)
);

NAND2xp5_ASAP7_75t_L g14336 ( 
.A(n_14199),
.B(n_7337),
.Y(n_14336)
);

AOI21xp33_ASAP7_75t_L g14337 ( 
.A1(n_14193),
.A2(n_7408),
.B(n_7368),
.Y(n_14337)
);

AOI21xp5_ASAP7_75t_L g14338 ( 
.A1(n_14233),
.A2(n_6795),
.B(n_6777),
.Y(n_14338)
);

INVx1_ASAP7_75t_L g14339 ( 
.A(n_14173),
.Y(n_14339)
);

INVx1_ASAP7_75t_L g14340 ( 
.A(n_14179),
.Y(n_14340)
);

NOR4xp75_ASAP7_75t_L g14341 ( 
.A(n_14248),
.B(n_14196),
.C(n_14157),
.D(n_14188),
.Y(n_14341)
);

AOI322xp5_ASAP7_75t_L g14342 ( 
.A1(n_14254),
.A2(n_14134),
.A3(n_14168),
.B1(n_14197),
.B2(n_14232),
.C1(n_14172),
.C2(n_14236),
.Y(n_14342)
);

OAI211xp5_ASAP7_75t_L g14343 ( 
.A1(n_14249),
.A2(n_14228),
.B(n_14164),
.C(n_14167),
.Y(n_14343)
);

AOI221xp5_ASAP7_75t_L g14344 ( 
.A1(n_14246),
.A2(n_14201),
.B1(n_14223),
.B2(n_14200),
.C(n_14149),
.Y(n_14344)
);

AND2x2_ASAP7_75t_L g14345 ( 
.A(n_14278),
.B(n_7209),
.Y(n_14345)
);

INVx1_ASAP7_75t_L g14346 ( 
.A(n_14250),
.Y(n_14346)
);

AOI222xp33_ASAP7_75t_L g14347 ( 
.A1(n_14339),
.A2(n_5966),
.B1(n_5945),
.B2(n_5971),
.C1(n_5967),
.C2(n_5963),
.Y(n_14347)
);

OAI22xp33_ASAP7_75t_L g14348 ( 
.A1(n_14340),
.A2(n_5834),
.B1(n_5855),
.B2(n_5852),
.Y(n_14348)
);

NAND4xp25_ASAP7_75t_L g14349 ( 
.A(n_14242),
.B(n_14243),
.C(n_14279),
.D(n_14244),
.Y(n_14349)
);

INVx1_ASAP7_75t_L g14350 ( 
.A(n_14316),
.Y(n_14350)
);

INVx1_ASAP7_75t_L g14351 ( 
.A(n_14317),
.Y(n_14351)
);

NOR3xp33_ASAP7_75t_L g14352 ( 
.A(n_14269),
.B(n_5852),
.C(n_5834),
.Y(n_14352)
);

HAxp5_ASAP7_75t_SL g14353 ( 
.A(n_14301),
.B(n_4326),
.CON(n_14353),
.SN(n_14353)
);

AOI211xp5_ASAP7_75t_L g14354 ( 
.A1(n_14302),
.A2(n_6777),
.B(n_6827),
.C(n_6823),
.Y(n_14354)
);

NAND4xp25_ASAP7_75t_L g14355 ( 
.A(n_14294),
.B(n_6335),
.C(n_6267),
.D(n_5747),
.Y(n_14355)
);

OAI211xp5_ASAP7_75t_SL g14356 ( 
.A1(n_14285),
.A2(n_6209),
.B(n_6220),
.C(n_6034),
.Y(n_14356)
);

AOI22xp33_ASAP7_75t_SL g14357 ( 
.A1(n_14257),
.A2(n_5706),
.B1(n_5752),
.B2(n_5747),
.Y(n_14357)
);

NOR3xp33_ASAP7_75t_L g14358 ( 
.A(n_14287),
.B(n_5910),
.C(n_5855),
.Y(n_14358)
);

OAI221xp5_ASAP7_75t_L g14359 ( 
.A1(n_14259),
.A2(n_5900),
.B1(n_5982),
.B2(n_6036),
.C(n_5910),
.Y(n_14359)
);

AOI322xp5_ASAP7_75t_L g14360 ( 
.A1(n_14247),
.A2(n_5889),
.A3(n_5817),
.B1(n_5915),
.B2(n_5921),
.C1(n_5849),
.C2(n_7364),
.Y(n_14360)
);

NAND2xp5_ASAP7_75t_L g14361 ( 
.A(n_14313),
.B(n_7337),
.Y(n_14361)
);

AOI21xp33_ASAP7_75t_L g14362 ( 
.A1(n_14315),
.A2(n_7408),
.B(n_7368),
.Y(n_14362)
);

OAI22xp5_ASAP7_75t_L g14363 ( 
.A1(n_14266),
.A2(n_6220),
.B1(n_6227),
.B2(n_6209),
.Y(n_14363)
);

INVx2_ASAP7_75t_L g14364 ( 
.A(n_14329),
.Y(n_14364)
);

AOI221xp5_ASAP7_75t_L g14365 ( 
.A1(n_14275),
.A2(n_14334),
.B1(n_14328),
.B2(n_14326),
.C(n_14331),
.Y(n_14365)
);

O2A1O1Ixp33_ASAP7_75t_L g14366 ( 
.A1(n_14314),
.A2(n_5921),
.B(n_5915),
.C(n_5382),
.Y(n_14366)
);

AO21x1_ASAP7_75t_L g14367 ( 
.A1(n_14300),
.A2(n_5982),
.B(n_5910),
.Y(n_14367)
);

XNOR2x1_ASAP7_75t_L g14368 ( 
.A(n_14265),
.B(n_6625),
.Y(n_14368)
);

A2O1A1Ixp33_ASAP7_75t_L g14369 ( 
.A1(n_14272),
.A2(n_6996),
.B(n_7206),
.C(n_7201),
.Y(n_14369)
);

AND2x2_ASAP7_75t_L g14370 ( 
.A(n_14289),
.B(n_7209),
.Y(n_14370)
);

NAND3xp33_ASAP7_75t_L g14371 ( 
.A(n_14252),
.B(n_4326),
.C(n_5884),
.Y(n_14371)
);

AOI221xp5_ASAP7_75t_L g14372 ( 
.A1(n_14319),
.A2(n_5971),
.B1(n_5972),
.B2(n_5967),
.C(n_5966),
.Y(n_14372)
);

AOI22xp5_ASAP7_75t_L g14373 ( 
.A1(n_14318),
.A2(n_6365),
.B1(n_6353),
.B2(n_6795),
.Y(n_14373)
);

AOI211x1_ASAP7_75t_L g14374 ( 
.A1(n_14283),
.A2(n_6393),
.B(n_6408),
.C(n_5973),
.Y(n_14374)
);

O2A1O1Ixp33_ASAP7_75t_L g14375 ( 
.A1(n_14253),
.A2(n_5382),
.B(n_5508),
.C(n_5449),
.Y(n_14375)
);

AOI21xp5_ASAP7_75t_L g14376 ( 
.A1(n_14256),
.A2(n_14323),
.B(n_14296),
.Y(n_14376)
);

NOR3xp33_ASAP7_75t_L g14377 ( 
.A(n_14251),
.B(n_5982),
.C(n_5910),
.Y(n_14377)
);

NOR2xp33_ASAP7_75t_R g14378 ( 
.A(n_14262),
.B(n_6181),
.Y(n_14378)
);

INVx2_ASAP7_75t_SL g14379 ( 
.A(n_14264),
.Y(n_14379)
);

AOI221xp5_ASAP7_75t_L g14380 ( 
.A1(n_14337),
.A2(n_5980),
.B1(n_5985),
.B2(n_5973),
.C(n_5972),
.Y(n_14380)
);

AOI221xp5_ASAP7_75t_L g14381 ( 
.A1(n_14261),
.A2(n_5999),
.B1(n_6022),
.B2(n_5985),
.C(n_5980),
.Y(n_14381)
);

NAND2xp5_ASAP7_75t_L g14382 ( 
.A(n_14292),
.B(n_7337),
.Y(n_14382)
);

AOI21xp5_ASAP7_75t_L g14383 ( 
.A1(n_14245),
.A2(n_6777),
.B(n_6022),
.Y(n_14383)
);

NOR4xp25_ASAP7_75t_L g14384 ( 
.A(n_14308),
.B(n_6308),
.C(n_6311),
.D(n_6227),
.Y(n_14384)
);

OAI321xp33_ASAP7_75t_L g14385 ( 
.A1(n_14336),
.A2(n_6308),
.A3(n_6311),
.B1(n_6227),
.B2(n_6072),
.C(n_6061),
.Y(n_14385)
);

O2A1O1Ixp33_ASAP7_75t_L g14386 ( 
.A1(n_14330),
.A2(n_5382),
.B(n_5508),
.C(n_5449),
.Y(n_14386)
);

O2A1O1Ixp33_ASAP7_75t_L g14387 ( 
.A1(n_14273),
.A2(n_5449),
.B(n_5508),
.C(n_6831),
.Y(n_14387)
);

INVx1_ASAP7_75t_L g14388 ( 
.A(n_14332),
.Y(n_14388)
);

OAI21xp33_ASAP7_75t_SL g14389 ( 
.A1(n_14295),
.A2(n_7264),
.B(n_7261),
.Y(n_14389)
);

NOR3xp33_ASAP7_75t_L g14390 ( 
.A(n_14310),
.B(n_5982),
.C(n_5910),
.Y(n_14390)
);

AOI211xp5_ASAP7_75t_L g14391 ( 
.A1(n_14309),
.A2(n_6827),
.B(n_6834),
.C(n_6823),
.Y(n_14391)
);

OAI21xp33_ASAP7_75t_SL g14392 ( 
.A1(n_14280),
.A2(n_7264),
.B(n_7261),
.Y(n_14392)
);

NOR2xp33_ASAP7_75t_L g14393 ( 
.A(n_14321),
.B(n_7117),
.Y(n_14393)
);

AOI221xp5_ASAP7_75t_L g14394 ( 
.A1(n_14290),
.A2(n_6068),
.B1(n_6072),
.B2(n_6061),
.C(n_5999),
.Y(n_14394)
);

NOR2xp33_ASAP7_75t_L g14395 ( 
.A(n_14327),
.B(n_7117),
.Y(n_14395)
);

AOI221xp5_ASAP7_75t_L g14396 ( 
.A1(n_14307),
.A2(n_6088),
.B1(n_6089),
.B2(n_6084),
.C(n_6068),
.Y(n_14396)
);

OAI21xp33_ASAP7_75t_SL g14397 ( 
.A1(n_14311),
.A2(n_7264),
.B(n_7261),
.Y(n_14397)
);

INVx1_ASAP7_75t_L g14398 ( 
.A(n_14291),
.Y(n_14398)
);

OAI211xp5_ASAP7_75t_L g14399 ( 
.A1(n_14268),
.A2(n_6036),
.B(n_6063),
.C(n_5982),
.Y(n_14399)
);

OAI221xp5_ASAP7_75t_L g14400 ( 
.A1(n_14258),
.A2(n_6063),
.B1(n_6095),
.B2(n_6085),
.C(n_6036),
.Y(n_14400)
);

AOI21xp33_ASAP7_75t_SL g14401 ( 
.A1(n_14284),
.A2(n_6662),
.B(n_6823),
.Y(n_14401)
);

AND2x4_ASAP7_75t_L g14402 ( 
.A(n_14255),
.B(n_5858),
.Y(n_14402)
);

AOI22xp5_ASAP7_75t_L g14403 ( 
.A1(n_14325),
.A2(n_6365),
.B1(n_6353),
.B2(n_6831),
.Y(n_14403)
);

AOI21xp33_ASAP7_75t_L g14404 ( 
.A1(n_14320),
.A2(n_7408),
.B(n_7378),
.Y(n_14404)
);

OAI21xp5_ASAP7_75t_L g14405 ( 
.A1(n_14324),
.A2(n_6764),
.B(n_6898),
.Y(n_14405)
);

INVx2_ASAP7_75t_L g14406 ( 
.A(n_14335),
.Y(n_14406)
);

AOI21xp33_ASAP7_75t_L g14407 ( 
.A1(n_14286),
.A2(n_14298),
.B(n_14276),
.Y(n_14407)
);

NAND2xp33_ASAP7_75t_R g14408 ( 
.A(n_14338),
.B(n_6831),
.Y(n_14408)
);

AOI221x1_ASAP7_75t_L g14409 ( 
.A1(n_14335),
.A2(n_6393),
.B1(n_6408),
.B2(n_6310),
.C(n_6089),
.Y(n_14409)
);

OAI21xp33_ASAP7_75t_L g14410 ( 
.A1(n_14299),
.A2(n_5955),
.B(n_5932),
.Y(n_14410)
);

OAI211xp5_ASAP7_75t_L g14411 ( 
.A1(n_14322),
.A2(n_14260),
.B(n_14333),
.C(n_14267),
.Y(n_14411)
);

O2A1O1Ixp33_ASAP7_75t_L g14412 ( 
.A1(n_14293),
.A2(n_5706),
.B(n_5752),
.C(n_5747),
.Y(n_14412)
);

AOI21xp5_ASAP7_75t_L g14413 ( 
.A1(n_14288),
.A2(n_6088),
.B(n_6084),
.Y(n_14413)
);

AOI221xp5_ASAP7_75t_L g14414 ( 
.A1(n_14281),
.A2(n_6125),
.B1(n_6127),
.B2(n_6106),
.C(n_6091),
.Y(n_14414)
);

OAI22xp33_ASAP7_75t_L g14415 ( 
.A1(n_14312),
.A2(n_6063),
.B1(n_6085),
.B2(n_6036),
.Y(n_14415)
);

AOI221xp5_ASAP7_75t_L g14416 ( 
.A1(n_14282),
.A2(n_6125),
.B1(n_6127),
.B2(n_6106),
.C(n_6091),
.Y(n_14416)
);

AOI221xp5_ASAP7_75t_L g14417 ( 
.A1(n_14306),
.A2(n_6139),
.B1(n_6134),
.B2(n_4788),
.C(n_4832),
.Y(n_14417)
);

OAI211xp5_ASAP7_75t_L g14418 ( 
.A1(n_14304),
.A2(n_6063),
.B(n_6085),
.C(n_6036),
.Y(n_14418)
);

NOR2xp33_ASAP7_75t_L g14419 ( 
.A(n_14303),
.B(n_7117),
.Y(n_14419)
);

AOI211xp5_ASAP7_75t_SL g14420 ( 
.A1(n_14305),
.A2(n_6310),
.B(n_6334),
.C(n_5561),
.Y(n_14420)
);

AOI211xp5_ASAP7_75t_L g14421 ( 
.A1(n_14297),
.A2(n_14263),
.B(n_14277),
.C(n_14270),
.Y(n_14421)
);

OAI211xp5_ASAP7_75t_SL g14422 ( 
.A1(n_14271),
.A2(n_6311),
.B(n_6308),
.C(n_5561),
.Y(n_14422)
);

NAND4xp75_ASAP7_75t_L g14423 ( 
.A(n_14274),
.B(n_6353),
.C(n_6334),
.D(n_6139),
.Y(n_14423)
);

AND2x2_ASAP7_75t_L g14424 ( 
.A(n_14254),
.B(n_7209),
.Y(n_14424)
);

AOI211xp5_ASAP7_75t_L g14425 ( 
.A1(n_14249),
.A2(n_6834),
.B(n_6827),
.C(n_6849),
.Y(n_14425)
);

NAND4xp25_ASAP7_75t_L g14426 ( 
.A(n_14254),
.B(n_5752),
.C(n_5762),
.D(n_5753),
.Y(n_14426)
);

AOI21xp5_ASAP7_75t_L g14427 ( 
.A1(n_14248),
.A2(n_6134),
.B(n_6898),
.Y(n_14427)
);

AOI221xp5_ASAP7_75t_L g14428 ( 
.A1(n_14249),
.A2(n_4788),
.B1(n_4832),
.B2(n_4829),
.C(n_4692),
.Y(n_14428)
);

AOI322xp5_ASAP7_75t_L g14429 ( 
.A1(n_14254),
.A2(n_6691),
.A3(n_6540),
.B1(n_6783),
.B2(n_6817),
.C1(n_6628),
.C2(n_5704),
.Y(n_14429)
);

OAI21xp33_ASAP7_75t_L g14430 ( 
.A1(n_14254),
.A2(n_5955),
.B(n_5932),
.Y(n_14430)
);

NAND4xp75_ASAP7_75t_L g14431 ( 
.A(n_14346),
.B(n_6404),
.C(n_6421),
.D(n_6372),
.Y(n_14431)
);

NAND2xp5_ASAP7_75t_L g14432 ( 
.A(n_14379),
.B(n_7209),
.Y(n_14432)
);

INVx2_ASAP7_75t_L g14433 ( 
.A(n_14406),
.Y(n_14433)
);

NOR3x1_ASAP7_75t_L g14434 ( 
.A(n_14349),
.B(n_6996),
.C(n_6834),
.Y(n_14434)
);

INVx1_ASAP7_75t_L g14435 ( 
.A(n_14364),
.Y(n_14435)
);

NOR2xp33_ASAP7_75t_L g14436 ( 
.A(n_14350),
.B(n_6625),
.Y(n_14436)
);

NOR3xp33_ASAP7_75t_L g14437 ( 
.A(n_14365),
.B(n_5438),
.C(n_6063),
.Y(n_14437)
);

INVx1_ASAP7_75t_L g14438 ( 
.A(n_14351),
.Y(n_14438)
);

NAND2xp5_ASAP7_75t_L g14439 ( 
.A(n_14376),
.B(n_7209),
.Y(n_14439)
);

NAND2xp5_ASAP7_75t_L g14440 ( 
.A(n_14424),
.B(n_7209),
.Y(n_14440)
);

AO22x2_ASAP7_75t_L g14441 ( 
.A1(n_14398),
.A2(n_6095),
.B1(n_6113),
.B2(n_6085),
.Y(n_14441)
);

NOR2x1p5_ASAP7_75t_L g14442 ( 
.A(n_14388),
.B(n_5752),
.Y(n_14442)
);

AND2x2_ASAP7_75t_L g14443 ( 
.A(n_14370),
.B(n_7193),
.Y(n_14443)
);

NAND3xp33_ASAP7_75t_SL g14444 ( 
.A(n_14341),
.B(n_4420),
.C(n_4376),
.Y(n_14444)
);

NAND3xp33_ASAP7_75t_L g14445 ( 
.A(n_14343),
.B(n_6628),
.C(n_6540),
.Y(n_14445)
);

AOI22xp5_ASAP7_75t_L g14446 ( 
.A1(n_14344),
.A2(n_14411),
.B1(n_14361),
.B2(n_14408),
.Y(n_14446)
);

AO22x2_ASAP7_75t_L g14447 ( 
.A1(n_14368),
.A2(n_6095),
.B1(n_6113),
.B2(n_6085),
.Y(n_14447)
);

NOR3xp33_ASAP7_75t_L g14448 ( 
.A(n_14407),
.B(n_6113),
.C(n_6095),
.Y(n_14448)
);

INVx1_ASAP7_75t_L g14449 ( 
.A(n_14421),
.Y(n_14449)
);

INVx1_ASAP7_75t_L g14450 ( 
.A(n_14382),
.Y(n_14450)
);

AOI22xp5_ASAP7_75t_L g14451 ( 
.A1(n_14393),
.A2(n_14430),
.B1(n_14371),
.B2(n_14423),
.Y(n_14451)
);

NAND2xp5_ASAP7_75t_L g14452 ( 
.A(n_14342),
.B(n_14395),
.Y(n_14452)
);

NOR2xp33_ASAP7_75t_L g14453 ( 
.A(n_14385),
.B(n_6625),
.Y(n_14453)
);

INVx1_ASAP7_75t_L g14454 ( 
.A(n_14387),
.Y(n_14454)
);

NAND4xp25_ASAP7_75t_L g14455 ( 
.A(n_14386),
.B(n_5762),
.C(n_5764),
.D(n_5753),
.Y(n_14455)
);

INVx2_ASAP7_75t_L g14456 ( 
.A(n_14402),
.Y(n_14456)
);

NOR2xp67_ASAP7_75t_L g14457 ( 
.A(n_14400),
.B(n_5884),
.Y(n_14457)
);

INVx1_ASAP7_75t_L g14458 ( 
.A(n_14378),
.Y(n_14458)
);

NAND3xp33_ASAP7_75t_L g14459 ( 
.A(n_14353),
.B(n_6628),
.C(n_6540),
.Y(n_14459)
);

NOR3xp33_ASAP7_75t_L g14460 ( 
.A(n_14396),
.B(n_6113),
.C(n_6095),
.Y(n_14460)
);

NAND4xp25_ASAP7_75t_L g14461 ( 
.A(n_14410),
.B(n_5762),
.C(n_5764),
.D(n_5753),
.Y(n_14461)
);

AND2x4_ASAP7_75t_L g14462 ( 
.A(n_14402),
.B(n_6540),
.Y(n_14462)
);

NAND3xp33_ASAP7_75t_SL g14463 ( 
.A(n_14367),
.B(n_4420),
.C(n_6113),
.Y(n_14463)
);

OAI21xp33_ASAP7_75t_L g14464 ( 
.A1(n_14384),
.A2(n_6691),
.B(n_6628),
.Y(n_14464)
);

NOR2x1_ASAP7_75t_L g14465 ( 
.A(n_14422),
.B(n_5753),
.Y(n_14465)
);

INVx2_ASAP7_75t_L g14466 ( 
.A(n_14374),
.Y(n_14466)
);

OAI21xp5_ASAP7_75t_SL g14467 ( 
.A1(n_14404),
.A2(n_6783),
.B(n_6691),
.Y(n_14467)
);

AOI22xp5_ASAP7_75t_L g14468 ( 
.A1(n_14419),
.A2(n_4692),
.B1(n_4829),
.B2(n_4788),
.Y(n_14468)
);

OAI221xp5_ASAP7_75t_SL g14469 ( 
.A1(n_14392),
.A2(n_6384),
.B1(n_6395),
.B2(n_6429),
.C(n_6390),
.Y(n_14469)
);

OAI321xp33_ASAP7_75t_L g14470 ( 
.A1(n_14415),
.A2(n_6943),
.A3(n_6773),
.B1(n_7055),
.B2(n_6797),
.C(n_6625),
.Y(n_14470)
);

NOR3xp33_ASAP7_75t_L g14471 ( 
.A(n_14380),
.B(n_6367),
.C(n_6662),
.Y(n_14471)
);

NAND4xp75_ASAP7_75t_L g14472 ( 
.A(n_14409),
.B(n_14383),
.C(n_14397),
.D(n_14427),
.Y(n_14472)
);

NAND2x1_ASAP7_75t_L g14473 ( 
.A(n_14390),
.B(n_6691),
.Y(n_14473)
);

NAND2xp5_ASAP7_75t_L g14474 ( 
.A(n_14394),
.B(n_7337),
.Y(n_14474)
);

INVx2_ASAP7_75t_SL g14475 ( 
.A(n_14363),
.Y(n_14475)
);

NOR4xp75_ASAP7_75t_L g14476 ( 
.A(n_14405),
.B(n_5955),
.C(n_6002),
.D(n_5932),
.Y(n_14476)
);

INVx1_ASAP7_75t_L g14477 ( 
.A(n_14413),
.Y(n_14477)
);

NAND2xp5_ASAP7_75t_SL g14478 ( 
.A(n_14357),
.B(n_6691),
.Y(n_14478)
);

INVx1_ASAP7_75t_L g14479 ( 
.A(n_14381),
.Y(n_14479)
);

NAND2xp5_ASAP7_75t_L g14480 ( 
.A(n_14362),
.B(n_7337),
.Y(n_14480)
);

OAI21xp5_ASAP7_75t_SL g14481 ( 
.A1(n_14377),
.A2(n_6817),
.B(n_6783),
.Y(n_14481)
);

NOR2x1_ASAP7_75t_L g14482 ( 
.A(n_14375),
.B(n_14426),
.Y(n_14482)
);

AOI22xp5_ASAP7_75t_L g14483 ( 
.A1(n_14373),
.A2(n_4692),
.B1(n_4829),
.B2(n_4788),
.Y(n_14483)
);

NAND3xp33_ASAP7_75t_SL g14484 ( 
.A(n_14352),
.B(n_4420),
.C(n_6367),
.Y(n_14484)
);

NOR3xp33_ASAP7_75t_L g14485 ( 
.A(n_14418),
.B(n_6367),
.C(n_6662),
.Y(n_14485)
);

NAND3xp33_ASAP7_75t_L g14486 ( 
.A(n_14369),
.B(n_6817),
.C(n_6783),
.Y(n_14486)
);

OAI21xp33_ASAP7_75t_L g14487 ( 
.A1(n_14403),
.A2(n_6817),
.B(n_6783),
.Y(n_14487)
);

NAND3xp33_ASAP7_75t_SL g14488 ( 
.A(n_14366),
.B(n_4420),
.C(n_6367),
.Y(n_14488)
);

AND2x2_ASAP7_75t_SL g14489 ( 
.A(n_14358),
.B(n_6817),
.Y(n_14489)
);

NOR2xp33_ASAP7_75t_L g14490 ( 
.A(n_14401),
.B(n_6797),
.Y(n_14490)
);

OR3x1_ASAP7_75t_L g14491 ( 
.A(n_14356),
.B(n_4993),
.C(n_4971),
.Y(n_14491)
);

NOR2xp33_ASAP7_75t_L g14492 ( 
.A(n_14399),
.B(n_6797),
.Y(n_14492)
);

NOR3xp33_ASAP7_75t_L g14493 ( 
.A(n_14348),
.B(n_6367),
.C(n_6670),
.Y(n_14493)
);

NAND2xp5_ASAP7_75t_SL g14494 ( 
.A(n_14428),
.B(n_5884),
.Y(n_14494)
);

NAND4xp75_ASAP7_75t_L g14495 ( 
.A(n_14345),
.B(n_6404),
.C(n_6421),
.D(n_6372),
.Y(n_14495)
);

AND2x4_ASAP7_75t_L g14496 ( 
.A(n_14412),
.B(n_5858),
.Y(n_14496)
);

INVx1_ASAP7_75t_L g14497 ( 
.A(n_14372),
.Y(n_14497)
);

NOR2x1_ASAP7_75t_L g14498 ( 
.A(n_14355),
.B(n_5762),
.Y(n_14498)
);

NOR2x1_ASAP7_75t_L g14499 ( 
.A(n_14420),
.B(n_5764),
.Y(n_14499)
);

NAND2xp5_ASAP7_75t_SL g14500 ( 
.A(n_14391),
.B(n_5884),
.Y(n_14500)
);

NOR2x1_ASAP7_75t_L g14501 ( 
.A(n_14359),
.B(n_5764),
.Y(n_14501)
);

NOR2x1_ASAP7_75t_L g14502 ( 
.A(n_14389),
.B(n_5771),
.Y(n_14502)
);

AOI211xp5_ASAP7_75t_L g14503 ( 
.A1(n_14438),
.A2(n_14414),
.B(n_14416),
.C(n_14417),
.Y(n_14503)
);

NOR3xp33_ASAP7_75t_L g14504 ( 
.A(n_14435),
.B(n_14425),
.C(n_14354),
.Y(n_14504)
);

NAND5xp2_ASAP7_75t_L g14505 ( 
.A(n_14449),
.B(n_14347),
.C(n_14429),
.D(n_14360),
.E(n_4420),
.Y(n_14505)
);

AND2x2_ASAP7_75t_L g14506 ( 
.A(n_14433),
.B(n_7193),
.Y(n_14506)
);

NAND3xp33_ASAP7_75t_L g14507 ( 
.A(n_14446),
.B(n_5591),
.C(n_5571),
.Y(n_14507)
);

XOR2xp5_ASAP7_75t_L g14508 ( 
.A(n_14452),
.B(n_5546),
.Y(n_14508)
);

AND2x4_ASAP7_75t_L g14509 ( 
.A(n_14456),
.B(n_5858),
.Y(n_14509)
);

NAND5xp2_ASAP7_75t_L g14510 ( 
.A(n_14454),
.B(n_5317),
.C(n_4708),
.D(n_5625),
.E(n_5586),
.Y(n_14510)
);

NAND3xp33_ASAP7_75t_L g14511 ( 
.A(n_14450),
.B(n_5591),
.C(n_5571),
.Y(n_14511)
);

INVx1_ASAP7_75t_L g14512 ( 
.A(n_14439),
.Y(n_14512)
);

NAND4xp75_ASAP7_75t_L g14513 ( 
.A(n_14458),
.B(n_6147),
.C(n_6150),
.D(n_6141),
.Y(n_14513)
);

AOI211xp5_ASAP7_75t_L g14514 ( 
.A1(n_14479),
.A2(n_4616),
.B(n_6819),
.C(n_6996),
.Y(n_14514)
);

NAND4xp25_ASAP7_75t_L g14515 ( 
.A(n_14482),
.B(n_5794),
.C(n_5820),
.D(n_5771),
.Y(n_14515)
);

NAND4xp25_ASAP7_75t_L g14516 ( 
.A(n_14436),
.B(n_5794),
.C(n_5820),
.D(n_5771),
.Y(n_14516)
);

AOI211xp5_ASAP7_75t_L g14517 ( 
.A1(n_14477),
.A2(n_4616),
.B(n_6842),
.C(n_6898),
.Y(n_14517)
);

AND2x4_ASAP7_75t_L g14518 ( 
.A(n_14475),
.B(n_5858),
.Y(n_14518)
);

O2A1O1Ixp33_ASAP7_75t_L g14519 ( 
.A1(n_14497),
.A2(n_14466),
.B(n_14500),
.C(n_14432),
.Y(n_14519)
);

AOI211xp5_ASAP7_75t_L g14520 ( 
.A1(n_14451),
.A2(n_6842),
.B(n_6903),
.C(n_6901),
.Y(n_14520)
);

AOI31xp33_ASAP7_75t_L g14521 ( 
.A1(n_14502),
.A2(n_6390),
.A3(n_6395),
.B(n_6384),
.Y(n_14521)
);

NOR3xp33_ASAP7_75t_L g14522 ( 
.A(n_14472),
.B(n_6671),
.C(n_6670),
.Y(n_14522)
);

OAI211xp5_ASAP7_75t_L g14523 ( 
.A1(n_14467),
.A2(n_5924),
.B(n_5926),
.C(n_4850),
.Y(n_14523)
);

NAND2xp5_ASAP7_75t_L g14524 ( 
.A(n_14457),
.B(n_7342),
.Y(n_14524)
);

NAND4xp25_ASAP7_75t_L g14525 ( 
.A(n_14453),
.B(n_5794),
.C(n_5820),
.D(n_5771),
.Y(n_14525)
);

OAI211xp5_ASAP7_75t_SL g14526 ( 
.A1(n_14480),
.A2(n_6040),
.B(n_6041),
.C(n_6021),
.Y(n_14526)
);

O2A1O1Ixp33_ASAP7_75t_L g14527 ( 
.A1(n_14440),
.A2(n_5820),
.B(n_5827),
.C(n_5794),
.Y(n_14527)
);

NAND3xp33_ASAP7_75t_L g14528 ( 
.A(n_14437),
.B(n_5591),
.C(n_5571),
.Y(n_14528)
);

AOI221xp5_ASAP7_75t_L g14529 ( 
.A1(n_14444),
.A2(n_5604),
.B1(n_5609),
.B2(n_5591),
.C(n_5571),
.Y(n_14529)
);

NAND4xp25_ASAP7_75t_L g14530 ( 
.A(n_14445),
.B(n_5844),
.C(n_5860),
.D(n_5827),
.Y(n_14530)
);

OAI211xp5_ASAP7_75t_SL g14531 ( 
.A1(n_14498),
.A2(n_6041),
.B(n_6066),
.C(n_6040),
.Y(n_14531)
);

OAI221xp5_ASAP7_75t_SL g14532 ( 
.A1(n_14461),
.A2(n_5860),
.B1(n_5869),
.B2(n_5844),
.C(n_5827),
.Y(n_14532)
);

OAI221xp5_ASAP7_75t_L g14533 ( 
.A1(n_14473),
.A2(n_6429),
.B1(n_6395),
.B2(n_6035),
.C(n_6043),
.Y(n_14533)
);

OAI221xp5_ASAP7_75t_L g14534 ( 
.A1(n_14492),
.A2(n_6429),
.B1(n_6035),
.B2(n_6043),
.C(n_6026),
.Y(n_14534)
);

NAND4xp25_ASAP7_75t_L g14535 ( 
.A(n_14490),
.B(n_5844),
.C(n_5860),
.D(n_5827),
.Y(n_14535)
);

OAI211xp5_ASAP7_75t_SL g14536 ( 
.A1(n_14494),
.A2(n_6041),
.B(n_6066),
.C(n_6040),
.Y(n_14536)
);

OAI211xp5_ASAP7_75t_SL g14537 ( 
.A1(n_14499),
.A2(n_14501),
.B(n_14474),
.C(n_14465),
.Y(n_14537)
);

OAI211xp5_ASAP7_75t_SL g14538 ( 
.A1(n_14478),
.A2(n_6066),
.B(n_6102),
.C(n_6041),
.Y(n_14538)
);

AND2x4_ASAP7_75t_L g14539 ( 
.A(n_14462),
.B(n_7359),
.Y(n_14539)
);

AOI221x1_ASAP7_75t_L g14540 ( 
.A1(n_14463),
.A2(n_5565),
.B1(n_5580),
.B2(n_5561),
.C(n_5558),
.Y(n_14540)
);

NAND3xp33_ASAP7_75t_SL g14541 ( 
.A(n_14485),
.B(n_6147),
.C(n_6141),
.Y(n_14541)
);

NAND2xp5_ASAP7_75t_L g14542 ( 
.A(n_14462),
.B(n_7342),
.Y(n_14542)
);

NAND2xp5_ASAP7_75t_L g14543 ( 
.A(n_14489),
.B(n_7342),
.Y(n_14543)
);

NOR3xp33_ASAP7_75t_SL g14544 ( 
.A(n_14484),
.B(n_7342),
.C(n_5365),
.Y(n_14544)
);

NAND2xp5_ASAP7_75t_L g14545 ( 
.A(n_14443),
.B(n_7342),
.Y(n_14545)
);

NOR2xp33_ASAP7_75t_R g14546 ( 
.A(n_14488),
.B(n_6181),
.Y(n_14546)
);

INVx1_ASAP7_75t_L g14547 ( 
.A(n_14491),
.Y(n_14547)
);

INVx1_ASAP7_75t_L g14548 ( 
.A(n_14495),
.Y(n_14548)
);

OA211x2_ASAP7_75t_L g14549 ( 
.A1(n_14464),
.A2(n_7342),
.B(n_7379),
.C(n_7258),
.Y(n_14549)
);

AOI211x1_ASAP7_75t_L g14550 ( 
.A1(n_14455),
.A2(n_6076),
.B(n_6093),
.C(n_6141),
.Y(n_14550)
);

AOI21xp5_ASAP7_75t_L g14551 ( 
.A1(n_14469),
.A2(n_6903),
.B(n_6901),
.Y(n_14551)
);

NOR2xp33_ASAP7_75t_L g14552 ( 
.A(n_14496),
.B(n_14459),
.Y(n_14552)
);

A2O1A1Ixp33_ASAP7_75t_L g14553 ( 
.A1(n_14496),
.A2(n_7206),
.B(n_7220),
.C(n_7201),
.Y(n_14553)
);

NOR3xp33_ASAP7_75t_L g14554 ( 
.A(n_14460),
.B(n_6671),
.C(n_6670),
.Y(n_14554)
);

NOR4xp25_ASAP7_75t_L g14555 ( 
.A(n_14481),
.B(n_6026),
.C(n_6035),
.D(n_6002),
.Y(n_14555)
);

NOR4xp25_ASAP7_75t_L g14556 ( 
.A(n_14486),
.B(n_6026),
.C(n_6043),
.D(n_6002),
.Y(n_14556)
);

NOR3xp33_ASAP7_75t_L g14557 ( 
.A(n_14493),
.B(n_14471),
.C(n_14448),
.Y(n_14557)
);

OAI211xp5_ASAP7_75t_SL g14558 ( 
.A1(n_14468),
.A2(n_6066),
.B(n_6102),
.C(n_6041),
.Y(n_14558)
);

NAND2xp5_ASAP7_75t_L g14559 ( 
.A(n_14442),
.B(n_7342),
.Y(n_14559)
);

OAI221xp5_ASAP7_75t_SL g14560 ( 
.A1(n_14487),
.A2(n_5869),
.B1(n_5872),
.B2(n_5860),
.C(n_5844),
.Y(n_14560)
);

AOI221x1_ASAP7_75t_L g14561 ( 
.A1(n_14447),
.A2(n_5565),
.B1(n_5580),
.B2(n_5561),
.C(n_5558),
.Y(n_14561)
);

AND2x4_ASAP7_75t_L g14562 ( 
.A(n_14509),
.B(n_14476),
.Y(n_14562)
);

INVx2_ASAP7_75t_L g14563 ( 
.A(n_14547),
.Y(n_14563)
);

INVx2_ASAP7_75t_L g14564 ( 
.A(n_14512),
.Y(n_14564)
);

NAND2xp33_ASAP7_75t_SL g14565 ( 
.A(n_14548),
.B(n_14447),
.Y(n_14565)
);

NOR2xp33_ASAP7_75t_L g14566 ( 
.A(n_14537),
.B(n_14431),
.Y(n_14566)
);

NOR3xp33_ASAP7_75t_L g14567 ( 
.A(n_14519),
.B(n_14470),
.C(n_14483),
.Y(n_14567)
);

NAND2xp5_ASAP7_75t_SL g14568 ( 
.A(n_14504),
.B(n_14434),
.Y(n_14568)
);

INVx1_ASAP7_75t_L g14569 ( 
.A(n_14552),
.Y(n_14569)
);

NAND4xp75_ASAP7_75t_L g14570 ( 
.A(n_14543),
.B(n_14441),
.C(n_6058),
.D(n_6052),
.Y(n_14570)
);

OAI211xp5_ASAP7_75t_L g14571 ( 
.A1(n_14503),
.A2(n_14441),
.B(n_5924),
.C(n_5926),
.Y(n_14571)
);

NAND3xp33_ASAP7_75t_L g14572 ( 
.A(n_14557),
.B(n_5926),
.C(n_5924),
.Y(n_14572)
);

INVx1_ASAP7_75t_L g14573 ( 
.A(n_14508),
.Y(n_14573)
);

NOR2x1_ASAP7_75t_L g14574 ( 
.A(n_14525),
.B(n_14505),
.Y(n_14574)
);

AND2x2_ASAP7_75t_L g14575 ( 
.A(n_14509),
.B(n_14518),
.Y(n_14575)
);

NAND4xp75_ASAP7_75t_L g14576 ( 
.A(n_14559),
.B(n_6058),
.C(n_6052),
.D(n_6147),
.Y(n_14576)
);

NAND2xp5_ASAP7_75t_L g14577 ( 
.A(n_14518),
.B(n_7193),
.Y(n_14577)
);

NOR2xp67_ASAP7_75t_L g14578 ( 
.A(n_14507),
.B(n_5924),
.Y(n_14578)
);

AO22x1_ASAP7_75t_L g14579 ( 
.A1(n_14522),
.A2(n_14554),
.B1(n_14524),
.B2(n_14506),
.Y(n_14579)
);

OR2x2_ASAP7_75t_L g14580 ( 
.A(n_14545),
.B(n_7193),
.Y(n_14580)
);

INVxp67_ASAP7_75t_L g14581 ( 
.A(n_14511),
.Y(n_14581)
);

INVx1_ASAP7_75t_L g14582 ( 
.A(n_14526),
.Y(n_14582)
);

OR2x2_ASAP7_75t_L g14583 ( 
.A(n_14541),
.B(n_7193),
.Y(n_14583)
);

AND2x2_ASAP7_75t_L g14584 ( 
.A(n_14544),
.B(n_6797),
.Y(n_14584)
);

OR2x2_ASAP7_75t_L g14585 ( 
.A(n_14528),
.B(n_7193),
.Y(n_14585)
);

INVx1_ASAP7_75t_L g14586 ( 
.A(n_14546),
.Y(n_14586)
);

NOR2x1_ASAP7_75t_L g14587 ( 
.A(n_14531),
.B(n_5869),
.Y(n_14587)
);

INVx2_ASAP7_75t_L g14588 ( 
.A(n_14542),
.Y(n_14588)
);

AND2x2_ASAP7_75t_L g14589 ( 
.A(n_14556),
.B(n_6797),
.Y(n_14589)
);

NAND4xp75_ASAP7_75t_L g14590 ( 
.A(n_14549),
.B(n_6058),
.C(n_6052),
.D(n_6150),
.Y(n_14590)
);

OAI21xp5_ASAP7_75t_SL g14591 ( 
.A1(n_14521),
.A2(n_14523),
.B(n_14535),
.Y(n_14591)
);

OAI21xp5_ASAP7_75t_L g14592 ( 
.A1(n_14555),
.A2(n_6675),
.B(n_6671),
.Y(n_14592)
);

NAND4xp75_ASAP7_75t_L g14593 ( 
.A(n_14550),
.B(n_6150),
.C(n_6172),
.D(n_6094),
.Y(n_14593)
);

INVx2_ASAP7_75t_L g14594 ( 
.A(n_14534),
.Y(n_14594)
);

AND2x4_ASAP7_75t_L g14595 ( 
.A(n_14540),
.B(n_5717),
.Y(n_14595)
);

NOR4xp25_ASAP7_75t_L g14596 ( 
.A(n_14536),
.B(n_6102),
.C(n_6168),
.D(n_6066),
.Y(n_14596)
);

NOR3xp33_ASAP7_75t_L g14597 ( 
.A(n_14538),
.B(n_4622),
.C(n_4608),
.Y(n_14597)
);

AOI22xp5_ASAP7_75t_L g14598 ( 
.A1(n_14530),
.A2(n_5591),
.B1(n_5604),
.B2(n_5571),
.Y(n_14598)
);

OAI221xp5_ASAP7_75t_L g14599 ( 
.A1(n_14532),
.A2(n_4708),
.B1(n_5317),
.B2(n_5872),
.C(n_5869),
.Y(n_14599)
);

INVx1_ASAP7_75t_L g14600 ( 
.A(n_14527),
.Y(n_14600)
);

AOI22xp5_ASAP7_75t_L g14601 ( 
.A1(n_14516),
.A2(n_5591),
.B1(n_5604),
.B2(n_5571),
.Y(n_14601)
);

INVx2_ASAP7_75t_L g14602 ( 
.A(n_14533),
.Y(n_14602)
);

INVx1_ASAP7_75t_L g14603 ( 
.A(n_14561),
.Y(n_14603)
);

INVx1_ASAP7_75t_L g14604 ( 
.A(n_14510),
.Y(n_14604)
);

INVx3_ASAP7_75t_L g14605 ( 
.A(n_14513),
.Y(n_14605)
);

NOR2xp67_ASAP7_75t_L g14606 ( 
.A(n_14515),
.B(n_5924),
.Y(n_14606)
);

INVx1_ASAP7_75t_L g14607 ( 
.A(n_14558),
.Y(n_14607)
);

INVx1_ASAP7_75t_L g14608 ( 
.A(n_14560),
.Y(n_14608)
);

NOR4xp75_ASAP7_75t_L g14609 ( 
.A(n_14568),
.B(n_14551),
.C(n_14517),
.D(n_14520),
.Y(n_14609)
);

AOI21x1_ASAP7_75t_L g14610 ( 
.A1(n_14569),
.A2(n_14539),
.B(n_14514),
.Y(n_14610)
);

NOR3xp33_ASAP7_75t_L g14611 ( 
.A(n_14564),
.B(n_14529),
.C(n_14539),
.Y(n_14611)
);

OR3x1_ASAP7_75t_L g14612 ( 
.A(n_14566),
.B(n_14553),
.C(n_5368),
.Y(n_14612)
);

AO211x2_ASAP7_75t_L g14613 ( 
.A1(n_14567),
.A2(n_14573),
.B(n_14604),
.C(n_14600),
.Y(n_14613)
);

AOI22xp5_ASAP7_75t_L g14614 ( 
.A1(n_14563),
.A2(n_5865),
.B1(n_6029),
.B2(n_5639),
.Y(n_14614)
);

NOR5xp2_ASAP7_75t_L g14615 ( 
.A(n_14581),
.B(n_4993),
.C(n_5036),
.D(n_5022),
.E(n_5016),
.Y(n_14615)
);

XNOR2xp5_ASAP7_75t_L g14616 ( 
.A(n_14575),
.B(n_6943),
.Y(n_14616)
);

NAND3xp33_ASAP7_75t_SL g14617 ( 
.A(n_14565),
.B(n_14588),
.C(n_14586),
.Y(n_14617)
);

NAND4xp75_ASAP7_75t_L g14618 ( 
.A(n_14574),
.B(n_6172),
.C(n_6093),
.D(n_6076),
.Y(n_14618)
);

AND2x4_ASAP7_75t_L g14619 ( 
.A(n_14562),
.B(n_7193),
.Y(n_14619)
);

AOI21xp5_ASAP7_75t_L g14620 ( 
.A1(n_14608),
.A2(n_5891),
.B(n_5622),
.Y(n_14620)
);

AND5x1_ASAP7_75t_L g14621 ( 
.A(n_14579),
.B(n_7258),
.C(n_7379),
.D(n_7096),
.E(n_7251),
.Y(n_14621)
);

NAND4xp75_ASAP7_75t_L g14622 ( 
.A(n_14603),
.B(n_6172),
.C(n_6093),
.D(n_6076),
.Y(n_14622)
);

OR5x1_ASAP7_75t_L g14623 ( 
.A(n_14571),
.B(n_7258),
.C(n_7379),
.D(n_6932),
.E(n_6939),
.Y(n_14623)
);

XNOR2xp5_ASAP7_75t_L g14624 ( 
.A(n_14605),
.B(n_6943),
.Y(n_14624)
);

NAND5xp2_ASAP7_75t_L g14625 ( 
.A(n_14591),
.B(n_5317),
.C(n_4708),
.D(n_4506),
.E(n_4520),
.Y(n_14625)
);

AND2x2_ASAP7_75t_SL g14626 ( 
.A(n_14594),
.B(n_4955),
.Y(n_14626)
);

NOR3xp33_ASAP7_75t_L g14627 ( 
.A(n_14602),
.B(n_6903),
.C(n_6901),
.Y(n_14627)
);

NAND4xp25_ASAP7_75t_SL g14628 ( 
.A(n_14582),
.B(n_6094),
.C(n_6261),
.D(n_6259),
.Y(n_14628)
);

NAND3xp33_ASAP7_75t_L g14629 ( 
.A(n_14607),
.B(n_5926),
.C(n_5924),
.Y(n_14629)
);

NAND3xp33_ASAP7_75t_L g14630 ( 
.A(n_14606),
.B(n_5926),
.C(n_5924),
.Y(n_14630)
);

AO211x2_ASAP7_75t_L g14631 ( 
.A1(n_14577),
.A2(n_5368),
.B(n_5374),
.C(n_5361),
.Y(n_14631)
);

NAND2xp5_ASAP7_75t_L g14632 ( 
.A(n_14570),
.B(n_7258),
.Y(n_14632)
);

NAND4xp25_ASAP7_75t_L g14633 ( 
.A(n_14584),
.B(n_5885),
.C(n_5886),
.D(n_5872),
.Y(n_14633)
);

AND2x2_ASAP7_75t_L g14634 ( 
.A(n_14589),
.B(n_6943),
.Y(n_14634)
);

XNOR2x1_ASAP7_75t_L g14635 ( 
.A(n_14590),
.B(n_6943),
.Y(n_14635)
);

NOR4xp25_ASAP7_75t_L g14636 ( 
.A(n_14580),
.B(n_6168),
.C(n_6204),
.D(n_6102),
.Y(n_14636)
);

NAND3xp33_ASAP7_75t_L g14637 ( 
.A(n_14578),
.B(n_5926),
.C(n_5924),
.Y(n_14637)
);

OAI211xp5_ASAP7_75t_SL g14638 ( 
.A1(n_14583),
.A2(n_6102),
.B(n_6204),
.C(n_6168),
.Y(n_14638)
);

NOR3xp33_ASAP7_75t_SL g14639 ( 
.A(n_14576),
.B(n_5377),
.C(n_5374),
.Y(n_14639)
);

OR4x2_ASAP7_75t_L g14640 ( 
.A(n_14587),
.B(n_7258),
.C(n_7379),
.D(n_6181),
.Y(n_14640)
);

NOR3xp33_ASAP7_75t_L g14641 ( 
.A(n_14593),
.B(n_6922),
.C(n_6920),
.Y(n_14641)
);

AND2x4_ASAP7_75t_L g14642 ( 
.A(n_14595),
.B(n_7258),
.Y(n_14642)
);

NOR3xp33_ASAP7_75t_SL g14643 ( 
.A(n_14572),
.B(n_5383),
.C(n_5377),
.Y(n_14643)
);

NOR4xp25_ASAP7_75t_L g14644 ( 
.A(n_14585),
.B(n_6204),
.C(n_6215),
.D(n_6168),
.Y(n_14644)
);

INVx1_ASAP7_75t_L g14645 ( 
.A(n_14597),
.Y(n_14645)
);

OAI211xp5_ASAP7_75t_L g14646 ( 
.A1(n_14596),
.A2(n_5924),
.B(n_5926),
.C(n_4850),
.Y(n_14646)
);

NAND3xp33_ASAP7_75t_SL g14647 ( 
.A(n_14592),
.B(n_4622),
.C(n_4608),
.Y(n_14647)
);

NOR3xp33_ASAP7_75t_L g14648 ( 
.A(n_14599),
.B(n_6922),
.C(n_6920),
.Y(n_14648)
);

NAND4xp25_ASAP7_75t_L g14649 ( 
.A(n_14598),
.B(n_14601),
.C(n_5885),
.D(n_5886),
.Y(n_14649)
);

NOR4xp25_ASAP7_75t_L g14650 ( 
.A(n_14569),
.B(n_6204),
.C(n_6215),
.D(n_6168),
.Y(n_14650)
);

OR2x2_ASAP7_75t_L g14651 ( 
.A(n_14563),
.B(n_7258),
.Y(n_14651)
);

NOR3xp33_ASAP7_75t_L g14652 ( 
.A(n_14569),
.B(n_6922),
.C(n_6920),
.Y(n_14652)
);

NAND4xp25_ASAP7_75t_L g14653 ( 
.A(n_14574),
.B(n_5885),
.C(n_5886),
.D(n_5872),
.Y(n_14653)
);

NOR2x1_ASAP7_75t_L g14654 ( 
.A(n_14563),
.B(n_5885),
.Y(n_14654)
);

INVx1_ASAP7_75t_L g14655 ( 
.A(n_14613),
.Y(n_14655)
);

HB1xp67_ASAP7_75t_L g14656 ( 
.A(n_14617),
.Y(n_14656)
);

NAND3xp33_ASAP7_75t_SL g14657 ( 
.A(n_14611),
.B(n_4622),
.C(n_4608),
.Y(n_14657)
);

OAI311xp33_ASAP7_75t_L g14658 ( 
.A1(n_14645),
.A2(n_6223),
.A3(n_6252),
.B1(n_6215),
.C1(n_6204),
.Y(n_14658)
);

OAI222xp33_ASAP7_75t_R g14659 ( 
.A1(n_14610),
.A2(n_4891),
.B1(n_4872),
.B2(n_4901),
.C1(n_4885),
.C2(n_4859),
.Y(n_14659)
);

NOR3xp33_ASAP7_75t_L g14660 ( 
.A(n_14638),
.B(n_4622),
.C(n_4608),
.Y(n_14660)
);

OAI221xp5_ASAP7_75t_L g14661 ( 
.A1(n_14654),
.A2(n_5317),
.B1(n_5926),
.B2(n_5886),
.C(n_5891),
.Y(n_14661)
);

NAND3xp33_ASAP7_75t_L g14662 ( 
.A(n_14634),
.B(n_5926),
.C(n_5591),
.Y(n_14662)
);

AOI221xp5_ASAP7_75t_L g14663 ( 
.A1(n_14644),
.A2(n_5604),
.B1(n_5609),
.B2(n_5591),
.C(n_5571),
.Y(n_14663)
);

NOR3xp33_ASAP7_75t_L g14664 ( 
.A(n_14647),
.B(n_4622),
.C(n_4608),
.Y(n_14664)
);

OAI22xp5_ASAP7_75t_SL g14665 ( 
.A1(n_14626),
.A2(n_5317),
.B1(n_7055),
.B2(n_6943),
.Y(n_14665)
);

AOI211xp5_ASAP7_75t_L g14666 ( 
.A1(n_14636),
.A2(n_5604),
.B(n_5609),
.C(n_5571),
.Y(n_14666)
);

AOI22xp5_ASAP7_75t_L g14667 ( 
.A1(n_14624),
.A2(n_5317),
.B1(n_5609),
.B2(n_5604),
.Y(n_14667)
);

NOR2x1_ASAP7_75t_L g14668 ( 
.A(n_14612),
.B(n_7143),
.Y(n_14668)
);

INVx1_ASAP7_75t_L g14669 ( 
.A(n_14609),
.Y(n_14669)
);

AOI221xp5_ASAP7_75t_L g14670 ( 
.A1(n_14632),
.A2(n_5614),
.B1(n_5635),
.B2(n_5609),
.C(n_5604),
.Y(n_14670)
);

OAI221xp5_ASAP7_75t_L g14671 ( 
.A1(n_14616),
.A2(n_5891),
.B1(n_6212),
.B2(n_5958),
.C(n_5622),
.Y(n_14671)
);

NAND5xp2_ASAP7_75t_L g14672 ( 
.A(n_14620),
.B(n_4506),
.C(n_4520),
.D(n_4507),
.E(n_4497),
.Y(n_14672)
);

AOI21xp5_ASAP7_75t_L g14673 ( 
.A1(n_14635),
.A2(n_5891),
.B(n_5622),
.Y(n_14673)
);

NAND2xp5_ASAP7_75t_L g14674 ( 
.A(n_14631),
.B(n_7055),
.Y(n_14674)
);

NOR2xp67_ASAP7_75t_L g14675 ( 
.A(n_14649),
.B(n_14630),
.Y(n_14675)
);

AND4x1_ASAP7_75t_L g14676 ( 
.A(n_14639),
.B(n_5856),
.C(n_5851),
.D(n_5647),
.Y(n_14676)
);

INVx2_ASAP7_75t_L g14677 ( 
.A(n_14651),
.Y(n_14677)
);

NOR2xp33_ASAP7_75t_L g14678 ( 
.A(n_14637),
.B(n_7055),
.Y(n_14678)
);

AND2x4_ASAP7_75t_L g14679 ( 
.A(n_14643),
.B(n_7096),
.Y(n_14679)
);

NAND3xp33_ASAP7_75t_SL g14680 ( 
.A(n_14641),
.B(n_14648),
.C(n_14614),
.Y(n_14680)
);

HB1xp67_ASAP7_75t_L g14681 ( 
.A(n_14633),
.Y(n_14681)
);

INVx1_ASAP7_75t_L g14682 ( 
.A(n_14646),
.Y(n_14682)
);

INVxp67_ASAP7_75t_SL g14683 ( 
.A(n_14615),
.Y(n_14683)
);

NAND3xp33_ASAP7_75t_SL g14684 ( 
.A(n_14650),
.B(n_4637),
.C(n_4058),
.Y(n_14684)
);

NAND3xp33_ASAP7_75t_SL g14685 ( 
.A(n_14627),
.B(n_4637),
.C(n_4058),
.Y(n_14685)
);

INVxp67_ASAP7_75t_L g14686 ( 
.A(n_14625),
.Y(n_14686)
);

NOR5xp2_ASAP7_75t_L g14687 ( 
.A(n_14629),
.B(n_5392),
.C(n_5397),
.D(n_5387),
.E(n_5383),
.Y(n_14687)
);

OAI221xp5_ASAP7_75t_R g14688 ( 
.A1(n_14652),
.A2(n_6087),
.B1(n_5995),
.B2(n_7379),
.C(n_6924),
.Y(n_14688)
);

AOI21xp5_ASAP7_75t_L g14689 ( 
.A1(n_14642),
.A2(n_5891),
.B(n_5622),
.Y(n_14689)
);

AOI221xp5_ASAP7_75t_L g14690 ( 
.A1(n_14640),
.A2(n_14642),
.B1(n_14653),
.B2(n_14628),
.C(n_14619),
.Y(n_14690)
);

INVx1_ASAP7_75t_L g14691 ( 
.A(n_14618),
.Y(n_14691)
);

NAND5xp2_ASAP7_75t_L g14692 ( 
.A(n_14655),
.B(n_14623),
.C(n_14621),
.D(n_14622),
.E(n_14619),
.Y(n_14692)
);

INVx1_ASAP7_75t_L g14693 ( 
.A(n_14656),
.Y(n_14693)
);

INVx1_ASAP7_75t_L g14694 ( 
.A(n_14669),
.Y(n_14694)
);

HB1xp67_ASAP7_75t_L g14695 ( 
.A(n_14677),
.Y(n_14695)
);

OA22x2_ASAP7_75t_L g14696 ( 
.A1(n_14686),
.A2(n_6923),
.B1(n_6932),
.B2(n_6924),
.Y(n_14696)
);

NAND2xp5_ASAP7_75t_SL g14697 ( 
.A(n_14691),
.B(n_5604),
.Y(n_14697)
);

INVx2_ASAP7_75t_L g14698 ( 
.A(n_14681),
.Y(n_14698)
);

NAND3xp33_ASAP7_75t_L g14699 ( 
.A(n_14690),
.B(n_5614),
.C(n_5609),
.Y(n_14699)
);

AOI22xp5_ASAP7_75t_SL g14700 ( 
.A1(n_14683),
.A2(n_4660),
.B1(n_5375),
.B2(n_5044),
.Y(n_14700)
);

NAND2xp5_ASAP7_75t_L g14701 ( 
.A(n_14675),
.B(n_7379),
.Y(n_14701)
);

INVx2_ASAP7_75t_L g14702 ( 
.A(n_14682),
.Y(n_14702)
);

INVx1_ASAP7_75t_SL g14703 ( 
.A(n_14668),
.Y(n_14703)
);

OAI22xp5_ASAP7_75t_L g14704 ( 
.A1(n_14674),
.A2(n_5609),
.B1(n_5635),
.B2(n_5614),
.Y(n_14704)
);

INVx2_ASAP7_75t_L g14705 ( 
.A(n_14679),
.Y(n_14705)
);

OAI221xp5_ASAP7_75t_L g14706 ( 
.A1(n_14680),
.A2(n_5958),
.B1(n_6212),
.B2(n_5622),
.C(n_4660),
.Y(n_14706)
);

AND2x2_ASAP7_75t_L g14707 ( 
.A(n_14678),
.B(n_7055),
.Y(n_14707)
);

XNOR2x1_ASAP7_75t_L g14708 ( 
.A(n_14679),
.B(n_7055),
.Y(n_14708)
);

AOI22xp5_ASAP7_75t_L g14709 ( 
.A1(n_14685),
.A2(n_5614),
.B1(n_5635),
.B2(n_5609),
.Y(n_14709)
);

A2O1A1Ixp33_ASAP7_75t_L g14710 ( 
.A1(n_14664),
.A2(n_6923),
.B(n_6932),
.C(n_6924),
.Y(n_14710)
);

INVx1_ASAP7_75t_L g14711 ( 
.A(n_14684),
.Y(n_14711)
);

AO22x2_ASAP7_75t_L g14712 ( 
.A1(n_14657),
.A2(n_5546),
.B1(n_5606),
.B2(n_5596),
.Y(n_14712)
);

AOI22xp5_ASAP7_75t_L g14713 ( 
.A1(n_14660),
.A2(n_5635),
.B1(n_5639),
.B2(n_5614),
.Y(n_14713)
);

INVx1_ASAP7_75t_L g14714 ( 
.A(n_14662),
.Y(n_14714)
);

INVx1_ASAP7_75t_L g14715 ( 
.A(n_14676),
.Y(n_14715)
);

XNOR2x1_ASAP7_75t_L g14716 ( 
.A(n_14667),
.B(n_6675),
.Y(n_14716)
);

OAI21xp33_ASAP7_75t_L g14717 ( 
.A1(n_14673),
.A2(n_6223),
.B(n_6215),
.Y(n_14717)
);

INVx1_ASAP7_75t_L g14718 ( 
.A(n_14672),
.Y(n_14718)
);

INVx2_ASAP7_75t_SL g14719 ( 
.A(n_14659),
.Y(n_14719)
);

OAI221xp5_ASAP7_75t_L g14720 ( 
.A1(n_14689),
.A2(n_6212),
.B1(n_5958),
.B2(n_4660),
.C(n_5025),
.Y(n_14720)
);

NAND3xp33_ASAP7_75t_SL g14721 ( 
.A(n_14687),
.B(n_4637),
.C(n_4058),
.Y(n_14721)
);

NAND2xp5_ASAP7_75t_L g14722 ( 
.A(n_14666),
.B(n_7379),
.Y(n_14722)
);

NAND2xp5_ASAP7_75t_L g14723 ( 
.A(n_14670),
.B(n_14665),
.Y(n_14723)
);

NAND4xp75_ASAP7_75t_L g14724 ( 
.A(n_14688),
.B(n_4885),
.C(n_4891),
.D(n_4872),
.Y(n_14724)
);

OAI22xp5_ASAP7_75t_L g14725 ( 
.A1(n_14693),
.A2(n_14661),
.B1(n_14663),
.B2(n_14671),
.Y(n_14725)
);

HB1xp67_ASAP7_75t_L g14726 ( 
.A(n_14695),
.Y(n_14726)
);

NOR2x1_ASAP7_75t_L g14727 ( 
.A(n_14694),
.B(n_14658),
.Y(n_14727)
);

INVx1_ASAP7_75t_L g14728 ( 
.A(n_14698),
.Y(n_14728)
);

INVx2_ASAP7_75t_L g14729 ( 
.A(n_14702),
.Y(n_14729)
);

AOI22xp5_ASAP7_75t_L g14730 ( 
.A1(n_14718),
.A2(n_5614),
.B1(n_5639),
.B2(n_5635),
.Y(n_14730)
);

AOI22xp5_ASAP7_75t_L g14731 ( 
.A1(n_14715),
.A2(n_5614),
.B1(n_5639),
.B2(n_5635),
.Y(n_14731)
);

INVx1_ASAP7_75t_L g14732 ( 
.A(n_14705),
.Y(n_14732)
);

INVx1_ASAP7_75t_L g14733 ( 
.A(n_14703),
.Y(n_14733)
);

INVxp67_ASAP7_75t_L g14734 ( 
.A(n_14714),
.Y(n_14734)
);

XOR2xp5_ASAP7_75t_L g14735 ( 
.A(n_14711),
.B(n_5614),
.Y(n_14735)
);

OAI22xp5_ASAP7_75t_L g14736 ( 
.A1(n_14719),
.A2(n_5639),
.B1(n_5667),
.B2(n_5635),
.Y(n_14736)
);

OAI22xp5_ASAP7_75t_SL g14737 ( 
.A1(n_14723),
.A2(n_5950),
.B1(n_6003),
.B2(n_5998),
.Y(n_14737)
);

INVx1_ASAP7_75t_L g14738 ( 
.A(n_14692),
.Y(n_14738)
);

XOR2xp5_ASAP7_75t_L g14739 ( 
.A(n_14697),
.B(n_5635),
.Y(n_14739)
);

INVx1_ASAP7_75t_L g14740 ( 
.A(n_14716),
.Y(n_14740)
);

INVx1_ASAP7_75t_L g14741 ( 
.A(n_14701),
.Y(n_14741)
);

AOI22xp5_ASAP7_75t_L g14742 ( 
.A1(n_14699),
.A2(n_5639),
.B1(n_5691),
.B2(n_5667),
.Y(n_14742)
);

INVx2_ASAP7_75t_L g14743 ( 
.A(n_14724),
.Y(n_14743)
);

INVx1_ASAP7_75t_L g14744 ( 
.A(n_14722),
.Y(n_14744)
);

INVx1_ASAP7_75t_L g14745 ( 
.A(n_14726),
.Y(n_14745)
);

HB1xp67_ASAP7_75t_L g14746 ( 
.A(n_14728),
.Y(n_14746)
);

INVx1_ASAP7_75t_L g14747 ( 
.A(n_14729),
.Y(n_14747)
);

NAND2xp33_ASAP7_75t_L g14748 ( 
.A(n_14733),
.B(n_14717),
.Y(n_14748)
);

NAND2xp5_ASAP7_75t_L g14749 ( 
.A(n_14738),
.B(n_14708),
.Y(n_14749)
);

OR3x1_ASAP7_75t_L g14750 ( 
.A(n_14732),
.B(n_14721),
.C(n_14712),
.Y(n_14750)
);

INVx1_ASAP7_75t_L g14751 ( 
.A(n_14734),
.Y(n_14751)
);

AOI21xp5_ASAP7_75t_L g14752 ( 
.A1(n_14727),
.A2(n_14712),
.B(n_14704),
.Y(n_14752)
);

OAI21xp5_ASAP7_75t_L g14753 ( 
.A1(n_14740),
.A2(n_14741),
.B(n_14744),
.Y(n_14753)
);

OA22x2_ASAP7_75t_L g14754 ( 
.A1(n_14743),
.A2(n_14707),
.B1(n_14713),
.B2(n_14709),
.Y(n_14754)
);

INVx1_ASAP7_75t_L g14755 ( 
.A(n_14725),
.Y(n_14755)
);

NAND4xp25_ASAP7_75t_L g14756 ( 
.A(n_14745),
.B(n_14735),
.C(n_14730),
.D(n_14720),
.Y(n_14756)
);

AOI22xp5_ASAP7_75t_L g14757 ( 
.A1(n_14746),
.A2(n_14739),
.B1(n_14736),
.B2(n_14731),
.Y(n_14757)
);

INVx2_ASAP7_75t_L g14758 ( 
.A(n_14751),
.Y(n_14758)
);

INVx1_ASAP7_75t_L g14759 ( 
.A(n_14747),
.Y(n_14759)
);

OAI221xp5_ASAP7_75t_L g14760 ( 
.A1(n_14753),
.A2(n_14700),
.B1(n_14706),
.B2(n_14742),
.C(n_14710),
.Y(n_14760)
);

NAND4xp25_ASAP7_75t_L g14761 ( 
.A(n_14755),
.B(n_14737),
.C(n_14696),
.D(n_5042),
.Y(n_14761)
);

INVx1_ASAP7_75t_L g14762 ( 
.A(n_14749),
.Y(n_14762)
);

INVx1_ASAP7_75t_L g14763 ( 
.A(n_14748),
.Y(n_14763)
);

NAND3xp33_ASAP7_75t_SL g14764 ( 
.A(n_14752),
.B(n_4637),
.C(n_4143),
.Y(n_14764)
);

XOR2xp5_ASAP7_75t_L g14765 ( 
.A(n_14754),
.B(n_14750),
.Y(n_14765)
);

NOR3x1_ASAP7_75t_L g14766 ( 
.A(n_14759),
.B(n_6939),
.C(n_6923),
.Y(n_14766)
);

INVx2_ASAP7_75t_L g14767 ( 
.A(n_14758),
.Y(n_14767)
);

OAI221xp5_ASAP7_75t_SL g14768 ( 
.A1(n_14765),
.A2(n_5044),
.B1(n_5069),
.B2(n_5042),
.C(n_5025),
.Y(n_14768)
);

OA22x2_ASAP7_75t_L g14769 ( 
.A1(n_14763),
.A2(n_14762),
.B1(n_14757),
.B2(n_14756),
.Y(n_14769)
);

AOI22x1_ASAP7_75t_L g14770 ( 
.A1(n_14760),
.A2(n_5639),
.B1(n_5691),
.B2(n_5667),
.Y(n_14770)
);

AND2x2_ASAP7_75t_SL g14771 ( 
.A(n_14761),
.B(n_4955),
.Y(n_14771)
);

OAI22xp5_ASAP7_75t_L g14772 ( 
.A1(n_14764),
.A2(n_4850),
.B1(n_6212),
.B2(n_5958),
.Y(n_14772)
);

HB1xp67_ASAP7_75t_L g14773 ( 
.A(n_14765),
.Y(n_14773)
);

OAI222xp33_ASAP7_75t_L g14774 ( 
.A1(n_14767),
.A2(n_4012),
.B1(n_4146),
.B2(n_4242),
.C1(n_4155),
.C2(n_4143),
.Y(n_14774)
);

INVx1_ASAP7_75t_L g14775 ( 
.A(n_14769),
.Y(n_14775)
);

INVx1_ASAP7_75t_L g14776 ( 
.A(n_14773),
.Y(n_14776)
);

OAI222xp33_ASAP7_75t_L g14777 ( 
.A1(n_14772),
.A2(n_4242),
.B1(n_4146),
.B2(n_4248),
.C1(n_4155),
.C2(n_4143),
.Y(n_14777)
);

OAI22xp5_ASAP7_75t_SL g14778 ( 
.A1(n_14775),
.A2(n_14771),
.B1(n_14770),
.B2(n_14768),
.Y(n_14778)
);

INVx1_ASAP7_75t_L g14779 ( 
.A(n_14776),
.Y(n_14779)
);

AOI22xp33_ASAP7_75t_L g14780 ( 
.A1(n_14779),
.A2(n_14777),
.B1(n_14774),
.B2(n_14766),
.Y(n_14780)
);

AOI21xp5_ASAP7_75t_L g14781 ( 
.A1(n_14778),
.A2(n_6212),
.B(n_5958),
.Y(n_14781)
);

NAND2xp5_ASAP7_75t_L g14782 ( 
.A(n_14780),
.B(n_4955),
.Y(n_14782)
);

NOR2xp33_ASAP7_75t_L g14783 ( 
.A(n_14781),
.B(n_4086),
.Y(n_14783)
);

OR2x6_ASAP7_75t_L g14784 ( 
.A(n_14782),
.B(n_5042),
.Y(n_14784)
);

INVx1_ASAP7_75t_L g14785 ( 
.A(n_14784),
.Y(n_14785)
);

OAI21xp33_ASAP7_75t_L g14786 ( 
.A1(n_14785),
.A2(n_14783),
.B(n_5561),
.Y(n_14786)
);

AOI221xp5_ASAP7_75t_L g14787 ( 
.A1(n_14786),
.A2(n_5691),
.B1(n_5740),
.B2(n_5667),
.C(n_5639),
.Y(n_14787)
);

AOI22xp5_ASAP7_75t_L g14788 ( 
.A1(n_14787),
.A2(n_5025),
.B1(n_5069),
.B2(n_5044),
.Y(n_14788)
);

AOI211xp5_ASAP7_75t_L g14789 ( 
.A1(n_14788),
.A2(n_5096),
.B(n_5112),
.C(n_5069),
.Y(n_14789)
);


endmodule