module fake_netlist_1_9974_n_14 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_14);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_9;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_3), .B(n_2), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_4), .B(n_6), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_10), .B(n_8), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
OAI22xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_9), .B1(n_1), .B2(n_2), .Y(n_13) );
OAI211xp5_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_0), .B(n_1), .C(n_12), .Y(n_14) );
endmodule