module fake_netlist_1_2238_n_695 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_695);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_695;
wire n_117;
wire n_663;
wire n_513;
wire n_361;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_476;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_285;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_L g79 ( .A(n_76), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_10), .Y(n_80) );
INVxp33_ASAP7_75t_SL g81 ( .A(n_4), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_46), .Y(n_82) );
OR2x2_ASAP7_75t_L g83 ( .A(n_24), .B(n_52), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_31), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_70), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_20), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_23), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_2), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_42), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_1), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_3), .Y(n_91) );
INVx1_ASAP7_75t_SL g92 ( .A(n_27), .Y(n_92) );
INVxp67_ASAP7_75t_L g93 ( .A(n_67), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_12), .Y(n_94) );
INVxp67_ASAP7_75t_L g95 ( .A(n_56), .Y(n_95) );
AND2x2_ASAP7_75t_L g96 ( .A(n_40), .B(n_75), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_10), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_6), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_44), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_65), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_71), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_72), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_32), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_69), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_68), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_55), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_48), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_36), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_59), .Y(n_109) );
INVxp67_ASAP7_75t_L g110 ( .A(n_17), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_63), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_29), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_61), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_0), .Y(n_114) );
INVxp33_ASAP7_75t_L g115 ( .A(n_19), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_16), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_57), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_53), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_35), .Y(n_119) );
INVxp33_ASAP7_75t_L g120 ( .A(n_77), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_39), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_22), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_37), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_13), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_15), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
INVx1_ASAP7_75t_SL g128 ( .A(n_107), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_115), .B(n_1), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_110), .B(n_2), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_80), .B(n_3), .Y(n_131) );
BUFx2_ASAP7_75t_L g132 ( .A(n_104), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
AOI22xp5_ASAP7_75t_L g134 ( .A1(n_81), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_87), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_99), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_97), .B(n_5), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_100), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_102), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_103), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_106), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_111), .B(n_117), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_121), .Y(n_143) );
BUFx2_ASAP7_75t_L g144 ( .A(n_122), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_88), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_88), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_123), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_91), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_83), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_98), .B(n_7), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_91), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_94), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_126), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_81), .B(n_7), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_83), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_116), .B(n_8), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_120), .B(n_8), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_114), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_114), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_124), .Y(n_162) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_124), .A2(n_38), .B(n_74), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_82), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_79), .B(n_9), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_85), .Y(n_166) );
OR2x6_ASAP7_75t_L g167 ( .A(n_96), .B(n_9), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_113), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_118), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_145), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_144), .B(n_122), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_144), .B(n_89), .Y(n_174) );
INVxp67_ASAP7_75t_L g175 ( .A(n_132), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_132), .B(n_105), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_167), .A2(n_105), .B1(n_119), .B2(n_101), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_145), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_164), .B(n_112), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_127), .B(n_101), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_157), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_127), .B(n_119), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_160), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_133), .B(n_108), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_149), .B(n_96), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_160), .A2(n_125), .B1(n_95), .B2(n_93), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_164), .B(n_92), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_160), .A2(n_109), .B1(n_107), .B2(n_90), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_163), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_133), .B(n_109), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_166), .B(n_90), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_149), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_160), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_166), .B(n_34), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_163), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_135), .B(n_11), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_161), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_135), .B(n_11), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_167), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_167), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_136), .B(n_17), .Y(n_202) );
INVx2_ASAP7_75t_SL g203 ( .A(n_157), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_161), .A2(n_18), .B1(n_19), .B2(n_78), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_136), .B(n_18), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_149), .B(n_21), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_138), .B(n_25), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_157), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_149), .B(n_26), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_146), .B(n_73), .Y(n_210) );
BUFx5_ASAP7_75t_L g211 ( .A(n_148), .Y(n_211) );
INVx1_ASAP7_75t_SL g212 ( .A(n_128), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_149), .B(n_28), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_138), .B(n_30), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_157), .B(n_33), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_161), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_161), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_139), .B(n_41), .Y(n_218) );
OR2x2_ASAP7_75t_L g219 ( .A(n_168), .B(n_43), .Y(n_219) );
NOR3xp33_ASAP7_75t_L g220 ( .A(n_156), .B(n_45), .C(n_47), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_154), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_139), .B(n_49), .Y(n_222) );
NAND3xp33_ASAP7_75t_L g223 ( .A(n_157), .B(n_50), .C(n_51), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_140), .B(n_54), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_140), .B(n_58), .Y(n_225) );
NOR2xp33_ASAP7_75t_SL g226 ( .A(n_167), .B(n_60), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_143), .B(n_62), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_148), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_163), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_191), .B(n_167), .Y(n_230) );
INVx1_ASAP7_75t_SL g231 ( .A(n_212), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_221), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_178), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_181), .B(n_169), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_178), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_221), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_182), .Y(n_237) );
AND2x6_ASAP7_75t_L g238 ( .A(n_200), .B(n_165), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_175), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_183), .B(n_169), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_174), .B(n_168), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_174), .B(n_165), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_177), .B(n_165), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_203), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_193), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_190), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_190), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_190), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_171), .B(n_142), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_208), .Y(n_250) );
INVx4_ASAP7_75t_L g251 ( .A(n_211), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_195), .A2(n_152), .B(n_151), .C(n_153), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_193), .Y(n_253) );
OR2x6_ASAP7_75t_L g254 ( .A(n_186), .B(n_165), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_170), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_192), .Y(n_256) );
INVx4_ASAP7_75t_L g257 ( .A(n_211), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_188), .B(n_143), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_188), .B(n_129), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_172), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_228), .A2(n_159), .B(n_153), .C(n_151), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_179), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_179), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_173), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_192), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_211), .B(n_147), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_211), .B(n_147), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_198), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_180), .B(n_152), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_186), .A2(n_163), .B(n_141), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_184), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_210), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_201), .A2(n_134), .B1(n_158), .B2(n_131), .Y(n_273) );
NOR2xp33_ASAP7_75t_SL g274 ( .A(n_226), .B(n_130), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_184), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_219), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_180), .B(n_141), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_216), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_185), .B(n_154), .Y(n_279) );
CKINVDCx16_ASAP7_75t_R g280 ( .A(n_176), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_211), .B(n_155), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_211), .B(n_155), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_197), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_190), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_196), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_187), .B(n_162), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_187), .B(n_137), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_194), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_194), .B(n_217), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_206), .A2(n_150), .B(n_162), .Y(n_290) );
INVx4_ASAP7_75t_L g291 ( .A(n_217), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_195), .B(n_64), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_196), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_231), .Y(n_294) );
CKINVDCx16_ASAP7_75t_R g295 ( .A(n_239), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_270), .A2(n_229), .B(n_196), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_235), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_256), .B(n_189), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_251), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_266), .A2(n_229), .B(n_196), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_243), .B(n_220), .Y(n_301) );
OR2x6_ASAP7_75t_L g302 ( .A(n_243), .B(n_189), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_267), .A2(n_229), .B(n_209), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_243), .B(n_205), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_280), .B(n_199), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_238), .A2(n_202), .B1(n_204), .B2(n_224), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_238), .A2(n_204), .B1(n_225), .B2(n_207), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_276), .B(n_206), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_259), .B(n_218), .Y(n_309) );
BUFx2_ASAP7_75t_SL g310 ( .A(n_251), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_252), .A2(n_214), .B(n_227), .C(n_222), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_279), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_279), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_255), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_246), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_251), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_246), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_259), .B(n_209), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_283), .B(n_229), .Y(n_319) );
NOR2x1_ASAP7_75t_SL g320 ( .A(n_254), .B(n_215), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_238), .A2(n_213), .B1(n_223), .B2(n_66), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_265), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_238), .A2(n_287), .B1(n_277), .B2(n_269), .Y(n_323) );
NAND2x1p5_ASAP7_75t_L g324 ( .A(n_257), .B(n_291), .Y(n_324) );
AOI21xp33_ASAP7_75t_L g325 ( .A1(n_230), .A2(n_272), .B(n_241), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_257), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_290), .A2(n_242), .B(n_282), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_269), .B(n_230), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_235), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_281), .A2(n_289), .B(n_252), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_265), .B(n_287), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_260), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_287), .B(n_258), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_254), .A2(n_240), .B1(n_234), .B2(n_286), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_291), .Y(n_335) );
OR2x6_ASAP7_75t_L g336 ( .A(n_254), .B(n_257), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_277), .B(n_249), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_264), .A2(n_268), .B(n_278), .Y(n_338) );
INVx5_ASAP7_75t_L g339 ( .A(n_291), .Y(n_339) );
AOI21xp33_ASAP7_75t_SL g340 ( .A1(n_273), .A2(n_249), .B(n_277), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_238), .A2(n_254), .B1(n_232), .B2(n_236), .Y(n_341) );
CKINVDCx11_ASAP7_75t_R g342 ( .A(n_263), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_233), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_233), .B(n_245), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_314), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_312), .B(n_275), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_328), .A2(n_275), .B1(n_263), .B2(n_262), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_294), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_315), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_315), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_342), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_315), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_328), .B(n_288), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_317), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_332), .Y(n_356) );
OAI31xp33_ASAP7_75t_L g357 ( .A1(n_298), .A2(n_261), .A3(n_274), .B(n_292), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_317), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_296), .A2(n_233), .B(n_288), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_295), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_317), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_316), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_316), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_302), .A2(n_271), .B1(n_288), .B2(n_262), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_339), .Y(n_365) );
A2O1A1Ixp33_ASAP7_75t_L g366 ( .A1(n_340), .A2(n_271), .B(n_262), .C(n_245), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_317), .Y(n_367) );
AO21x2_ASAP7_75t_L g368 ( .A1(n_296), .A2(n_237), .B(n_244), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_323), .B(n_313), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_324), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_324), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_299), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_338), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_299), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_338), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_310), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_333), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_371), .Y(n_378) );
NAND2x1_ASAP7_75t_L g379 ( .A(n_370), .B(n_326), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_359), .Y(n_380) );
NOR2x1_ASAP7_75t_SL g381 ( .A(n_370), .B(n_336), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_377), .B(n_323), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_377), .B(n_302), .Y(n_383) );
OA21x2_ASAP7_75t_L g384 ( .A1(n_359), .A2(n_303), .B(n_300), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_359), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_349), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_369), .B(n_346), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_369), .A2(n_302), .B1(n_301), .B2(n_322), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_369), .B(n_331), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_345), .Y(n_390) );
AOI33xp33_ASAP7_75t_L g391 ( .A1(n_345), .A2(n_305), .A3(n_337), .B1(n_341), .B2(n_301), .B3(n_318), .Y(n_391) );
INVxp67_ASAP7_75t_L g392 ( .A(n_346), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_356), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_349), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_356), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_365), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_373), .Y(n_397) );
OAI211xp5_ASAP7_75t_L g398 ( .A1(n_364), .A2(n_341), .B(n_325), .C(n_304), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_346), .B(n_336), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_371), .B(n_336), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_373), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_365), .Y(n_402) );
NAND3xp33_ASAP7_75t_L g403 ( .A(n_357), .B(n_307), .C(n_306), .Y(n_403) );
NAND2x1_ASAP7_75t_L g404 ( .A(n_370), .B(n_326), .Y(n_404) );
NOR4xp25_ASAP7_75t_SL g405 ( .A(n_351), .B(n_311), .C(n_343), .D(n_308), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_397), .Y(n_406) );
AO21x2_ASAP7_75t_L g407 ( .A1(n_403), .A2(n_366), .B(n_375), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_387), .B(n_348), .Y(n_408) );
AND4x1_ASAP7_75t_L g409 ( .A(n_391), .B(n_364), .C(n_376), .D(n_357), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_378), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_397), .Y(n_411) );
OAI21x1_ASAP7_75t_L g412 ( .A1(n_380), .A2(n_375), .B(n_300), .Y(n_412) );
INVx5_ASAP7_75t_L g413 ( .A(n_378), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_401), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_401), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_387), .B(n_348), .Y(n_416) );
O2A1O1Ixp5_ASAP7_75t_L g417 ( .A1(n_398), .A2(n_403), .B(n_385), .C(n_380), .Y(n_417) );
INVx2_ASAP7_75t_SL g418 ( .A(n_378), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_390), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_382), .B(n_363), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_387), .B(n_368), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
OAI211xp5_ASAP7_75t_L g423 ( .A1(n_388), .A2(n_348), .B(n_376), .C(n_304), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_380), .Y(n_424) );
AOI21xp33_ASAP7_75t_L g425 ( .A1(n_398), .A2(n_334), .B(n_308), .Y(n_425) );
NAND3xp33_ASAP7_75t_SL g426 ( .A(n_405), .B(n_360), .C(n_347), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_390), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_396), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_386), .B(n_368), .Y(n_429) );
INVxp67_ASAP7_75t_L g430 ( .A(n_402), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_385), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_393), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_393), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_392), .A2(n_347), .B1(n_309), .B2(n_366), .C(n_308), .Y(n_434) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_385), .B(n_362), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_386), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_402), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_379), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_382), .B(n_362), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_421), .B(n_406), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_424), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_424), .Y(n_443) );
NAND2x1_ASAP7_75t_L g444 ( .A(n_438), .B(n_395), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_419), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_408), .B(n_389), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_408), .B(n_389), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_421), .B(n_383), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_416), .B(n_382), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_413), .B(n_395), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_416), .B(n_383), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_421), .B(n_383), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_419), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_406), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_406), .Y(n_455) );
OAI21xp33_ASAP7_75t_L g456 ( .A1(n_423), .A2(n_321), .B(n_399), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_424), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_413), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_427), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_415), .B(n_399), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_427), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_415), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_431), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_437), .B(n_392), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_431), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_431), .Y(n_466) );
NOR2xp33_ASAP7_75t_SL g467 ( .A(n_413), .B(n_400), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_423), .A2(n_330), .B(n_327), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_437), .B(n_399), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_436), .Y(n_470) );
OR2x6_ASAP7_75t_L g471 ( .A(n_410), .B(n_404), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_436), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_432), .B(n_400), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_432), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_433), .B(n_363), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_433), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_422), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_430), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_420), .B(n_337), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_420), .B(n_381), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_440), .B(n_381), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_440), .B(n_405), .Y(n_482) );
INVx3_ASAP7_75t_L g483 ( .A(n_413), .Y(n_483) );
INVxp67_ASAP7_75t_L g484 ( .A(n_422), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_428), .B(n_394), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_415), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_428), .B(n_394), .Y(n_487) );
INVxp33_ASAP7_75t_L g488 ( .A(n_410), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_411), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_441), .B(n_429), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_442), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_441), .B(n_429), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_445), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_453), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_456), .A2(n_426), .B1(n_434), .B2(n_439), .Y(n_495) );
OAI222xp33_ASAP7_75t_L g496 ( .A1(n_446), .A2(n_434), .B1(n_430), .B2(n_413), .C1(n_418), .C2(n_439), .Y(n_496) );
INVx2_ASAP7_75t_SL g497 ( .A(n_483), .Y(n_497) );
INVxp33_ASAP7_75t_L g498 ( .A(n_467), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_448), .B(n_429), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_448), .B(n_414), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_452), .B(n_411), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_459), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_446), .B(n_426), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_442), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_443), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_452), .B(n_414), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_454), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_460), .B(n_429), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_483), .Y(n_509) );
INVx2_ASAP7_75t_SL g510 ( .A(n_483), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_461), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_474), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_460), .B(n_429), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_443), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_476), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_489), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_454), .B(n_435), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_455), .B(n_435), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_455), .B(n_435), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_447), .B(n_439), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_447), .B(n_418), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_478), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_469), .B(n_407), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_462), .B(n_407), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_458), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_462), .B(n_407), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_473), .B(n_418), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_449), .B(n_436), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_469), .B(n_407), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_457), .Y(n_530) );
INVxp67_ASAP7_75t_SL g531 ( .A(n_485), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_457), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_486), .B(n_438), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_458), .B(n_413), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_485), .B(n_412), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_450), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_487), .B(n_412), .Y(n_537) );
INVxp67_ASAP7_75t_SL g538 ( .A(n_487), .Y(n_538) );
OAI221xp5_ASAP7_75t_L g539 ( .A1(n_482), .A2(n_409), .B1(n_425), .B2(n_417), .C(n_321), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_486), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_464), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_464), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_470), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_463), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_475), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_488), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_480), .A2(n_425), .B1(n_413), .B2(n_354), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_525), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_542), .B(n_477), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_522), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_541), .B(n_484), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_531), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_493), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_509), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_494), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_545), .B(n_451), .Y(n_556) );
NOR2x1_ASAP7_75t_L g557 ( .A(n_534), .B(n_471), .Y(n_557) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_495), .A2(n_481), .B1(n_471), .B2(n_488), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_502), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_546), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_511), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_500), .B(n_472), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_512), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_515), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_498), .A2(n_471), .B1(n_444), .B2(n_479), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_499), .B(n_471), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_501), .B(n_472), .Y(n_567) );
OAI31xp33_ASAP7_75t_L g568 ( .A1(n_503), .A2(n_438), .A3(n_470), .B(n_409), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_516), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_500), .B(n_506), .Y(n_570) );
INVx3_ASAP7_75t_L g571 ( .A(n_533), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_507), .Y(n_572) );
NAND2xp33_ASAP7_75t_SL g573 ( .A(n_498), .B(n_444), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_499), .B(n_466), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_538), .B(n_466), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_536), .B(n_468), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_535), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_496), .B(n_438), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_521), .B(n_463), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_520), .B(n_465), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_507), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_534), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_539), .B(n_465), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_492), .B(n_412), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_540), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_492), .B(n_417), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_497), .B(n_394), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_527), .B(n_404), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_535), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_517), .Y(n_590) );
AOI21xp33_ASAP7_75t_SL g591 ( .A1(n_497), .A2(n_384), .B(n_374), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_517), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_518), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_510), .B(n_379), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_518), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_519), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_519), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_528), .B(n_384), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_537), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_537), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g601 ( .A(n_558), .B(n_510), .C(n_526), .Y(n_601) );
NAND3xp33_ASAP7_75t_SL g602 ( .A(n_568), .B(n_547), .C(n_523), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_583), .A2(n_490), .B1(n_533), .B2(n_513), .Y(n_603) );
AND4x1_ASAP7_75t_L g604 ( .A(n_557), .B(n_513), .C(n_508), .D(n_526), .Y(n_604) );
AOI221xp5_ASAP7_75t_L g605 ( .A1(n_576), .A2(n_490), .B1(n_524), .B2(n_523), .C(n_529), .Y(n_605) );
INVxp67_ASAP7_75t_L g606 ( .A(n_552), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_599), .B(n_524), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_566), .B(n_490), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_583), .A2(n_533), .B1(n_508), .B2(n_529), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_576), .B(n_543), .C(n_544), .Y(n_610) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_578), .B(n_588), .C(n_565), .D(n_560), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_548), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_550), .B(n_543), .Y(n_613) );
AND4x1_ASAP7_75t_L g614 ( .A(n_578), .B(n_330), .C(n_327), .D(n_354), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_589), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_574), .B(n_544), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_570), .B(n_532), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_553), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_577), .B(n_532), .Y(n_619) );
NAND4xp25_ASAP7_75t_SL g620 ( .A(n_554), .B(n_491), .C(n_514), .D(n_505), .Y(n_620) );
NAND5xp2_ASAP7_75t_L g621 ( .A(n_588), .B(n_303), .C(n_354), .D(n_319), .E(n_320), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_558), .A2(n_530), .B1(n_514), .B2(n_505), .Y(n_622) );
NOR3x1_ASAP7_75t_L g623 ( .A(n_549), .B(n_530), .C(n_504), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_573), .B(n_504), .Y(n_624) );
NAND4xp25_ASAP7_75t_L g625 ( .A(n_551), .B(n_491), .C(n_329), .D(n_297), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_582), .A2(n_372), .B(n_374), .C(n_386), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_570), .B(n_372), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_591), .B(n_384), .C(n_374), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_555), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_600), .B(n_593), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_556), .B(n_372), .Y(n_631) );
AOI211x1_ASAP7_75t_SL g632 ( .A1(n_587), .A2(n_358), .B(n_355), .C(n_353), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_579), .A2(n_372), .B1(n_368), .B2(n_335), .C(n_344), .Y(n_633) );
NAND2xp33_ASAP7_75t_L g634 ( .A(n_573), .B(n_358), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_559), .Y(n_635) );
AOI211x1_ASAP7_75t_L g636 ( .A1(n_561), .A2(n_250), .B(n_384), .C(n_253), .Y(n_636) );
OAI221xp5_ASAP7_75t_SL g637 ( .A1(n_586), .A2(n_372), .B1(n_349), .B2(n_367), .C(n_361), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_563), .Y(n_638) );
INVx6_ASAP7_75t_L g639 ( .A(n_619), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_611), .B(n_594), .C(n_587), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_605), .A2(n_564), .B1(n_569), .B2(n_579), .C(n_596), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g642 ( .A(n_602), .B(n_594), .C(n_571), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_601), .A2(n_584), .B1(n_590), .B2(n_597), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_605), .A2(n_592), .B1(n_595), .B2(n_600), .C(n_585), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_621), .A2(n_571), .B1(n_580), .B2(n_598), .Y(n_645) );
NOR2xp33_ASAP7_75t_SL g646 ( .A(n_612), .B(n_562), .Y(n_646) );
INVxp67_ASAP7_75t_L g647 ( .A(n_615), .Y(n_647) );
OAI32xp33_ASAP7_75t_L g648 ( .A1(n_606), .A2(n_575), .A3(n_567), .B1(n_572), .B2(n_581), .Y(n_648) );
NOR2x1_ASAP7_75t_SL g649 ( .A(n_624), .B(n_368), .Y(n_649) );
NOR2xp67_ASAP7_75t_L g650 ( .A(n_620), .B(n_358), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_609), .B(n_384), .Y(n_651) );
AOI32xp33_ASAP7_75t_L g652 ( .A1(n_634), .A2(n_367), .A3(n_361), .B1(n_355), .B2(n_353), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_614), .B(n_367), .C(n_361), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_618), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g655 ( .A1(n_633), .A2(n_344), .B1(n_353), .B2(n_352), .C1(n_350), .C2(n_355), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_623), .B(n_352), .Y(n_656) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_628), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_617), .B(n_352), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_629), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g660 ( .A1(n_603), .A2(n_339), .B1(n_350), .B2(n_247), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_637), .A2(n_339), .B1(n_350), .B2(n_247), .Y(n_661) );
NAND4xp25_ASAP7_75t_SL g662 ( .A(n_641), .B(n_633), .C(n_622), .D(n_604), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_642), .A2(n_627), .B1(n_613), .B2(n_631), .Y(n_663) );
OAI222xp33_ASAP7_75t_R g664 ( .A1(n_643), .A2(n_638), .B1(n_635), .B2(n_610), .C1(n_625), .C2(n_636), .Y(n_664) );
NOR2x1_ASAP7_75t_L g665 ( .A(n_653), .B(n_626), .Y(n_665) );
NOR3xp33_ASAP7_75t_L g666 ( .A(n_640), .B(n_626), .C(n_630), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_644), .B(n_607), .Y(n_667) );
AOI211xp5_ASAP7_75t_L g668 ( .A1(n_648), .A2(n_608), .B(n_616), .C(n_632), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_647), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_657), .B(n_339), .C(n_246), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_639), .B(n_293), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_654), .A2(n_271), .B1(n_246), .B2(n_247), .C(n_248), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_645), .B(n_247), .Y(n_673) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_657), .B(n_248), .C(n_284), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_659), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_675), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_669), .A2(n_639), .B1(n_650), .B2(n_656), .Y(n_677) );
AO21x2_ASAP7_75t_L g678 ( .A1(n_666), .A2(n_649), .B(n_651), .Y(n_678) );
XNOR2xp5_ASAP7_75t_L g679 ( .A(n_663), .B(n_660), .Y(n_679) );
XNOR2xp5_ASAP7_75t_L g680 ( .A(n_668), .B(n_658), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_662), .A2(n_646), .B1(n_657), .B2(n_655), .Y(n_681) );
INVx4_ASAP7_75t_L g682 ( .A(n_671), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g683 ( .A1(n_667), .A2(n_661), .B1(n_652), .B2(n_284), .Y(n_683) );
OR4x1_ASAP7_75t_L g684 ( .A(n_681), .B(n_664), .C(n_665), .D(n_666), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_676), .Y(n_685) );
AOI311xp33_ASAP7_75t_L g686 ( .A1(n_677), .A2(n_673), .A3(n_672), .B(n_670), .C(n_674), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_679), .B(n_293), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_680), .A2(n_248), .B1(n_284), .B2(n_285), .Y(n_688) );
OAI222xp33_ASAP7_75t_L g689 ( .A1(n_685), .A2(n_682), .B1(n_683), .B2(n_678), .C1(n_245), .C2(n_285), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_687), .B(n_682), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_688), .B(n_248), .Y(n_691) );
XNOR2xp5_ASAP7_75t_L g692 ( .A(n_690), .B(n_688), .Y(n_692) );
INVx4_ASAP7_75t_L g693 ( .A(n_691), .Y(n_693) );
OAI222xp33_ASAP7_75t_L g694 ( .A1(n_692), .A2(n_684), .B1(n_689), .B2(n_686), .C1(n_284), .C2(n_293), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_694), .A2(n_285), .B1(n_293), .B2(n_693), .C(n_684), .Y(n_695) );
endmodule