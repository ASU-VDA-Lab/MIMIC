module real_jpeg_33640_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_0),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_0),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_1),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_1),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_1),
.A2(n_142),
.B1(n_189),
.B2(n_192),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_1),
.A2(n_142),
.B1(n_286),
.B2(n_288),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_2),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_3),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_3),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_4),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_5),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_5),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_5),
.A2(n_133),
.B1(n_217),
.B2(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_5),
.A2(n_133),
.B1(n_320),
.B2(n_324),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_5),
.A2(n_133),
.B1(n_368),
.B2(n_373),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_6),
.A2(n_145),
.B1(n_146),
.B2(n_152),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_6),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_6),
.A2(n_145),
.B1(n_203),
.B2(n_206),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_6),
.A2(n_145),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_6),
.A2(n_145),
.B1(n_377),
.B2(n_378),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_7),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_8),
.A2(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_8),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_8),
.A2(n_139),
.B1(n_174),
.B2(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_8),
.A2(n_174),
.B1(n_343),
.B2(n_348),
.Y(n_342)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_9),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_10),
.A2(n_48),
.B1(n_51),
.B2(n_56),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_10),
.A2(n_56),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_11),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_11),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_12),
.Y(n_102)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_13),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_14),
.A2(n_118),
.B(n_123),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_14),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_14),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_14),
.B(n_181),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_14),
.A2(n_75),
.B1(n_367),
.B2(n_385),
.Y(n_384)
);

OAI32xp33_ASAP7_75t_L g408 ( 
.A1(n_14),
.A2(n_156),
.A3(n_293),
.B1(n_409),
.B2(n_410),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_14),
.A2(n_152),
.B1(n_261),
.B2(n_414),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_15),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_15),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_15),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_16),
.A2(n_35),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_264),
.Y(n_17)
);

NAND2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_262),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_238),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_20),
.B(n_238),
.Y(n_263)
);

XNOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_183),
.Y(n_20)
);

XNOR2x1_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_91),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_67),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_34),
.B1(n_47),
.B2(n_57),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_24),
.A2(n_47),
.B1(n_57),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_24),
.A2(n_57),
.B1(n_138),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_24),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_24),
.A2(n_57),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_24),
.B(n_261),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_25),
.Y(n_417)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AO21x2_ASAP7_75t_L g57 ( 
.A1(n_26),
.A2(n_58),
.B(n_63),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_26)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_27),
.Y(n_391)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_28),
.Y(n_255)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_29),
.Y(n_235)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B(n_41),
.Y(n_34)
);

BUFx2_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_38),
.Y(n_317)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_42),
.Y(n_141)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_46),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_46),
.Y(n_280)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_46),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_50),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_54),
.Y(n_360)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_55),
.Y(n_314)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_57),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_62),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_63),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_75),
.B1(n_81),
.B2(n_88),
.Y(n_67)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_68),
.Y(n_227)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_69),
.Y(n_330)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_70),
.Y(n_236)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_70),
.Y(n_372)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_75),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_75),
.A2(n_342),
.B1(n_350),
.B2(n_352),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_75),
.A2(n_367),
.B1(n_376),
.B2(n_381),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_78),
.Y(n_289)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_80),
.Y(n_258)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_80),
.Y(n_287)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_80),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_80),
.Y(n_349)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_80),
.Y(n_375)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_89),
.Y(n_259)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g291 ( 
.A(n_90),
.Y(n_291)
);

INVx8_ASAP7_75t_L g381 ( 
.A(n_90),
.Y(n_381)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_136),
.C(n_143),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_93),
.B(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_117),
.B1(n_128),
.B2(n_129),
.Y(n_93)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_94),
.Y(n_199)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_108),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_101),
.B1(n_103),
.B2(n_105),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_100),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_100),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_102),
.Y(n_216)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

AOI22x1_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_114),
.B2(n_116),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_112),
.Y(n_219)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_112),
.Y(n_300)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_118),
.Y(n_222)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AO21x1_ASAP7_75t_L g211 ( 
.A1(n_123),
.A2(n_212),
.B(n_220),
.Y(n_211)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_128),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_128),
.B(n_261),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g198 ( 
.A(n_129),
.Y(n_198)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_136),
.A2(n_137),
.B1(n_143),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_155),
.B1(n_173),
.B2(n_180),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_144),
.A2(n_155),
.B1(n_180),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_151),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_173),
.B1(n_188),
.B2(n_194),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_155),
.A2(n_194),
.B1(n_246),
.B2(n_413),
.Y(n_412)
);

AO21x2_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_161),
.B(n_166),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_156),
.A2(n_293),
.B(n_299),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_171),
.Y(n_166)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

XNOR2x1_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_210),
.Y(n_183)
);

OAI21x1_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_195),
.B(n_209),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_197),
.Y(n_209)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_191),
.Y(n_414)
);

INVx3_ASAP7_75t_SL g224 ( 
.A(n_192),
.Y(n_224)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22x1_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_225),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_211),
.A2(n_225),
.B1(n_226),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_221),
.C(n_223),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_233),
.B2(n_237),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_229),
.B(n_261),
.Y(n_388)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_231),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_232),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_237),
.B1(n_253),
.B2(n_259),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_237),
.A2(n_253),
.B1(n_285),
.B2(n_290),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_237),
.A2(n_395),
.B1(n_396),
.B2(n_397),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.C(n_244),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_244),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_251),
.C(n_260),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_252),
.B1(n_260),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_294),
.Y(n_293)
);

NAND3xp33_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_300),
.C(n_301),
.Y(n_299)
);

OAI21xp33_ASAP7_75t_SL g311 ( 
.A1(n_261),
.A2(n_312),
.B(n_315),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_261),
.B(n_316),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_304),
.B(n_427),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_268),
.B(n_270),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_275),
.C(n_281),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_271),
.A2(n_272),
.B1(n_421),
.B2(n_422),
.Y(n_420)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_275),
.A2(n_281),
.B1(n_282),
.B2(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_275),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_277),
.A2(n_318),
.B1(n_416),
.B2(n_417),
.Y(n_415)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_280),
.Y(n_358)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_292),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_283),
.A2(n_284),
.B1(n_292),
.B2(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_285),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_287),
.Y(n_338)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_300),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_301),
.Y(n_410)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_419),
.B(n_426),
.Y(n_304)
);

AOI21x1_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_403),
.B(n_418),
.Y(n_305)
);

OAI21x1_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_363),
.B(n_402),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_340),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_308),
.B(n_340),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_327),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_309),
.A2(n_310),
.B1(n_327),
.B2(n_328),
.Y(n_400)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_318),
.B1(n_319),
.B2(n_326),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_315),
.Y(n_335)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_319),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_335),
.B1(n_336),
.B2(n_339),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_353),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_341),
.B(n_355),
.C(n_361),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_342),
.Y(n_396)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_346),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_349),
.Y(n_380)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_355),
.B1(n_361),
.B2(n_362),
.Y(n_353)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_354),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_355),
.Y(n_362)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_357),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_364),
.A2(n_393),
.B(n_401),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_383),
.B(n_392),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_382),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_366),
.B(n_382),
.Y(n_392)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_376),
.Y(n_395)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_400),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_394),
.B(n_400),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

NOR2x1_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_405),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_411),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_415),
.C(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.Y(n_411)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_412),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_424),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_420),
.B(n_424),
.Y(n_426)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);


endmodule