module fake_jpeg_25646_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_8),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_21),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_62),
.Y(n_80)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_58),
.B(n_67),
.Y(n_99)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx5_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_38),
.Y(n_76)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_33),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_25),
.B1(n_35),
.B2(n_26),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_49),
.B1(n_48),
.B2(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_21),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_75),
.A2(n_79),
.B1(n_94),
.B2(n_101),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_76),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_81),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_49),
.B1(n_45),
.B2(n_26),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_83),
.B(n_86),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_17),
.B1(n_31),
.B2(n_24),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_96),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_23),
.B(n_28),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_87),
.B(n_88),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_28),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_90),
.Y(n_147)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_93),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_26),
.B1(n_35),
.B2(n_42),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_70),
.B(n_34),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_95),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_63),
.B(n_37),
.CI(n_41),
.CON(n_96),
.SN(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g146 ( 
.A(n_97),
.Y(n_146)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_45),
.B1(n_35),
.B2(n_38),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_104),
.B1(n_22),
.B2(n_46),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_66),
.A2(n_33),
.B1(n_24),
.B2(n_34),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_65),
.A2(n_40),
.B1(n_47),
.B2(n_29),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_6),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_80),
.Y(n_116)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_30),
.Y(n_107)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_0),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_40),
.B1(n_29),
.B2(n_3),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g110 ( 
.A(n_68),
.Y(n_110)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_59),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_116),
.B(n_30),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_84),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_126),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_37),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_30),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_75),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_136),
.A2(n_82),
.B1(n_109),
.B2(n_98),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_92),
.A2(n_113),
.B1(n_90),
.B2(n_97),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_85),
.B1(n_103),
.B2(n_73),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_91),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_148),
.B(n_151),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_100),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_150),
.A2(n_160),
.B(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_91),
.Y(n_151)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_153),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_100),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_157),
.B1(n_110),
.B2(n_146),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_94),
.B1(n_112),
.B2(n_82),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_146),
.B1(n_142),
.B2(n_123),
.Y(n_183)
);

AO22x2_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_43),
.B1(n_44),
.B2(n_89),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_159),
.A2(n_142),
.B1(n_138),
.B2(n_132),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_162),
.Y(n_184)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_166),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_116),
.B(n_143),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_44),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_167),
.A2(n_170),
.B(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_128),
.B(n_27),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_122),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_85),
.B1(n_121),
.B2(n_118),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_89),
.Y(n_172)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

AND2x6_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_14),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_145),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_181),
.B(n_190),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_183),
.A2(n_211),
.B1(n_197),
.B2(n_178),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_147),
.B(n_123),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_185),
.A2(n_205),
.B(n_175),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_168),
.B(n_150),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_194),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_188),
.A2(n_193),
.B1(n_209),
.B2(n_167),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_138),
.C(n_44),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_137),
.Y(n_194)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_207),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_41),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_169),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_150),
.A2(n_132),
.B(n_144),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_201),
.A2(n_203),
.B(n_175),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_202),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_155),
.A2(n_149),
.B(n_160),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_156),
.B(n_8),
.Y(n_205)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_159),
.A2(n_118),
.B1(n_121),
.B2(n_141),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_141),
.B1(n_144),
.B2(n_46),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_185),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

XOR2x1_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_216),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_161),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_220),
.B(n_224),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_179),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_222),
.Y(n_242)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_223),
.A2(n_241),
.B1(n_211),
.B2(n_210),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_172),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_208),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_226),
.Y(n_243)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_164),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_227),
.B(n_228),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_153),
.B(n_159),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_191),
.B(n_176),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_232),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_199),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_159),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_236),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_184),
.B(n_177),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_237),
.A2(n_238),
.B1(n_206),
.B2(n_200),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_203),
.A2(n_173),
.B1(n_174),
.B2(n_18),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_184),
.B(n_162),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_240),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_187),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_204),
.A2(n_163),
.B1(n_32),
.B2(n_19),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_19),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_223),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_194),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_181),
.C(n_187),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_234),
.C(n_230),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_265),
.B1(n_237),
.B2(n_231),
.Y(n_272)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_219),
.A2(n_180),
.B(n_182),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_259),
.Y(n_279)
);

A2O1A1O1Ixp25_ASAP7_75t_L g259 ( 
.A1(n_230),
.A2(n_180),
.B(n_205),
.C(n_191),
.D(n_182),
.Y(n_259)
);

NOR4xp25_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_196),
.C(n_41),
.D(n_27),
.Y(n_261)
);

NAND3xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_22),
.C(n_11),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_213),
.B(n_196),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_240),
.C(n_226),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_27),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_241),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_264),
.A2(n_260),
.B1(n_259),
.B2(n_258),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_222),
.A2(n_46),
.B1(n_32),
.B2(n_19),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_235),
.B(n_229),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_266),
.B(n_271),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_280),
.C(n_256),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_275),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_276),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_250),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_274),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_264),
.B(n_214),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_277),
.B(n_278),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_247),
.B(n_214),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_217),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_218),
.C(n_32),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_242),
.C(n_253),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_283),
.A2(n_249),
.B1(n_265),
.B2(n_248),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_255),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_275),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_291),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_288),
.A2(n_295),
.B1(n_282),
.B2(n_270),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_245),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_293),
.A2(n_9),
.B(n_2),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_243),
.B1(n_257),
.B2(n_242),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_257),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_298),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_243),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_218),
.C(n_6),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_283),
.C(n_271),
.Y(n_309)
);

NOR2xp67_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_279),
.Y(n_304)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_305),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_306),
.B(n_297),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_273),
.Y(n_307)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_267),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_309),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_281),
.B(n_8),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_313),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_14),
.C(n_12),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_299),
.C(n_290),
.Y(n_317)
);

OAI31xp33_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_298),
.A3(n_300),
.B(n_299),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_312),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_303),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_319),
.C(n_311),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_290),
.C(n_301),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_314),
.B(n_319),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_323),
.B(n_325),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_328),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_310),
.B(n_302),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_317),
.B(n_302),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_327),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_318),
.C(n_309),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_320),
.B(n_312),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_329),
.B(n_320),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_9),
.C(n_3),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_335),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_9),
.C(n_4),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_331),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_330),
.B(n_4),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_5),
.B(n_0),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_340),
.B(n_0),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_4),
.Y(n_342)
);


endmodule