module fake_jpeg_7962_n_261 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_261);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_0),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_18),
.Y(n_47)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NAND2x1_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

NAND2x1_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_20),
.Y(n_53)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_44),
.B1(n_25),
.B2(n_13),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_19),
.B(n_16),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_53),
.B(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_14),
.B1(n_23),
.B2(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_59),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_57),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx2_ASAP7_75t_SL g91 ( 
.A(n_60),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_71),
.B1(n_53),
.B2(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_73),
.Y(n_77)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_75),
.B(n_80),
.Y(n_100)
);

XNOR2x1_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_90),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_82),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_88),
.B1(n_38),
.B2(n_49),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_53),
.B1(n_35),
.B2(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_89),
.B1(n_92),
.B2(n_33),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_70),
.B1(n_35),
.B2(n_62),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_51),
.B1(n_54),
.B2(n_39),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_27),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_70),
.B1(n_43),
.B2(n_38),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_106),
.B1(n_108),
.B2(n_111),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_28),
.B(n_13),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_107),
.B(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_107),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_68),
.B1(n_39),
.B2(n_48),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_28),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_48),
.B1(n_61),
.B2(n_64),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_79),
.B1(n_78),
.B2(n_33),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_72),
.B1(n_67),
.B2(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_32),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_85),
.Y(n_130)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_120),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_122),
.B(n_123),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_77),
.B1(n_75),
.B2(n_74),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_125),
.B1(n_102),
.B2(n_101),
.Y(n_137)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_127),
.B(n_128),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_77),
.B1(n_93),
.B2(n_37),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_27),
.Y(n_135)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_95),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_132),
.B1(n_134),
.B2(n_85),
.Y(n_153)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_79),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_37),
.B1(n_78),
.B2(n_25),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_156),
.Y(n_162)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_138),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_143),
.B(n_146),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_109),
.B1(n_104),
.B2(n_96),
.Y(n_139)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_113),
.B(n_19),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_104),
.B1(n_113),
.B2(n_32),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_120),
.B1(n_115),
.B2(n_126),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_13),
.B1(n_26),
.B2(n_21),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_153),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_152),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_21),
.B1(n_26),
.B2(n_22),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_24),
.Y(n_168)
);

XOR2x2_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_19),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_121),
.C(n_123),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_169),
.C(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_167),
.Y(n_190)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_127),
.B(n_122),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_164),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_129),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_172),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_168),
.B(n_155),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_118),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_118),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_134),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

OAI221xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_22),
.B1(n_17),
.B2(n_15),
.C(n_23),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_174),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_151),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_182),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_135),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_181),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_154),
.B1(n_142),
.B2(n_146),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_183),
.A2(n_187),
.B1(n_195),
.B2(n_157),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_139),
.C(n_143),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_171),
.C(n_173),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_21),
.B1(n_15),
.B2(n_17),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_36),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_191),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_162),
.B(n_10),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_178),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_23),
.B1(n_14),
.B2(n_17),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_36),
.B1(n_32),
.B2(n_14),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_166),
.B1(n_177),
.B2(n_170),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_196),
.A2(n_180),
.B1(n_186),
.B2(n_184),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_169),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_199),
.C(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_171),
.B(n_164),
.Y(n_202)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_204),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_157),
.B(n_168),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_11),
.Y(n_222)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_162),
.C(n_172),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_55),
.C(n_36),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_0),
.C(n_1),
.Y(n_220)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_191),
.B1(n_55),
.B2(n_2),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_216),
.A2(n_8),
.B1(n_7),
.B2(n_2),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_12),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_222),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_208),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_197),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_223),
.C(n_210),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_198),
.B(n_12),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_210),
.C(n_209),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_11),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_212),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_225),
.B(n_234),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_228),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_211),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_213),
.C(n_230),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_196),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_229),
.A2(n_216),
.B1(n_224),
.B2(n_221),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_220),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_232),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_7),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_0),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_1),
.B(n_3),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_239),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_223),
.C(n_218),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_231),
.B(n_229),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_240),
.B(n_241),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_1),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_244),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_248),
.B(n_238),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_233),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_241),
.Y(n_250)
);

AOI21x1_ASAP7_75t_L g253 ( 
.A1(n_250),
.A2(n_4),
.B(n_5),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_252),
.C(n_247),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_247),
.B(n_236),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_253),
.A2(n_254),
.B(n_246),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_249),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_255),
.A2(n_256),
.B(n_6),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_257),
.Y(n_258)
);

O2A1O1Ixp33_ASAP7_75t_SL g259 ( 
.A1(n_258),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_5),
.C(n_6),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_6),
.Y(n_261)
);


endmodule