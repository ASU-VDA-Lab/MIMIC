module fake_jpeg_2953_n_120 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_19),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_9),
.A2(n_11),
.B(n_15),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_47),
.Y(n_52)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_38),
.Y(n_48)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_50),
.Y(n_54)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_50),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_41),
.B1(n_38),
.B2(n_34),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_56),
.B(n_61),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_37),
.B1(n_34),
.B2(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_35),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_36),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_37),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_41),
.C(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_68),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_69),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_0),
.C(n_1),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_71),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_49),
.B1(n_37),
.B2(n_39),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_18),
.B1(n_29),
.B2(n_28),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_7),
.B(n_8),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_39),
.B1(n_2),
.B2(n_3),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_39),
.B1(n_5),
.B2(n_6),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_20),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_10),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_83),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_82),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_7),
.Y(n_82)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_71),
.CI(n_10),
.CON(n_87),
.SN(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_90),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_8),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_92),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_11),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_13),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_96),
.B(n_21),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_16),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_103),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_84),
.B1(n_86),
.B2(n_83),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_107),
.B1(n_22),
.B2(n_26),
.Y(n_111)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_27),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_75),
.B(n_76),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_90),
.B(n_23),
.C(n_25),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_108),
.B(n_112),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_111),
.A2(n_104),
.B(n_106),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_109),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_113),
.C(n_108),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_100),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_98),
.B(n_110),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_30),
.Y(n_120)
);


endmodule