module fake_jpeg_12247_n_38 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_1),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_20),
.B1(n_19),
.B2(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_17),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_17),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_16),
.C(n_14),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_18),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_28),
.B1(n_29),
.B2(n_23),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_31),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_21),
.C(n_14),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_21),
.B1(n_13),
.B2(n_3),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_33),
.B1(n_4),
.B2(n_6),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_29),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_33)
);

AOI21x1_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_31),
.B(n_33),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_34),
.B1(n_8),
.B2(n_7),
.Y(n_37)
);

OA21x2_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_7),
.B(n_34),
.Y(n_38)
);


endmodule