module fake_jpeg_1600_n_509 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_509);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_509;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_352;
wire n_350;
wire n_150;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_46),
.B(n_50),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_47),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_64),
.Y(n_115)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_55),
.B(n_79),
.Y(n_154)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_16),
.B(n_7),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_73),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_31),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_17),
.B(n_0),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_18),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_77),
.B(n_85),
.Y(n_137)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_33),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_18),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_36),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_93),
.Y(n_149)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g113 ( 
.A(n_87),
.Y(n_113)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_7),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_95),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_17),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_26),
.B(n_0),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_26),
.B(n_0),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_32),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_21),
.B(n_7),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_12),
.Y(n_134)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_58),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_103),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_97),
.A2(n_29),
.B1(n_24),
.B2(n_28),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_105),
.A2(n_41),
.B1(n_28),
.B2(n_24),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_32),
.B1(n_29),
.B2(n_44),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_120),
.A2(n_20),
.B1(n_40),
.B2(n_39),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_51),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_134),
.Y(n_160)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_54),
.Y(n_142)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_59),
.B(n_66),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_158),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_56),
.A2(n_32),
.B1(n_29),
.B2(n_44),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_146),
.A2(n_32),
.B1(n_20),
.B2(n_63),
.Y(n_198)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_73),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_46),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_97),
.A2(n_46),
.B1(n_87),
.B2(n_49),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_157),
.A2(n_53),
.B1(n_62),
.B2(n_89),
.Y(n_204)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_111),
.A2(n_38),
.B1(n_93),
.B2(n_55),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_161),
.A2(n_168),
.B1(n_204),
.B2(n_146),
.Y(n_206)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_163),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_115),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_164),
.B(n_179),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_120),
.A2(n_38),
.B1(n_41),
.B2(n_23),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_170),
.Y(n_235)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_182),
.B(n_201),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

CKINVDCx12_ASAP7_75t_R g186 ( 
.A(n_136),
.Y(n_186)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_79),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_190),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_109),
.B(n_88),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_61),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_20),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_110),
.B(n_92),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_203),
.Y(n_211)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_104),
.Y(n_196)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_101),
.Y(n_197)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_198),
.A2(n_202),
.B1(n_205),
.B2(n_125),
.Y(n_214)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

BUFx8_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_122),
.B(n_90),
.Y(n_201)
);

CKINVDCx9p33_ASAP7_75t_R g202 ( 
.A(n_136),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_106),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_223),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_139),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_239),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_133),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_171),
.B1(n_160),
.B2(n_203),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_113),
.B1(n_187),
.B2(n_183),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_238),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_166),
.B(n_100),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_166),
.B(n_167),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_202),
.A2(n_117),
.B1(n_140),
.B2(n_127),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_242),
.Y(n_298)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_244),
.A2(n_263),
.B1(n_268),
.B2(n_165),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_193),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_246),
.B(n_247),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_193),
.Y(n_247)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_211),
.A2(n_113),
.B1(n_121),
.B2(n_138),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_259),
.Y(n_279)
);

AO22x2_ASAP7_75t_L g252 ( 
.A1(n_206),
.A2(n_167),
.B1(n_187),
.B2(n_183),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_267),
.Y(n_273)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_207),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_253),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_219),
.A2(n_162),
.B1(n_177),
.B2(n_184),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_258),
.B1(n_232),
.B2(n_220),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_215),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_257),
.B(n_266),
.Y(n_293)
);

OAI22x1_ASAP7_75t_L g258 ( 
.A1(n_211),
.A2(n_180),
.B1(n_170),
.B2(n_173),
.Y(n_258)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_178),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_219),
.A2(n_180),
.B(n_145),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_260),
.A2(n_225),
.B(n_68),
.Y(n_291)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_231),
.A2(n_23),
.B1(n_174),
.B2(n_172),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_209),
.B(n_200),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_78),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_230),
.A2(n_199),
.B1(n_196),
.B2(n_173),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_208),
.B(n_135),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_269),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_275),
.Y(n_323)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_245),
.A2(n_211),
.B(n_235),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_282),
.B(n_286),
.Y(n_324)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_284),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_249),
.A2(n_220),
.B(n_235),
.Y(n_285)
);

OR2x6_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_291),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_247),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_222),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_292),
.C(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_289),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_218),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_245),
.A2(n_226),
.B1(n_207),
.B2(n_121),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_294),
.A2(n_250),
.B1(n_258),
.B2(n_249),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_254),
.B(n_234),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_264),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_248),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_257),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_267),
.Y(n_297)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_301),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_302),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_293),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_303),
.B(n_310),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_270),
.A2(n_244),
.B1(n_259),
.B2(n_255),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_304),
.A2(n_306),
.B1(n_312),
.B2(n_320),
.Y(n_337)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_279),
.A2(n_245),
.B1(n_265),
.B2(n_255),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_287),
.C(n_297),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_328),
.C(n_280),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_288),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_288),
.Y(n_311)
);

NOR3xp33_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_319),
.C(n_329),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_279),
.A2(n_255),
.B1(n_252),
.B2(n_267),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_274),
.Y(n_313)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_313),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_274),
.B(n_284),
.Y(n_314)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_314),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_252),
.Y(n_318)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_318),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_299),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_213),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_321),
.B(n_216),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_273),
.A2(n_252),
.B1(n_243),
.B2(n_262),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_330),
.B1(n_298),
.B2(n_212),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_294),
.A2(n_225),
.B1(n_229),
.B2(n_216),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_326),
.A2(n_232),
.B(n_277),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_252),
.Y(n_327)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_327),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_278),
.B(n_280),
.C(n_282),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_299),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_273),
.A2(n_229),
.B1(n_234),
.B2(n_233),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_272),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_332),
.B(n_333),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_215),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_338),
.Y(n_363)
);

OAI32xp33_ASAP7_75t_L g336 ( 
.A1(n_318),
.A2(n_273),
.A3(n_281),
.B1(n_289),
.B2(n_271),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_336),
.B(n_341),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_300),
.B(n_291),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_308),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_346),
.C(n_348),
.Y(n_364)
);

AO21x1_ASAP7_75t_L g341 ( 
.A1(n_309),
.A2(n_285),
.B(n_277),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_343),
.A2(n_344),
.B1(n_353),
.B2(n_358),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_305),
.B(n_221),
.C(n_224),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_212),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_347),
.B(n_354),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_221),
.C(n_210),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_302),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_349),
.B(n_350),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_330),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_313),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_307),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_327),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_210),
.Y(n_354)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_357),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_317),
.B(n_298),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_312),
.A2(n_185),
.B1(n_205),
.B2(n_197),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_359),
.A2(n_320),
.B1(n_329),
.B2(n_319),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_317),
.B(n_232),
.Y(n_361)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_361),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_356),
.A2(n_306),
.B1(n_316),
.B2(n_323),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_365),
.A2(n_369),
.B1(n_359),
.B2(n_344),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_325),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_368),
.B(n_380),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_337),
.A2(n_323),
.B1(n_309),
.B2(n_311),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_371),
.A2(n_374),
.B1(n_382),
.B2(n_384),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_342),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_386),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_337),
.A2(n_309),
.B1(n_307),
.B2(n_322),
.Y(n_374)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_375),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_334),
.B(n_322),
.C(n_309),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_379),
.C(n_348),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_309),
.C(n_140),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_309),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_331),
.Y(n_381)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_381),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_356),
.A2(n_138),
.B1(n_148),
.B2(n_151),
.Y(n_382)
);

XOR2x2_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_217),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_351),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_360),
.A2(n_148),
.B1(n_106),
.B2(n_128),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_340),
.B(n_217),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_346),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_357),
.B(n_22),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_335),
.Y(n_387)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_387),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_335),
.B(n_39),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_8),
.Y(n_411)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_352),
.Y(n_389)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_389),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_393),
.B(n_379),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_394),
.B(n_382),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_364),
.B(n_360),
.C(n_345),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_400),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_397),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_364),
.B(n_345),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_399),
.B(n_403),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_372),
.A2(n_341),
.B(n_343),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_372),
.A2(n_341),
.B(n_355),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_401),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_402),
.A2(n_405),
.B1(n_413),
.B2(n_414),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_336),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_366),
.B(n_349),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_406),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_365),
.A2(n_358),
.B1(n_155),
.B2(n_152),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_169),
.C(n_165),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_407),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_114),
.C(n_47),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_408),
.B(n_409),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_114),
.C(n_152),
.Y(n_409)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_411),
.Y(n_428)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_378),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_362),
.A2(n_155),
.B1(n_151),
.B2(n_131),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_145),
.Y(n_454)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_416),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_392),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_419),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_380),
.C(n_371),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_421),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_374),
.C(n_383),
.Y(n_421)
);

XNOR2x2_ASAP7_75t_SL g423 ( 
.A(n_403),
.B(n_370),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_427),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_367),
.C(n_385),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_425),
.B(n_430),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_391),
.B(n_381),
.C(n_384),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_390),
.A2(n_150),
.B1(n_129),
.B2(n_94),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_431),
.B(n_433),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_432),
.A2(n_435),
.B1(n_413),
.B2(n_395),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_398),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_405),
.A2(n_107),
.B1(n_131),
.B2(n_128),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_418),
.B(n_401),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_439),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_409),
.C(n_391),
.Y(n_439)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_408),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_454),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_417),
.Y(n_442)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_442),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_406),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_443),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_425),
.A2(n_400),
.B(n_393),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_447),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_395),
.C(n_107),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_448),
.C(n_449),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_424),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_429),
.B(n_48),
.C(n_84),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_430),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_451),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_419),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_442),
.A2(n_434),
.B(n_423),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_455),
.A2(n_457),
.B(n_467),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_445),
.A2(n_434),
.B(n_422),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_461),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_438),
.A2(n_415),
.B1(n_428),
.B2(n_74),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_447),
.A2(n_118),
.B1(n_69),
.B2(n_60),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_463),
.A2(n_96),
.B1(n_76),
.B2(n_58),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_441),
.B(n_83),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_466),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_437),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_437),
.A2(n_118),
.B(n_145),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_67),
.C(n_82),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_9),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_468),
.B(n_448),
.Y(n_471)
);

OAI21x1_ASAP7_75t_SL g489 ( 
.A1(n_471),
.A2(n_472),
.B(n_473),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_465),
.A2(n_446),
.B(n_453),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_470),
.B(n_454),
.Y(n_473)
);

MAJx2_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_65),
.C(n_81),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_476),
.B(n_478),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_459),
.A2(n_42),
.B1(n_40),
.B2(n_15),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_456),
.A2(n_42),
.B(n_76),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_479),
.A2(n_483),
.B(n_14),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_480),
.B(n_482),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_455),
.C(n_461),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_9),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_15),
.C(n_45),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_493),
.Y(n_497)
);

AOI322xp5_ASAP7_75t_L g487 ( 
.A1(n_474),
.A2(n_462),
.A3(n_464),
.B1(n_469),
.B2(n_15),
.C1(n_45),
.C2(n_8),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_487),
.A2(n_488),
.B(n_490),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_474),
.B(n_462),
.C(n_15),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_15),
.C(n_45),
.Y(n_490)
);

FAx1_ASAP7_75t_SL g491 ( 
.A(n_477),
.B(n_6),
.CI(n_11),
.CON(n_491),
.SN(n_491)
);

A2O1A1O1Ixp25_ASAP7_75t_L g496 ( 
.A1(n_491),
.A2(n_5),
.B(n_6),
.C(n_9),
.D(n_11),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_473),
.C(n_14),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_492),
.A2(n_491),
.B(n_6),
.Y(n_499)
);

AOI21x1_ASAP7_75t_L g494 ( 
.A1(n_489),
.A2(n_6),
.B(n_10),
.Y(n_494)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_494),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_485),
.A2(n_484),
.B(n_487),
.Y(n_495)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_495),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_496),
.B(n_499),
.Y(n_500)
);

AOI322xp5_ASAP7_75t_L g502 ( 
.A1(n_497),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_9),
.C1(n_11),
.C2(n_498),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_502),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_503),
.B(n_11),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_505),
.B(n_500),
.C(n_501),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_506),
.B(n_504),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_507),
.B(n_2),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_3),
.Y(n_509)
);


endmodule